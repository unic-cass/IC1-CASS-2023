VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_io__corner_bus_overlay
  CLASS PAD ;
  FOREIGN sky130_fd_io__corner_bus_overlay ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 203.665 ;
  SYMMETRY X Y R90 ;
  PIN VSSA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 51.400 23.155 60.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 40.500 1.335 43.750 ;
    END
    PORT
      LAYER met5 ;
        RECT 36.840 0.000 40.085 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 47.735 0.000 56.735 26.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.400 19.575 51.730 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 40.400 1.335 43.850 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 55.310 21.550 56.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 60.070 23.175 60.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.405 0.000 56.735 26.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.645 0.000 52.825 21.555 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.735 0.000 40.185 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.735 0.000 48.065 23.240 ;
    END
  END VSSA
  PIN VSSIO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 179.450 1.435 203.665 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.600 1.600 34.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 25.935 0.000 30.385 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 175.785 0.000 200.000 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.500 1.600 34.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 179.450 1.435 203.665 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.785 0.000 200.000 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.835 0.000 30.485 1.270 ;
    END
  END VSSIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 35.650 1.385 38.900 ;
    END
    PORT
      LAYER met5 ;
        RECT 31.985 0.000 35.235 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 35.550 1.385 39.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.885 0.000 35.335 1.270 ;
    END
  END VSWITCH
  PIN VSSD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.350 1.475 49.800 ;
    END
    PORT
      LAYER met5 ;
        RECT 41.685 0.000 46.135 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.250 1.475 49.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.585 0.000 46.235 1.270 ;
    END
  END VSSD
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.000 1.625 66.250 ;
    END
    PORT
      LAYER met5 ;
        RECT 58.335 0.000 62.585 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 61.900 1.625 66.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.235 0.000 62.685 1.270 ;
    END
  END VSSIO_Q
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 67.850 1.480 72.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 64.185 0.000 68.435 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 67.750 1.480 72.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.085 0.000 68.535 1.270 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 73.700 2.645 98.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.550 1.525 28.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 19.885 0.000 24.335 1.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 70.035 0.000 94.985 1.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.450 1.525 28.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 73.700 2.645 98.665 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.035 0.000 95.000 1.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.785 0.000 24.435 1.270 ;
    END
  END VDDIO
  PIN VDDA
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 18.700 1.470 21.950 ;
    END
    PORT
      LAYER met5 ;
        RECT 15.035 0.000 18.285 1.255 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 18.600 1.470 22.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.935 0.000 18.385 1.255 ;
    END
  END VDDA
  PIN VCCHIB
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 5.800 2.350 11.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.135 0.000 7.385 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 5.700 2.350 11.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.035 0.000 7.485 1.270 ;
    END
  END VCCHIB
  PIN VCCD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 12.650 3.785 17.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 8.985 0.000 13.435 1.270 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.550 3.785 17.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.885 0.000 13.535 1.270 ;
    END
  END VCCD
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 56.790 22.910 59.770 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.125 0.000 56.105 18.475 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 52.030 20.935 55.010 ;
    END
    PORT
      LAYER met4 ;
        RECT 48.365 0.000 51.345 20.875 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met4 ;
        RECT 1.835 179.050 200.000 203.665 ;
        RECT 0.000 99.065 200.000 179.050 ;
        RECT 3.045 73.300 200.000 99.065 ;
        RECT 0.000 72.600 200.000 73.300 ;
        RECT 1.880 67.350 200.000 72.600 ;
        RECT 0.000 66.750 200.000 67.350 ;
        RECT 2.025 61.500 200.000 66.750 ;
        RECT 0.000 60.800 200.000 61.500 ;
        RECT 23.575 59.670 200.000 60.800 ;
        RECT 23.310 56.390 200.000 59.670 ;
        RECT 21.950 54.910 200.000 56.390 ;
        RECT 21.335 51.630 200.000 54.910 ;
        RECT 19.975 51.000 200.000 51.630 ;
        RECT 0.000 50.300 200.000 51.000 ;
        RECT 1.875 44.850 200.000 50.300 ;
        RECT 0.000 44.250 200.000 44.850 ;
        RECT 1.735 40.000 200.000 44.250 ;
        RECT 0.000 39.400 200.000 40.000 ;
        RECT 1.785 35.150 200.000 39.400 ;
        RECT 0.000 34.550 200.000 35.150 ;
        RECT 2.000 29.100 200.000 34.550 ;
        RECT 0.000 28.500 200.000 29.100 ;
        RECT 1.925 27.240 200.000 28.500 ;
        RECT 1.925 23.640 56.005 27.240 ;
        RECT 1.925 23.050 47.335 23.640 ;
        RECT 0.000 22.450 47.335 23.050 ;
        RECT 1.870 18.200 47.335 22.450 ;
        RECT 48.465 21.955 56.005 23.640 ;
        RECT 48.465 21.275 51.245 21.955 ;
        RECT 53.225 18.875 56.005 21.955 ;
        RECT 0.000 17.600 47.335 18.200 ;
        RECT 4.185 12.150 47.335 17.600 ;
        RECT 0.000 11.550 47.335 12.150 ;
        POLYGON 0.000 5.700 0.400 5.700 0.400 5.300 ;
        RECT 0.400 5.300 2.035 5.700 ;
        RECT 2.750 5.300 47.335 11.550 ;
        RECT 0.000 1.670 47.335 5.300 ;
        RECT 0.000 1.255 1.635 1.670 ;
        RECT 7.885 1.255 8.485 1.670 ;
        RECT 13.935 1.655 19.385 1.670 ;
        RECT 13.935 1.255 14.535 1.655 ;
        RECT 18.785 1.255 19.385 1.655 ;
        RECT 24.835 1.255 25.435 1.670 ;
        RECT 30.885 1.255 31.485 1.670 ;
        RECT 35.735 1.255 36.335 1.670 ;
        RECT 40.585 1.255 41.185 1.670 ;
        RECT 46.635 1.255 47.335 1.670 ;
        RECT 57.135 1.920 200.000 27.240 ;
        RECT 57.135 1.670 69.635 1.920 ;
        RECT 57.135 1.255 57.835 1.670 ;
        RECT 63.085 1.255 63.685 1.670 ;
        RECT 68.935 1.255 69.635 1.670 ;
        RECT 95.400 1.670 200.000 1.920 ;
        RECT 95.400 1.255 175.385 1.670 ;
      LAYER met5 ;
        RECT 3.035 177.850 200.000 203.665 ;
        RECT 0.000 100.250 200.000 177.850 ;
        RECT 4.245 72.100 200.000 100.250 ;
        RECT 3.080 67.850 200.000 72.100 ;
        RECT 3.225 62.000 200.000 67.850 ;
        RECT 24.755 49.800 200.000 62.000 ;
        RECT 3.075 43.750 200.000 49.800 ;
        RECT 2.935 40.500 200.000 43.750 ;
        RECT 2.985 35.650 200.000 40.500 ;
        RECT 3.200 28.420 200.000 35.650 ;
        RECT 3.200 28.000 46.135 28.420 ;
        RECT 3.125 21.950 46.135 28.000 ;
        RECT 3.070 18.700 46.135 21.950 ;
        RECT 5.385 11.050 46.135 18.700 ;
        POLYGON 0.000 5.800 1.600 5.800 1.600 4.200 ;
        RECT 1.600 4.200 2.135 5.800 ;
        RECT 3.950 4.200 46.135 11.050 ;
        RECT 0.000 2.870 46.135 4.200 ;
        RECT 58.335 3.120 200.000 28.420 ;
        RECT 58.335 2.870 68.435 3.120 ;
        RECT 96.585 2.870 200.000 3.120 ;
        RECT 0.000 0.000 0.535 2.870 ;
        RECT 15.035 2.855 18.285 2.870 ;
        RECT 96.585 0.000 174.185 2.870 ;
  END
END sky130_fd_io__corner_bus_overlay

#--------EOF---------

MACRO sky130_fd_io__overlay_gpiov2
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_gpiov2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.200 104.560 73.800 166.960 ;
    END
  END PAD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 175.785 80.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 25.935 80.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 25.835 80.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 175.785 80.000 200.000 ;
    END
  END VSSIO
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 78.730 19.885 80.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 70.035 80.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 70.035 80.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 19.785 80.000 24.435 ;
    END
  END VDDIO
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 78.730 2.135 80.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 2.035 80.000 7.485 ;
    END
  END VCCHIB
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 78.730 64.185 80.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 64.085 80.000 68.535 ;
    END
  END VDDIO_Q
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 78.730 8.985 80.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 8.885 80.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
  END VCCD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 78.730 36.840 80.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 78.730 47.735 80.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 80.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 80.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 36.735 80.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 51.645 80.000 52.825 ;
    END
  END VSSA
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 78.730 31.985 80.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 31.885 80.000 35.335 ;
    END
  END VSWITCH
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 78.730 58.335 80.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 58.235 80.000 62.685 ;
    END
  END VSSIO_Q
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 78.730 41.685 80.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.730 41.585 80.000 46.235 ;
    END
  END VSSD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 78.970 15.035 80.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.970 14.935 80.000 18.385 ;
    END
  END VDDA
  PIN AMUXBUS_A
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 80.000 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 80.000 51.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met4 ;
        RECT 1.670 175.385 78.330 200.000 ;
        RECT 0.965 95.400 78.970 175.385 ;
        RECT 1.670 69.635 78.330 95.400 ;
        RECT 0.965 68.935 78.970 69.635 ;
        RECT 1.670 63.685 78.330 68.935 ;
        RECT 0.965 63.085 78.970 63.685 ;
        RECT 1.670 57.835 78.330 63.085 ;
        RECT 0.965 57.135 78.970 57.835 ;
        RECT 1.670 51.745 78.330 52.725 ;
        RECT 0.965 46.635 78.970 47.335 ;
        RECT 1.670 41.185 78.330 46.635 ;
        RECT 0.965 40.585 78.970 41.185 ;
        RECT 1.670 36.335 78.330 40.585 ;
        RECT 0.965 35.735 78.970 36.335 ;
        RECT 1.670 31.485 78.330 35.735 ;
        RECT 0.965 30.885 78.970 31.485 ;
        RECT 1.670 25.435 78.330 30.885 ;
        RECT 0.965 24.835 78.970 25.435 ;
        RECT 1.670 19.385 78.330 24.835 ;
        RECT 0.965 18.785 78.970 19.385 ;
        RECT 1.365 14.535 78.570 18.785 ;
        RECT 0.965 13.935 78.970 14.535 ;
        RECT 1.670 8.485 78.330 13.935 ;
        RECT 0.965 7.885 78.970 8.485 ;
        RECT 1.670 2.035 78.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 77.130 200.000 ;
        RECT 0.000 168.560 80.000 174.185 ;
        RECT 0.000 102.960 9.600 168.560 ;
        RECT 75.400 102.960 80.000 168.560 ;
        RECT 0.000 96.585 80.000 102.960 ;
        RECT 2.870 36.840 77.130 96.585 ;
        RECT 0.000 36.835 80.000 36.840 ;
        RECT 2.870 18.285 77.130 36.835 ;
        RECT 2.565 15.035 77.370 18.285 ;
        RECT 2.870 2.135 77.130 15.035 ;
  END
END sky130_fd_io__overlay_gpiov2

#--------EOF---------

MACRO sky130_fd_io__overlay_vccd_hvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vccd_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
  END VDDIO
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
  END VCCHIB
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
  END VSSA
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 8.890 74.290 13.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 13.260 74.200 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 12.830 74.200 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 12.400 74.200 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 11.970 74.200 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 11.540 74.200 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 11.110 74.200 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 10.680 74.200 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 10.250 74.200 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 9.820 74.200 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 9.390 74.200 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 8.960 74.200 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 13.260 73.795 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 12.830 73.795 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 12.400 73.795 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 11.970 73.795 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 11.540 73.795 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 11.110 73.795 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 10.680 73.795 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 10.250 73.795 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 9.820 73.795 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 9.390 73.795 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 8.960 73.795 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 13.260 73.390 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 12.830 73.390 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 12.400 73.390 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 11.970 73.390 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 11.540 73.390 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 11.110 73.390 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 10.680 73.390 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 10.250 73.390 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 9.820 73.390 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 9.390 73.390 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 8.960 73.390 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 13.260 72.985 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 12.830 72.985 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 12.400 72.985 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 11.970 72.985 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 11.540 72.985 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 11.110 72.985 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 10.680 72.985 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 10.250 72.985 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 9.820 72.985 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 9.390 72.985 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 8.960 72.985 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 13.260 72.580 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 12.830 72.580 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 12.400 72.580 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 11.970 72.580 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 11.540 72.580 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 11.110 72.580 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 10.680 72.580 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 10.250 72.580 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 9.820 72.580 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 9.390 72.580 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 8.960 72.580 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 13.260 72.175 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 12.830 72.175 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 12.400 72.175 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 11.970 72.175 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 11.540 72.175 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 11.110 72.175 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 10.680 72.175 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 10.250 72.175 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 9.820 72.175 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 9.390 72.175 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 8.960 72.175 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 13.260 71.770 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 12.830 71.770 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 12.400 71.770 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 11.970 71.770 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 11.540 71.770 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 11.110 71.770 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 10.680 71.770 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 10.250 71.770 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 9.820 71.770 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 9.390 71.770 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 8.960 71.770 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 13.260 71.365 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 12.830 71.365 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 12.400 71.365 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 11.970 71.365 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 11.540 71.365 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 11.110 71.365 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 10.680 71.365 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 10.250 71.365 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 9.820 71.365 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 9.390 71.365 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 8.960 71.365 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 13.260 70.960 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 12.830 70.960 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 12.400 70.960 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 11.970 70.960 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 11.540 70.960 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 11.110 70.960 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 10.680 70.960 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 10.250 70.960 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 9.820 70.960 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 9.390 70.960 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 8.960 70.960 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 13.260 70.555 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 12.830 70.555 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 12.400 70.555 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 11.970 70.555 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 11.540 70.555 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 11.110 70.555 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 10.680 70.555 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 10.250 70.555 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 9.820 70.555 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 9.390 70.555 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 8.960 70.555 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 13.260 70.150 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 12.830 70.150 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 12.400 70.150 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 11.970 70.150 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 11.540 70.150 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 11.110 70.150 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 10.680 70.150 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 10.250 70.150 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 9.820 70.150 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 9.390 70.150 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 8.960 70.150 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 13.260 69.745 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 12.830 69.745 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 12.400 69.745 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 11.970 69.745 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 11.540 69.745 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 11.110 69.745 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 10.680 69.745 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 10.250 69.745 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 9.820 69.745 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 9.390 69.745 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 8.960 69.745 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 13.260 69.340 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 12.830 69.340 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 12.400 69.340 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 11.970 69.340 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 11.540 69.340 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 11.110 69.340 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 10.680 69.340 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 10.250 69.340 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 9.820 69.340 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 9.390 69.340 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 8.960 69.340 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 13.260 68.935 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 12.830 68.935 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 12.400 68.935 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 11.970 68.935 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 11.540 68.935 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 11.110 68.935 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 10.680 68.935 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 10.250 68.935 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 9.820 68.935 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 9.390 68.935 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 8.960 68.935 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 13.260 68.530 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 12.830 68.530 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 12.400 68.530 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 11.970 68.530 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 11.540 68.530 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 11.110 68.530 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 10.680 68.530 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 10.250 68.530 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 9.820 68.530 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 9.390 68.530 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 8.960 68.530 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 13.260 68.125 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 12.830 68.125 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 12.400 68.125 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 11.970 68.125 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 11.540 68.125 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 11.110 68.125 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 10.680 68.125 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 10.250 68.125 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 9.820 68.125 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 9.390 68.125 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 8.960 68.125 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 13.260 67.720 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 12.830 67.720 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 12.400 67.720 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 11.970 67.720 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 11.540 67.720 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 11.110 67.720 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 10.680 67.720 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 10.250 67.720 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 9.820 67.720 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 9.390 67.720 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 8.960 67.720 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 13.260 67.315 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 12.830 67.315 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 12.400 67.315 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 11.970 67.315 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 11.540 67.315 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 11.110 67.315 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 10.680 67.315 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 10.250 67.315 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 9.820 67.315 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 9.390 67.315 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 8.960 67.315 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 13.260 66.910 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 12.830 66.910 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 12.400 66.910 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 11.970 66.910 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 11.540 66.910 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 11.110 66.910 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 10.680 66.910 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 10.250 66.910 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 9.820 66.910 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 9.390 66.910 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 8.960 66.910 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 13.260 66.505 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 12.830 66.505 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 12.400 66.505 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 11.970 66.505 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 11.540 66.505 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 11.110 66.505 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 10.680 66.505 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 10.250 66.505 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 9.820 66.505 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 9.390 66.505 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 8.960 66.505 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 13.260 66.100 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 12.830 66.100 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 12.400 66.100 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 11.970 66.100 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 11.540 66.100 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 11.110 66.100 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 10.680 66.100 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 10.250 66.100 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 9.820 66.100 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 9.390 66.100 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 8.960 66.100 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 13.260 65.695 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 12.830 65.695 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 12.400 65.695 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 11.970 65.695 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 11.540 65.695 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 11.110 65.695 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 10.680 65.695 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 10.250 65.695 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 9.820 65.695 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 9.390 65.695 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 8.960 65.695 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 13.260 65.290 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 12.830 65.290 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 12.400 65.290 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 11.970 65.290 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 11.540 65.290 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 11.110 65.290 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 10.680 65.290 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 10.250 65.290 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 9.820 65.290 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 9.390 65.290 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 8.960 65.290 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 13.260 64.885 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 12.830 64.885 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 12.400 64.885 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 11.970 64.885 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 11.540 64.885 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 11.110 64.885 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 10.680 64.885 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 10.250 64.885 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 9.820 64.885 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 9.390 64.885 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 8.960 64.885 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 13.260 64.480 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 12.830 64.480 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 12.400 64.480 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 11.970 64.480 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 11.540 64.480 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 11.110 64.480 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 10.680 64.480 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 10.250 64.480 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 9.820 64.480 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 9.390 64.480 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 8.960 64.480 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 13.260 64.075 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 12.830 64.075 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 12.400 64.075 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 11.970 64.075 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 11.540 64.075 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 11.110 64.075 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 10.680 64.075 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 10.250 64.075 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 9.820 64.075 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 9.390 64.075 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 8.960 64.075 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 13.260 63.670 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 12.830 63.670 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 12.400 63.670 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 11.970 63.670 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 11.540 63.670 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 11.110 63.670 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 10.680 63.670 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 10.250 63.670 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 9.820 63.670 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 9.390 63.670 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 8.960 63.670 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 13.260 63.265 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 12.830 63.265 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 12.400 63.265 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 11.970 63.265 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 11.540 63.265 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 11.110 63.265 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 10.680 63.265 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 10.250 63.265 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 9.820 63.265 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 9.390 63.265 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 8.960 63.265 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 13.260 62.860 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 12.830 62.860 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 12.400 62.860 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 11.970 62.860 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 11.540 62.860 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 11.110 62.860 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 10.680 62.860 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 10.250 62.860 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 9.820 62.860 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 9.390 62.860 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 8.960 62.860 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 13.260 62.455 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 12.830 62.455 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 12.400 62.455 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 11.970 62.455 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 11.540 62.455 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 11.110 62.455 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 10.680 62.455 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 10.250 62.455 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 9.820 62.455 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 9.390 62.455 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 8.960 62.455 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 13.260 62.050 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 12.830 62.050 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 12.400 62.050 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 11.970 62.050 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 11.540 62.050 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 11.110 62.050 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 10.680 62.050 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 10.250 62.050 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 9.820 62.050 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 9.390 62.050 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 8.960 62.050 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 13.260 61.645 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 12.830 61.645 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 12.400 61.645 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 11.970 61.645 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 11.540 61.645 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 11.110 61.645 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 10.680 61.645 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 10.250 61.645 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 9.820 61.645 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 9.390 61.645 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 8.960 61.645 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 13.260 61.240 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 12.830 61.240 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 12.400 61.240 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 11.970 61.240 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 11.540 61.240 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 11.110 61.240 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 10.680 61.240 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 10.250 61.240 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 9.820 61.240 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 9.390 61.240 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 8.960 61.240 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 13.260 60.835 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 12.830 60.835 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 12.400 60.835 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 11.970 60.835 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 11.540 60.835 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 11.110 60.835 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 10.680 60.835 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 10.250 60.835 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 9.820 60.835 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 9.390 60.835 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 8.960 60.835 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 13.260 60.430 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 12.830 60.430 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 12.400 60.430 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 11.970 60.430 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 11.540 60.430 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 11.110 60.430 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 10.680 60.430 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 10.250 60.430 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 9.820 60.430 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 9.390 60.430 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 8.960 60.430 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 13.260 60.025 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 12.830 60.025 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 12.400 60.025 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 11.970 60.025 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 11.540 60.025 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 11.110 60.025 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 10.680 60.025 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 10.250 60.025 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 9.820 60.025 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 9.390 60.025 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 8.960 60.025 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 13.260 59.620 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 12.830 59.620 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 12.400 59.620 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 11.970 59.620 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 11.540 59.620 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 11.110 59.620 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 10.680 59.620 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 10.250 59.620 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 9.820 59.620 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 9.390 59.620 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 8.960 59.620 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 13.260 59.215 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 12.830 59.215 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 12.400 59.215 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 11.970 59.215 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 11.540 59.215 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 11.110 59.215 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 10.680 59.215 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 10.250 59.215 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 9.820 59.215 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 9.390 59.215 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 8.960 59.215 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 13.260 58.810 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 12.830 58.810 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 12.400 58.810 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 11.970 58.810 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 11.540 58.810 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 11.110 58.810 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 10.680 58.810 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 10.250 58.810 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 9.820 58.810 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 9.390 58.810 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 8.960 58.810 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 13.260 58.405 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 12.830 58.405 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 12.400 58.405 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 11.970 58.405 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 11.540 58.405 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 11.110 58.405 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 10.680 58.405 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 10.250 58.405 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 9.820 58.405 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 9.390 58.405 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 8.960 58.405 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 13.260 58.000 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 12.830 58.000 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 12.400 58.000 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 11.970 58.000 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 11.540 58.000 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 11.110 58.000 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 10.680 58.000 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 10.250 58.000 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 9.820 58.000 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 9.390 58.000 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 8.960 58.000 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 13.260 57.595 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 12.830 57.595 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 12.400 57.595 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 11.970 57.595 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 11.540 57.595 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 11.110 57.595 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 10.680 57.595 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 10.250 57.595 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 9.820 57.595 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 9.390 57.595 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 8.960 57.595 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 13.260 57.190 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 12.830 57.190 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 12.400 57.190 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 11.970 57.190 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 11.540 57.190 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 11.110 57.190 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 10.680 57.190 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 10.250 57.190 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 9.820 57.190 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 9.390 57.190 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 8.960 57.190 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 13.260 56.785 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 12.830 56.785 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 12.400 56.785 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 11.970 56.785 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 11.540 56.785 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 11.110 56.785 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 10.680 56.785 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 10.250 56.785 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 9.820 56.785 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 9.390 56.785 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 8.960 56.785 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 13.260 56.380 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 12.830 56.380 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 12.400 56.380 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 11.970 56.380 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 11.540 56.380 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 11.110 56.380 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 10.680 56.380 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 10.250 56.380 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 9.820 56.380 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 9.390 56.380 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 8.960 56.380 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 13.260 55.975 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 12.830 55.975 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 12.400 55.975 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 11.970 55.975 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 11.540 55.975 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 11.110 55.975 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 10.680 55.975 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 10.250 55.975 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 9.820 55.975 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 9.390 55.975 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 8.960 55.975 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 13.260 55.570 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 12.830 55.570 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 12.400 55.570 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 11.970 55.570 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 11.540 55.570 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 11.110 55.570 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 10.680 55.570 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 10.250 55.570 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 9.820 55.570 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 9.390 55.570 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 8.960 55.570 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 13.260 55.165 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 12.830 55.165 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 12.400 55.165 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 11.970 55.165 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 11.540 55.165 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 11.110 55.165 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 10.680 55.165 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 10.250 55.165 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 9.820 55.165 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 9.390 55.165 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 8.960 55.165 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 13.260 54.760 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 12.830 54.760 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 12.400 54.760 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 11.970 54.760 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 11.540 54.760 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 11.110 54.760 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 10.680 54.760 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 10.250 54.760 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 9.820 54.760 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 9.390 54.760 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 8.960 54.760 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 13.260 54.355 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 12.830 54.355 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 12.400 54.355 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 11.970 54.355 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 11.540 54.355 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 11.110 54.355 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 10.680 54.355 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 10.250 54.355 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 9.820 54.355 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 9.390 54.355 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 8.960 54.355 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 13.260 53.950 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 12.830 53.950 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 12.400 53.950 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 11.970 53.950 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 11.540 53.950 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 11.110 53.950 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 10.680 53.950 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 10.250 53.950 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 9.820 53.950 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 9.390 53.950 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 8.960 53.950 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 13.260 53.545 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 12.830 53.545 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 12.400 53.545 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 11.970 53.545 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 11.540 53.545 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 11.110 53.545 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 10.680 53.545 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 10.250 53.545 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 9.820 53.545 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 9.390 53.545 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 8.960 53.545 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 13.260 53.140 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 12.830 53.140 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 12.400 53.140 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 11.970 53.140 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 11.540 53.140 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 11.110 53.140 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 10.680 53.140 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 10.250 53.140 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 9.820 53.140 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 9.390 53.140 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 8.960 53.140 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 13.260 52.730 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 12.830 52.730 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 12.400 52.730 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 11.970 52.730 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 11.540 52.730 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 11.110 52.730 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 10.680 52.730 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 10.250 52.730 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 9.820 52.730 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 9.390 52.730 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 8.960 52.730 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 13.260 52.320 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 12.830 52.320 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 12.400 52.320 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 11.970 52.320 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 11.540 52.320 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 11.110 52.320 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 10.680 52.320 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 10.250 52.320 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 9.820 52.320 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 9.390 52.320 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 8.960 52.320 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 13.260 51.910 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 12.830 51.910 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 12.400 51.910 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 11.970 51.910 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 11.540 51.910 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 11.110 51.910 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 10.680 51.910 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 10.250 51.910 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 9.820 51.910 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 9.390 51.910 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 8.960 51.910 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 13.260 51.500 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 12.830 51.500 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 12.400 51.500 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 11.970 51.500 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 11.540 51.500 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 11.110 51.500 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 10.680 51.500 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 10.250 51.500 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 9.820 51.500 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 9.390 51.500 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 8.960 51.500 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 13.260 51.090 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 12.830 51.090 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 12.400 51.090 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 11.970 51.090 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 11.540 51.090 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 11.110 51.090 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 10.680 51.090 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 10.250 51.090 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 9.820 51.090 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 9.390 51.090 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 8.960 51.090 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 13.260 50.680 13.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 12.830 50.680 13.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 12.400 50.680 12.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 11.970 50.680 12.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 11.540 50.680 11.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 11.110 50.680 11.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 10.680 50.680 10.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 10.250 50.680 10.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 9.820 50.680 10.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 9.390 50.680 9.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 8.960 50.680 9.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 13.200 24.365 13.520 ;
      LAYER met4 ;
        RECT 24.045 13.200 24.365 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 12.770 24.365 13.090 ;
      LAYER met4 ;
        RECT 24.045 12.770 24.365 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 12.340 24.365 12.660 ;
      LAYER met4 ;
        RECT 24.045 12.340 24.365 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 11.910 24.365 12.230 ;
      LAYER met4 ;
        RECT 24.045 11.910 24.365 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 11.480 24.365 11.800 ;
      LAYER met4 ;
        RECT 24.045 11.480 24.365 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 11.050 24.365 11.370 ;
      LAYER met4 ;
        RECT 24.045 11.050 24.365 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 10.620 24.365 10.940 ;
      LAYER met4 ;
        RECT 24.045 10.620 24.365 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 10.190 24.365 10.510 ;
      LAYER met4 ;
        RECT 24.045 10.190 24.365 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 9.760 24.365 10.080 ;
      LAYER met4 ;
        RECT 24.045 9.760 24.365 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 9.330 24.365 9.650 ;
      LAYER met4 ;
        RECT 24.045 9.330 24.365 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 8.900 24.365 9.220 ;
      LAYER met4 ;
        RECT 24.045 8.900 24.365 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 13.200 23.960 13.520 ;
      LAYER met4 ;
        RECT 23.640 13.200 23.960 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 12.770 23.960 13.090 ;
      LAYER met4 ;
        RECT 23.640 12.770 23.960 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 12.340 23.960 12.660 ;
      LAYER met4 ;
        RECT 23.640 12.340 23.960 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 11.910 23.960 12.230 ;
      LAYER met4 ;
        RECT 23.640 11.910 23.960 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 11.480 23.960 11.800 ;
      LAYER met4 ;
        RECT 23.640 11.480 23.960 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 11.050 23.960 11.370 ;
      LAYER met4 ;
        RECT 23.640 11.050 23.960 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 10.620 23.960 10.940 ;
      LAYER met4 ;
        RECT 23.640 10.620 23.960 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 10.190 23.960 10.510 ;
      LAYER met4 ;
        RECT 23.640 10.190 23.960 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 9.760 23.960 10.080 ;
      LAYER met4 ;
        RECT 23.640 9.760 23.960 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 9.330 23.960 9.650 ;
      LAYER met4 ;
        RECT 23.640 9.330 23.960 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 8.900 23.960 9.220 ;
      LAYER met4 ;
        RECT 23.640 8.900 23.960 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 13.200 23.555 13.520 ;
      LAYER met4 ;
        RECT 23.235 13.200 23.555 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 12.770 23.555 13.090 ;
      LAYER met4 ;
        RECT 23.235 12.770 23.555 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 12.340 23.555 12.660 ;
      LAYER met4 ;
        RECT 23.235 12.340 23.555 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 11.910 23.555 12.230 ;
      LAYER met4 ;
        RECT 23.235 11.910 23.555 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 11.480 23.555 11.800 ;
      LAYER met4 ;
        RECT 23.235 11.480 23.555 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 11.050 23.555 11.370 ;
      LAYER met4 ;
        RECT 23.235 11.050 23.555 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 10.620 23.555 10.940 ;
      LAYER met4 ;
        RECT 23.235 10.620 23.555 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 10.190 23.555 10.510 ;
      LAYER met4 ;
        RECT 23.235 10.190 23.555 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 9.760 23.555 10.080 ;
      LAYER met4 ;
        RECT 23.235 9.760 23.555 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 9.330 23.555 9.650 ;
      LAYER met4 ;
        RECT 23.235 9.330 23.555 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 8.900 23.555 9.220 ;
      LAYER met4 ;
        RECT 23.235 8.900 23.555 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 13.200 23.150 13.520 ;
      LAYER met4 ;
        RECT 22.830 13.200 23.150 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 12.770 23.150 13.090 ;
      LAYER met4 ;
        RECT 22.830 12.770 23.150 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 12.340 23.150 12.660 ;
      LAYER met4 ;
        RECT 22.830 12.340 23.150 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 11.910 23.150 12.230 ;
      LAYER met4 ;
        RECT 22.830 11.910 23.150 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 11.480 23.150 11.800 ;
      LAYER met4 ;
        RECT 22.830 11.480 23.150 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 11.050 23.150 11.370 ;
      LAYER met4 ;
        RECT 22.830 11.050 23.150 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 10.620 23.150 10.940 ;
      LAYER met4 ;
        RECT 22.830 10.620 23.150 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 10.190 23.150 10.510 ;
      LAYER met4 ;
        RECT 22.830 10.190 23.150 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 9.760 23.150 10.080 ;
      LAYER met4 ;
        RECT 22.830 9.760 23.150 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 9.330 23.150 9.650 ;
      LAYER met4 ;
        RECT 22.830 9.330 23.150 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 8.900 23.150 9.220 ;
      LAYER met4 ;
        RECT 22.830 8.900 23.150 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 13.200 22.745 13.520 ;
      LAYER met4 ;
        RECT 22.425 13.200 22.745 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 12.770 22.745 13.090 ;
      LAYER met4 ;
        RECT 22.425 12.770 22.745 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 12.340 22.745 12.660 ;
      LAYER met4 ;
        RECT 22.425 12.340 22.745 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 11.910 22.745 12.230 ;
      LAYER met4 ;
        RECT 22.425 11.910 22.745 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 11.480 22.745 11.800 ;
      LAYER met4 ;
        RECT 22.425 11.480 22.745 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 11.050 22.745 11.370 ;
      LAYER met4 ;
        RECT 22.425 11.050 22.745 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 10.620 22.745 10.940 ;
      LAYER met4 ;
        RECT 22.425 10.620 22.745 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 10.190 22.745 10.510 ;
      LAYER met4 ;
        RECT 22.425 10.190 22.745 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 9.760 22.745 10.080 ;
      LAYER met4 ;
        RECT 22.425 9.760 22.745 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 9.330 22.745 9.650 ;
      LAYER met4 ;
        RECT 22.425 9.330 22.745 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 8.900 22.745 9.220 ;
      LAYER met4 ;
        RECT 22.425 8.900 22.745 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 13.200 22.340 13.520 ;
      LAYER met4 ;
        RECT 22.020 13.200 22.340 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 12.770 22.340 13.090 ;
      LAYER met4 ;
        RECT 22.020 12.770 22.340 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 12.340 22.340 12.660 ;
      LAYER met4 ;
        RECT 22.020 12.340 22.340 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 11.910 22.340 12.230 ;
      LAYER met4 ;
        RECT 22.020 11.910 22.340 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 11.480 22.340 11.800 ;
      LAYER met4 ;
        RECT 22.020 11.480 22.340 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 11.050 22.340 11.370 ;
      LAYER met4 ;
        RECT 22.020 11.050 22.340 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 10.620 22.340 10.940 ;
      LAYER met4 ;
        RECT 22.020 10.620 22.340 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 10.190 22.340 10.510 ;
      LAYER met4 ;
        RECT 22.020 10.190 22.340 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 9.760 22.340 10.080 ;
      LAYER met4 ;
        RECT 22.020 9.760 22.340 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 9.330 22.340 9.650 ;
      LAYER met4 ;
        RECT 22.020 9.330 22.340 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 8.900 22.340 9.220 ;
      LAYER met4 ;
        RECT 22.020 8.900 22.340 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 13.200 21.935 13.520 ;
      LAYER met4 ;
        RECT 21.615 13.200 21.935 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 12.770 21.935 13.090 ;
      LAYER met4 ;
        RECT 21.615 12.770 21.935 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 12.340 21.935 12.660 ;
      LAYER met4 ;
        RECT 21.615 12.340 21.935 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 11.910 21.935 12.230 ;
      LAYER met4 ;
        RECT 21.615 11.910 21.935 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 11.480 21.935 11.800 ;
      LAYER met4 ;
        RECT 21.615 11.480 21.935 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 11.050 21.935 11.370 ;
      LAYER met4 ;
        RECT 21.615 11.050 21.935 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 10.620 21.935 10.940 ;
      LAYER met4 ;
        RECT 21.615 10.620 21.935 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 10.190 21.935 10.510 ;
      LAYER met4 ;
        RECT 21.615 10.190 21.935 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 9.760 21.935 10.080 ;
      LAYER met4 ;
        RECT 21.615 9.760 21.935 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 9.330 21.935 9.650 ;
      LAYER met4 ;
        RECT 21.615 9.330 21.935 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 8.900 21.935 9.220 ;
      LAYER met4 ;
        RECT 21.615 8.900 21.935 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 13.200 21.530 13.520 ;
      LAYER met4 ;
        RECT 21.210 13.200 21.530 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 12.770 21.530 13.090 ;
      LAYER met4 ;
        RECT 21.210 12.770 21.530 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 12.340 21.530 12.660 ;
      LAYER met4 ;
        RECT 21.210 12.340 21.530 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 11.910 21.530 12.230 ;
      LAYER met4 ;
        RECT 21.210 11.910 21.530 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 11.480 21.530 11.800 ;
      LAYER met4 ;
        RECT 21.210 11.480 21.530 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 11.050 21.530 11.370 ;
      LAYER met4 ;
        RECT 21.210 11.050 21.530 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 10.620 21.530 10.940 ;
      LAYER met4 ;
        RECT 21.210 10.620 21.530 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 10.190 21.530 10.510 ;
      LAYER met4 ;
        RECT 21.210 10.190 21.530 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 9.760 21.530 10.080 ;
      LAYER met4 ;
        RECT 21.210 9.760 21.530 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 9.330 21.530 9.650 ;
      LAYER met4 ;
        RECT 21.210 9.330 21.530 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 8.900 21.530 9.220 ;
      LAYER met4 ;
        RECT 21.210 8.900 21.530 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 13.200 21.125 13.520 ;
      LAYER met4 ;
        RECT 20.805 13.200 21.125 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 12.770 21.125 13.090 ;
      LAYER met4 ;
        RECT 20.805 12.770 21.125 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 12.340 21.125 12.660 ;
      LAYER met4 ;
        RECT 20.805 12.340 21.125 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 11.910 21.125 12.230 ;
      LAYER met4 ;
        RECT 20.805 11.910 21.125 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 11.480 21.125 11.800 ;
      LAYER met4 ;
        RECT 20.805 11.480 21.125 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 11.050 21.125 11.370 ;
      LAYER met4 ;
        RECT 20.805 11.050 21.125 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 10.620 21.125 10.940 ;
      LAYER met4 ;
        RECT 20.805 10.620 21.125 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 10.190 21.125 10.510 ;
      LAYER met4 ;
        RECT 20.805 10.190 21.125 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 9.760 21.125 10.080 ;
      LAYER met4 ;
        RECT 20.805 9.760 21.125 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 9.330 21.125 9.650 ;
      LAYER met4 ;
        RECT 20.805 9.330 21.125 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 8.900 21.125 9.220 ;
      LAYER met4 ;
        RECT 20.805 8.900 21.125 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 13.200 20.720 13.520 ;
      LAYER met4 ;
        RECT 20.400 13.200 20.720 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 12.770 20.720 13.090 ;
      LAYER met4 ;
        RECT 20.400 12.770 20.720 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 12.340 20.720 12.660 ;
      LAYER met4 ;
        RECT 20.400 12.340 20.720 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 11.910 20.720 12.230 ;
      LAYER met4 ;
        RECT 20.400 11.910 20.720 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 11.480 20.720 11.800 ;
      LAYER met4 ;
        RECT 20.400 11.480 20.720 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 11.050 20.720 11.370 ;
      LAYER met4 ;
        RECT 20.400 11.050 20.720 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 10.620 20.720 10.940 ;
      LAYER met4 ;
        RECT 20.400 10.620 20.720 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 10.190 20.720 10.510 ;
      LAYER met4 ;
        RECT 20.400 10.190 20.720 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 9.760 20.720 10.080 ;
      LAYER met4 ;
        RECT 20.400 9.760 20.720 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 9.330 20.720 9.650 ;
      LAYER met4 ;
        RECT 20.400 9.330 20.720 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 8.900 20.720 9.220 ;
      LAYER met4 ;
        RECT 20.400 8.900 20.720 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 13.200 20.315 13.520 ;
      LAYER met4 ;
        RECT 19.995 13.200 20.315 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 12.770 20.315 13.090 ;
      LAYER met4 ;
        RECT 19.995 12.770 20.315 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 12.340 20.315 12.660 ;
      LAYER met4 ;
        RECT 19.995 12.340 20.315 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 11.910 20.315 12.230 ;
      LAYER met4 ;
        RECT 19.995 11.910 20.315 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 11.480 20.315 11.800 ;
      LAYER met4 ;
        RECT 19.995 11.480 20.315 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 11.050 20.315 11.370 ;
      LAYER met4 ;
        RECT 19.995 11.050 20.315 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 10.620 20.315 10.940 ;
      LAYER met4 ;
        RECT 19.995 10.620 20.315 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 10.190 20.315 10.510 ;
      LAYER met4 ;
        RECT 19.995 10.190 20.315 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 9.760 20.315 10.080 ;
      LAYER met4 ;
        RECT 19.995 9.760 20.315 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 9.330 20.315 9.650 ;
      LAYER met4 ;
        RECT 19.995 9.330 20.315 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 8.900 20.315 9.220 ;
      LAYER met4 ;
        RECT 19.995 8.900 20.315 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 13.200 19.910 13.520 ;
      LAYER met4 ;
        RECT 19.590 13.200 19.910 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 12.770 19.910 13.090 ;
      LAYER met4 ;
        RECT 19.590 12.770 19.910 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 12.340 19.910 12.660 ;
      LAYER met4 ;
        RECT 19.590 12.340 19.910 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 11.910 19.910 12.230 ;
      LAYER met4 ;
        RECT 19.590 11.910 19.910 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 11.480 19.910 11.800 ;
      LAYER met4 ;
        RECT 19.590 11.480 19.910 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 11.050 19.910 11.370 ;
      LAYER met4 ;
        RECT 19.590 11.050 19.910 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 10.620 19.910 10.940 ;
      LAYER met4 ;
        RECT 19.590 10.620 19.910 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 10.190 19.910 10.510 ;
      LAYER met4 ;
        RECT 19.590 10.190 19.910 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 9.760 19.910 10.080 ;
      LAYER met4 ;
        RECT 19.590 9.760 19.910 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 9.330 19.910 9.650 ;
      LAYER met4 ;
        RECT 19.590 9.330 19.910 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 8.900 19.910 9.220 ;
      LAYER met4 ;
        RECT 19.590 8.900 19.910 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 13.200 19.505 13.520 ;
      LAYER met4 ;
        RECT 19.185 13.200 19.505 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 12.770 19.505 13.090 ;
      LAYER met4 ;
        RECT 19.185 12.770 19.505 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 12.340 19.505 12.660 ;
      LAYER met4 ;
        RECT 19.185 12.340 19.505 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 11.910 19.505 12.230 ;
      LAYER met4 ;
        RECT 19.185 11.910 19.505 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 11.480 19.505 11.800 ;
      LAYER met4 ;
        RECT 19.185 11.480 19.505 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 11.050 19.505 11.370 ;
      LAYER met4 ;
        RECT 19.185 11.050 19.505 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 10.620 19.505 10.940 ;
      LAYER met4 ;
        RECT 19.185 10.620 19.505 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 10.190 19.505 10.510 ;
      LAYER met4 ;
        RECT 19.185 10.190 19.505 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 9.760 19.505 10.080 ;
      LAYER met4 ;
        RECT 19.185 9.760 19.505 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 9.330 19.505 9.650 ;
      LAYER met4 ;
        RECT 19.185 9.330 19.505 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 8.900 19.505 9.220 ;
      LAYER met4 ;
        RECT 19.185 8.900 19.505 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 13.200 19.100 13.520 ;
      LAYER met4 ;
        RECT 18.780 13.200 19.100 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 12.770 19.100 13.090 ;
      LAYER met4 ;
        RECT 18.780 12.770 19.100 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 12.340 19.100 12.660 ;
      LAYER met4 ;
        RECT 18.780 12.340 19.100 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 11.910 19.100 12.230 ;
      LAYER met4 ;
        RECT 18.780 11.910 19.100 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 11.480 19.100 11.800 ;
      LAYER met4 ;
        RECT 18.780 11.480 19.100 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 11.050 19.100 11.370 ;
      LAYER met4 ;
        RECT 18.780 11.050 19.100 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 10.620 19.100 10.940 ;
      LAYER met4 ;
        RECT 18.780 10.620 19.100 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 10.190 19.100 10.510 ;
      LAYER met4 ;
        RECT 18.780 10.190 19.100 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 9.760 19.100 10.080 ;
      LAYER met4 ;
        RECT 18.780 9.760 19.100 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 9.330 19.100 9.650 ;
      LAYER met4 ;
        RECT 18.780 9.330 19.100 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 8.900 19.100 9.220 ;
      LAYER met4 ;
        RECT 18.780 8.900 19.100 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 13.200 18.695 13.520 ;
      LAYER met4 ;
        RECT 18.375 13.200 18.695 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 12.770 18.695 13.090 ;
      LAYER met4 ;
        RECT 18.375 12.770 18.695 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 12.340 18.695 12.660 ;
      LAYER met4 ;
        RECT 18.375 12.340 18.695 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 11.910 18.695 12.230 ;
      LAYER met4 ;
        RECT 18.375 11.910 18.695 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 11.480 18.695 11.800 ;
      LAYER met4 ;
        RECT 18.375 11.480 18.695 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 11.050 18.695 11.370 ;
      LAYER met4 ;
        RECT 18.375 11.050 18.695 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 10.620 18.695 10.940 ;
      LAYER met4 ;
        RECT 18.375 10.620 18.695 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 10.190 18.695 10.510 ;
      LAYER met4 ;
        RECT 18.375 10.190 18.695 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 9.760 18.695 10.080 ;
      LAYER met4 ;
        RECT 18.375 9.760 18.695 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 9.330 18.695 9.650 ;
      LAYER met4 ;
        RECT 18.375 9.330 18.695 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 8.900 18.695 9.220 ;
      LAYER met4 ;
        RECT 18.375 8.900 18.695 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 13.200 18.290 13.520 ;
      LAYER met4 ;
        RECT 17.970 13.200 18.290 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 12.770 18.290 13.090 ;
      LAYER met4 ;
        RECT 17.970 12.770 18.290 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 12.340 18.290 12.660 ;
      LAYER met4 ;
        RECT 17.970 12.340 18.290 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 11.910 18.290 12.230 ;
      LAYER met4 ;
        RECT 17.970 11.910 18.290 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 11.480 18.290 11.800 ;
      LAYER met4 ;
        RECT 17.970 11.480 18.290 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 11.050 18.290 11.370 ;
      LAYER met4 ;
        RECT 17.970 11.050 18.290 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 10.620 18.290 10.940 ;
      LAYER met4 ;
        RECT 17.970 10.620 18.290 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 10.190 18.290 10.510 ;
      LAYER met4 ;
        RECT 17.970 10.190 18.290 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 9.760 18.290 10.080 ;
      LAYER met4 ;
        RECT 17.970 9.760 18.290 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 9.330 18.290 9.650 ;
      LAYER met4 ;
        RECT 17.970 9.330 18.290 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 8.900 18.290 9.220 ;
      LAYER met4 ;
        RECT 17.970 8.900 18.290 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 13.200 17.885 13.520 ;
      LAYER met4 ;
        RECT 17.565 13.200 17.885 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 12.770 17.885 13.090 ;
      LAYER met4 ;
        RECT 17.565 12.770 17.885 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 12.340 17.885 12.660 ;
      LAYER met4 ;
        RECT 17.565 12.340 17.885 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 11.910 17.885 12.230 ;
      LAYER met4 ;
        RECT 17.565 11.910 17.885 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 11.480 17.885 11.800 ;
      LAYER met4 ;
        RECT 17.565 11.480 17.885 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 11.050 17.885 11.370 ;
      LAYER met4 ;
        RECT 17.565 11.050 17.885 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 10.620 17.885 10.940 ;
      LAYER met4 ;
        RECT 17.565 10.620 17.885 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 10.190 17.885 10.510 ;
      LAYER met4 ;
        RECT 17.565 10.190 17.885 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 9.760 17.885 10.080 ;
      LAYER met4 ;
        RECT 17.565 9.760 17.885 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 9.330 17.885 9.650 ;
      LAYER met4 ;
        RECT 17.565 9.330 17.885 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 8.900 17.885 9.220 ;
      LAYER met4 ;
        RECT 17.565 8.900 17.885 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 13.200 17.480 13.520 ;
      LAYER met4 ;
        RECT 17.160 13.200 17.480 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 12.770 17.480 13.090 ;
      LAYER met4 ;
        RECT 17.160 12.770 17.480 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 12.340 17.480 12.660 ;
      LAYER met4 ;
        RECT 17.160 12.340 17.480 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 11.910 17.480 12.230 ;
      LAYER met4 ;
        RECT 17.160 11.910 17.480 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 11.480 17.480 11.800 ;
      LAYER met4 ;
        RECT 17.160 11.480 17.480 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 11.050 17.480 11.370 ;
      LAYER met4 ;
        RECT 17.160 11.050 17.480 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 10.620 17.480 10.940 ;
      LAYER met4 ;
        RECT 17.160 10.620 17.480 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 10.190 17.480 10.510 ;
      LAYER met4 ;
        RECT 17.160 10.190 17.480 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 9.760 17.480 10.080 ;
      LAYER met4 ;
        RECT 17.160 9.760 17.480 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 9.330 17.480 9.650 ;
      LAYER met4 ;
        RECT 17.160 9.330 17.480 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 8.900 17.480 9.220 ;
      LAYER met4 ;
        RECT 17.160 8.900 17.480 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 13.200 17.075 13.520 ;
      LAYER met4 ;
        RECT 16.755 13.200 17.075 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 12.770 17.075 13.090 ;
      LAYER met4 ;
        RECT 16.755 12.770 17.075 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 12.340 17.075 12.660 ;
      LAYER met4 ;
        RECT 16.755 12.340 17.075 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 11.910 17.075 12.230 ;
      LAYER met4 ;
        RECT 16.755 11.910 17.075 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 11.480 17.075 11.800 ;
      LAYER met4 ;
        RECT 16.755 11.480 17.075 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 11.050 17.075 11.370 ;
      LAYER met4 ;
        RECT 16.755 11.050 17.075 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 10.620 17.075 10.940 ;
      LAYER met4 ;
        RECT 16.755 10.620 17.075 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 10.190 17.075 10.510 ;
      LAYER met4 ;
        RECT 16.755 10.190 17.075 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 9.760 17.075 10.080 ;
      LAYER met4 ;
        RECT 16.755 9.760 17.075 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 9.330 17.075 9.650 ;
      LAYER met4 ;
        RECT 16.755 9.330 17.075 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 8.900 17.075 9.220 ;
      LAYER met4 ;
        RECT 16.755 8.900 17.075 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 13.200 16.670 13.520 ;
      LAYER met4 ;
        RECT 16.350 13.200 16.670 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 12.770 16.670 13.090 ;
      LAYER met4 ;
        RECT 16.350 12.770 16.670 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 12.340 16.670 12.660 ;
      LAYER met4 ;
        RECT 16.350 12.340 16.670 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 11.910 16.670 12.230 ;
      LAYER met4 ;
        RECT 16.350 11.910 16.670 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 11.480 16.670 11.800 ;
      LAYER met4 ;
        RECT 16.350 11.480 16.670 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 11.050 16.670 11.370 ;
      LAYER met4 ;
        RECT 16.350 11.050 16.670 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 10.620 16.670 10.940 ;
      LAYER met4 ;
        RECT 16.350 10.620 16.670 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 10.190 16.670 10.510 ;
      LAYER met4 ;
        RECT 16.350 10.190 16.670 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 9.760 16.670 10.080 ;
      LAYER met4 ;
        RECT 16.350 9.760 16.670 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 9.330 16.670 9.650 ;
      LAYER met4 ;
        RECT 16.350 9.330 16.670 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 8.900 16.670 9.220 ;
      LAYER met4 ;
        RECT 16.350 8.900 16.670 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 13.200 16.265 13.520 ;
      LAYER met4 ;
        RECT 15.945 13.200 16.265 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 12.770 16.265 13.090 ;
      LAYER met4 ;
        RECT 15.945 12.770 16.265 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 12.340 16.265 12.660 ;
      LAYER met4 ;
        RECT 15.945 12.340 16.265 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 11.910 16.265 12.230 ;
      LAYER met4 ;
        RECT 15.945 11.910 16.265 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 11.480 16.265 11.800 ;
      LAYER met4 ;
        RECT 15.945 11.480 16.265 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 11.050 16.265 11.370 ;
      LAYER met4 ;
        RECT 15.945 11.050 16.265 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 10.620 16.265 10.940 ;
      LAYER met4 ;
        RECT 15.945 10.620 16.265 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 10.190 16.265 10.510 ;
      LAYER met4 ;
        RECT 15.945 10.190 16.265 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 9.760 16.265 10.080 ;
      LAYER met4 ;
        RECT 15.945 9.760 16.265 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 9.330 16.265 9.650 ;
      LAYER met4 ;
        RECT 15.945 9.330 16.265 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 8.900 16.265 9.220 ;
      LAYER met4 ;
        RECT 15.945 8.900 16.265 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 13.200 15.860 13.520 ;
      LAYER met4 ;
        RECT 15.540 13.200 15.860 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 12.770 15.860 13.090 ;
      LAYER met4 ;
        RECT 15.540 12.770 15.860 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 12.340 15.860 12.660 ;
      LAYER met4 ;
        RECT 15.540 12.340 15.860 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 11.910 15.860 12.230 ;
      LAYER met4 ;
        RECT 15.540 11.910 15.860 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 11.480 15.860 11.800 ;
      LAYER met4 ;
        RECT 15.540 11.480 15.860 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 11.050 15.860 11.370 ;
      LAYER met4 ;
        RECT 15.540 11.050 15.860 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 10.620 15.860 10.940 ;
      LAYER met4 ;
        RECT 15.540 10.620 15.860 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 10.190 15.860 10.510 ;
      LAYER met4 ;
        RECT 15.540 10.190 15.860 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 9.760 15.860 10.080 ;
      LAYER met4 ;
        RECT 15.540 9.760 15.860 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 9.330 15.860 9.650 ;
      LAYER met4 ;
        RECT 15.540 9.330 15.860 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 8.900 15.860 9.220 ;
      LAYER met4 ;
        RECT 15.540 8.900 15.860 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 13.200 15.455 13.520 ;
      LAYER met4 ;
        RECT 15.135 13.200 15.455 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 12.770 15.455 13.090 ;
      LAYER met4 ;
        RECT 15.135 12.770 15.455 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 12.340 15.455 12.660 ;
      LAYER met4 ;
        RECT 15.135 12.340 15.455 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 11.910 15.455 12.230 ;
      LAYER met4 ;
        RECT 15.135 11.910 15.455 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 11.480 15.455 11.800 ;
      LAYER met4 ;
        RECT 15.135 11.480 15.455 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 11.050 15.455 11.370 ;
      LAYER met4 ;
        RECT 15.135 11.050 15.455 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 10.620 15.455 10.940 ;
      LAYER met4 ;
        RECT 15.135 10.620 15.455 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 10.190 15.455 10.510 ;
      LAYER met4 ;
        RECT 15.135 10.190 15.455 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 9.760 15.455 10.080 ;
      LAYER met4 ;
        RECT 15.135 9.760 15.455 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 9.330 15.455 9.650 ;
      LAYER met4 ;
        RECT 15.135 9.330 15.455 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 8.900 15.455 9.220 ;
      LAYER met4 ;
        RECT 15.135 8.900 15.455 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 13.200 15.050 13.520 ;
      LAYER met4 ;
        RECT 14.730 13.200 15.050 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 12.770 15.050 13.090 ;
      LAYER met4 ;
        RECT 14.730 12.770 15.050 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 12.340 15.050 12.660 ;
      LAYER met4 ;
        RECT 14.730 12.340 15.050 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 11.910 15.050 12.230 ;
      LAYER met4 ;
        RECT 14.730 11.910 15.050 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 11.480 15.050 11.800 ;
      LAYER met4 ;
        RECT 14.730 11.480 15.050 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 11.050 15.050 11.370 ;
      LAYER met4 ;
        RECT 14.730 11.050 15.050 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 10.620 15.050 10.940 ;
      LAYER met4 ;
        RECT 14.730 10.620 15.050 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 10.190 15.050 10.510 ;
      LAYER met4 ;
        RECT 14.730 10.190 15.050 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 9.760 15.050 10.080 ;
      LAYER met4 ;
        RECT 14.730 9.760 15.050 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 9.330 15.050 9.650 ;
      LAYER met4 ;
        RECT 14.730 9.330 15.050 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 8.900 15.050 9.220 ;
      LAYER met4 ;
        RECT 14.730 8.900 15.050 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 13.200 14.645 13.520 ;
      LAYER met4 ;
        RECT 14.325 13.200 14.645 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 12.770 14.645 13.090 ;
      LAYER met4 ;
        RECT 14.325 12.770 14.645 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 12.340 14.645 12.660 ;
      LAYER met4 ;
        RECT 14.325 12.340 14.645 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 11.910 14.645 12.230 ;
      LAYER met4 ;
        RECT 14.325 11.910 14.645 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 11.480 14.645 11.800 ;
      LAYER met4 ;
        RECT 14.325 11.480 14.645 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 11.050 14.645 11.370 ;
      LAYER met4 ;
        RECT 14.325 11.050 14.645 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 10.620 14.645 10.940 ;
      LAYER met4 ;
        RECT 14.325 10.620 14.645 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 10.190 14.645 10.510 ;
      LAYER met4 ;
        RECT 14.325 10.190 14.645 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 9.760 14.645 10.080 ;
      LAYER met4 ;
        RECT 14.325 9.760 14.645 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 9.330 14.645 9.650 ;
      LAYER met4 ;
        RECT 14.325 9.330 14.645 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 8.900 14.645 9.220 ;
      LAYER met4 ;
        RECT 14.325 8.900 14.645 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 13.200 14.240 13.520 ;
      LAYER met4 ;
        RECT 13.920 13.200 14.240 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 12.770 14.240 13.090 ;
      LAYER met4 ;
        RECT 13.920 12.770 14.240 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 12.340 14.240 12.660 ;
      LAYER met4 ;
        RECT 13.920 12.340 14.240 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 11.910 14.240 12.230 ;
      LAYER met4 ;
        RECT 13.920 11.910 14.240 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 11.480 14.240 11.800 ;
      LAYER met4 ;
        RECT 13.920 11.480 14.240 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 11.050 14.240 11.370 ;
      LAYER met4 ;
        RECT 13.920 11.050 14.240 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 10.620 14.240 10.940 ;
      LAYER met4 ;
        RECT 13.920 10.620 14.240 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 10.190 14.240 10.510 ;
      LAYER met4 ;
        RECT 13.920 10.190 14.240 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 9.760 14.240 10.080 ;
      LAYER met4 ;
        RECT 13.920 9.760 14.240 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 9.330 14.240 9.650 ;
      LAYER met4 ;
        RECT 13.920 9.330 14.240 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 8.900 14.240 9.220 ;
      LAYER met4 ;
        RECT 13.920 8.900 14.240 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 13.200 13.835 13.520 ;
      LAYER met4 ;
        RECT 13.515 13.200 13.835 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 12.770 13.835 13.090 ;
      LAYER met4 ;
        RECT 13.515 12.770 13.835 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 12.340 13.835 12.660 ;
      LAYER met4 ;
        RECT 13.515 12.340 13.835 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 11.910 13.835 12.230 ;
      LAYER met4 ;
        RECT 13.515 11.910 13.835 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 11.480 13.835 11.800 ;
      LAYER met4 ;
        RECT 13.515 11.480 13.835 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 11.050 13.835 11.370 ;
      LAYER met4 ;
        RECT 13.515 11.050 13.835 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 10.620 13.835 10.940 ;
      LAYER met4 ;
        RECT 13.515 10.620 13.835 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 10.190 13.835 10.510 ;
      LAYER met4 ;
        RECT 13.515 10.190 13.835 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 9.760 13.835 10.080 ;
      LAYER met4 ;
        RECT 13.515 9.760 13.835 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 9.330 13.835 9.650 ;
      LAYER met4 ;
        RECT 13.515 9.330 13.835 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 8.900 13.835 9.220 ;
      LAYER met4 ;
        RECT 13.515 8.900 13.835 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 13.200 13.430 13.520 ;
      LAYER met4 ;
        RECT 13.110 13.200 13.430 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 12.770 13.430 13.090 ;
      LAYER met4 ;
        RECT 13.110 12.770 13.430 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 12.340 13.430 12.660 ;
      LAYER met4 ;
        RECT 13.110 12.340 13.430 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 11.910 13.430 12.230 ;
      LAYER met4 ;
        RECT 13.110 11.910 13.430 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 11.480 13.430 11.800 ;
      LAYER met4 ;
        RECT 13.110 11.480 13.430 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 11.050 13.430 11.370 ;
      LAYER met4 ;
        RECT 13.110 11.050 13.430 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 10.620 13.430 10.940 ;
      LAYER met4 ;
        RECT 13.110 10.620 13.430 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 10.190 13.430 10.510 ;
      LAYER met4 ;
        RECT 13.110 10.190 13.430 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 9.760 13.430 10.080 ;
      LAYER met4 ;
        RECT 13.110 9.760 13.430 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 9.330 13.430 9.650 ;
      LAYER met4 ;
        RECT 13.110 9.330 13.430 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 8.900 13.430 9.220 ;
      LAYER met4 ;
        RECT 13.110 8.900 13.430 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 13.200 13.025 13.520 ;
      LAYER met4 ;
        RECT 12.705 13.200 13.025 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 12.770 13.025 13.090 ;
      LAYER met4 ;
        RECT 12.705 12.770 13.025 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 12.340 13.025 12.660 ;
      LAYER met4 ;
        RECT 12.705 12.340 13.025 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 11.910 13.025 12.230 ;
      LAYER met4 ;
        RECT 12.705 11.910 13.025 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 11.480 13.025 11.800 ;
      LAYER met4 ;
        RECT 12.705 11.480 13.025 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 11.050 13.025 11.370 ;
      LAYER met4 ;
        RECT 12.705 11.050 13.025 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 10.620 13.025 10.940 ;
      LAYER met4 ;
        RECT 12.705 10.620 13.025 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 10.190 13.025 10.510 ;
      LAYER met4 ;
        RECT 12.705 10.190 13.025 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 9.760 13.025 10.080 ;
      LAYER met4 ;
        RECT 12.705 9.760 13.025 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 9.330 13.025 9.650 ;
      LAYER met4 ;
        RECT 12.705 9.330 13.025 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 8.900 13.025 9.220 ;
      LAYER met4 ;
        RECT 12.705 8.900 13.025 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 13.200 12.620 13.520 ;
      LAYER met4 ;
        RECT 12.300 13.200 12.620 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 12.770 12.620 13.090 ;
      LAYER met4 ;
        RECT 12.300 12.770 12.620 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 12.340 12.620 12.660 ;
      LAYER met4 ;
        RECT 12.300 12.340 12.620 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 11.910 12.620 12.230 ;
      LAYER met4 ;
        RECT 12.300 11.910 12.620 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 11.480 12.620 11.800 ;
      LAYER met4 ;
        RECT 12.300 11.480 12.620 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 11.050 12.620 11.370 ;
      LAYER met4 ;
        RECT 12.300 11.050 12.620 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 10.620 12.620 10.940 ;
      LAYER met4 ;
        RECT 12.300 10.620 12.620 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 10.190 12.620 10.510 ;
      LAYER met4 ;
        RECT 12.300 10.190 12.620 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 9.760 12.620 10.080 ;
      LAYER met4 ;
        RECT 12.300 9.760 12.620 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 9.330 12.620 9.650 ;
      LAYER met4 ;
        RECT 12.300 9.330 12.620 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 8.900 12.620 9.220 ;
      LAYER met4 ;
        RECT 12.300 8.900 12.620 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 13.200 12.215 13.520 ;
      LAYER met4 ;
        RECT 11.895 13.200 12.215 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 12.770 12.215 13.090 ;
      LAYER met4 ;
        RECT 11.895 12.770 12.215 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 12.340 12.215 12.660 ;
      LAYER met4 ;
        RECT 11.895 12.340 12.215 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 11.910 12.215 12.230 ;
      LAYER met4 ;
        RECT 11.895 11.910 12.215 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 11.480 12.215 11.800 ;
      LAYER met4 ;
        RECT 11.895 11.480 12.215 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 11.050 12.215 11.370 ;
      LAYER met4 ;
        RECT 11.895 11.050 12.215 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 10.620 12.215 10.940 ;
      LAYER met4 ;
        RECT 11.895 10.620 12.215 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 10.190 12.215 10.510 ;
      LAYER met4 ;
        RECT 11.895 10.190 12.215 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 9.760 12.215 10.080 ;
      LAYER met4 ;
        RECT 11.895 9.760 12.215 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 9.330 12.215 9.650 ;
      LAYER met4 ;
        RECT 11.895 9.330 12.215 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 8.900 12.215 9.220 ;
      LAYER met4 ;
        RECT 11.895 8.900 12.215 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 13.200 11.810 13.520 ;
      LAYER met4 ;
        RECT 11.490 13.200 11.810 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 12.770 11.810 13.090 ;
      LAYER met4 ;
        RECT 11.490 12.770 11.810 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 12.340 11.810 12.660 ;
      LAYER met4 ;
        RECT 11.490 12.340 11.810 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 11.910 11.810 12.230 ;
      LAYER met4 ;
        RECT 11.490 11.910 11.810 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 11.480 11.810 11.800 ;
      LAYER met4 ;
        RECT 11.490 11.480 11.810 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 11.050 11.810 11.370 ;
      LAYER met4 ;
        RECT 11.490 11.050 11.810 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 10.620 11.810 10.940 ;
      LAYER met4 ;
        RECT 11.490 10.620 11.810 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 10.190 11.810 10.510 ;
      LAYER met4 ;
        RECT 11.490 10.190 11.810 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 9.760 11.810 10.080 ;
      LAYER met4 ;
        RECT 11.490 9.760 11.810 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 9.330 11.810 9.650 ;
      LAYER met4 ;
        RECT 11.490 9.330 11.810 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 8.900 11.810 9.220 ;
      LAYER met4 ;
        RECT 11.490 8.900 11.810 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 13.200 11.405 13.520 ;
      LAYER met4 ;
        RECT 11.085 13.200 11.405 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 12.770 11.405 13.090 ;
      LAYER met4 ;
        RECT 11.085 12.770 11.405 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 12.340 11.405 12.660 ;
      LAYER met4 ;
        RECT 11.085 12.340 11.405 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 11.910 11.405 12.230 ;
      LAYER met4 ;
        RECT 11.085 11.910 11.405 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 11.480 11.405 11.800 ;
      LAYER met4 ;
        RECT 11.085 11.480 11.405 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 11.050 11.405 11.370 ;
      LAYER met4 ;
        RECT 11.085 11.050 11.405 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 10.620 11.405 10.940 ;
      LAYER met4 ;
        RECT 11.085 10.620 11.405 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 10.190 11.405 10.510 ;
      LAYER met4 ;
        RECT 11.085 10.190 11.405 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 9.760 11.405 10.080 ;
      LAYER met4 ;
        RECT 11.085 9.760 11.405 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 9.330 11.405 9.650 ;
      LAYER met4 ;
        RECT 11.085 9.330 11.405 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 8.900 11.405 9.220 ;
      LAYER met4 ;
        RECT 11.085 8.900 11.405 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 13.200 11.000 13.520 ;
      LAYER met4 ;
        RECT 10.680 13.200 11.000 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 12.770 11.000 13.090 ;
      LAYER met4 ;
        RECT 10.680 12.770 11.000 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 12.340 11.000 12.660 ;
      LAYER met4 ;
        RECT 10.680 12.340 11.000 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 11.910 11.000 12.230 ;
      LAYER met4 ;
        RECT 10.680 11.910 11.000 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 11.480 11.000 11.800 ;
      LAYER met4 ;
        RECT 10.680 11.480 11.000 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 11.050 11.000 11.370 ;
      LAYER met4 ;
        RECT 10.680 11.050 11.000 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 10.620 11.000 10.940 ;
      LAYER met4 ;
        RECT 10.680 10.620 11.000 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 10.190 11.000 10.510 ;
      LAYER met4 ;
        RECT 10.680 10.190 11.000 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 9.760 11.000 10.080 ;
      LAYER met4 ;
        RECT 10.680 9.760 11.000 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 9.330 11.000 9.650 ;
      LAYER met4 ;
        RECT 10.680 9.330 11.000 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 8.900 11.000 9.220 ;
      LAYER met4 ;
        RECT 10.680 8.900 11.000 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 13.200 10.595 13.520 ;
      LAYER met4 ;
        RECT 10.275 13.200 10.595 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 12.770 10.595 13.090 ;
      LAYER met4 ;
        RECT 10.275 12.770 10.595 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 12.340 10.595 12.660 ;
      LAYER met4 ;
        RECT 10.275 12.340 10.595 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 11.910 10.595 12.230 ;
      LAYER met4 ;
        RECT 10.275 11.910 10.595 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 11.480 10.595 11.800 ;
      LAYER met4 ;
        RECT 10.275 11.480 10.595 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 11.050 10.595 11.370 ;
      LAYER met4 ;
        RECT 10.275 11.050 10.595 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 10.620 10.595 10.940 ;
      LAYER met4 ;
        RECT 10.275 10.620 10.595 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 10.190 10.595 10.510 ;
      LAYER met4 ;
        RECT 10.275 10.190 10.595 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 9.760 10.595 10.080 ;
      LAYER met4 ;
        RECT 10.275 9.760 10.595 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 9.330 10.595 9.650 ;
      LAYER met4 ;
        RECT 10.275 9.330 10.595 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 8.900 10.595 9.220 ;
      LAYER met4 ;
        RECT 10.275 8.900 10.595 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 13.200 10.190 13.520 ;
      LAYER met4 ;
        RECT 9.870 13.200 10.190 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 12.770 10.190 13.090 ;
      LAYER met4 ;
        RECT 9.870 12.770 10.190 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 12.340 10.190 12.660 ;
      LAYER met4 ;
        RECT 9.870 12.340 10.190 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 11.910 10.190 12.230 ;
      LAYER met4 ;
        RECT 9.870 11.910 10.190 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 11.480 10.190 11.800 ;
      LAYER met4 ;
        RECT 9.870 11.480 10.190 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 11.050 10.190 11.370 ;
      LAYER met4 ;
        RECT 9.870 11.050 10.190 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 10.620 10.190 10.940 ;
      LAYER met4 ;
        RECT 9.870 10.620 10.190 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 10.190 10.190 10.510 ;
      LAYER met4 ;
        RECT 9.870 10.190 10.190 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 9.760 10.190 10.080 ;
      LAYER met4 ;
        RECT 9.870 9.760 10.190 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 9.330 10.190 9.650 ;
      LAYER met4 ;
        RECT 9.870 9.330 10.190 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 8.900 10.190 9.220 ;
      LAYER met4 ;
        RECT 9.870 8.900 10.190 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 13.200 9.785 13.520 ;
      LAYER met4 ;
        RECT 9.465 13.200 9.785 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 12.770 9.785 13.090 ;
      LAYER met4 ;
        RECT 9.465 12.770 9.785 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 12.340 9.785 12.660 ;
      LAYER met4 ;
        RECT 9.465 12.340 9.785 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 11.910 9.785 12.230 ;
      LAYER met4 ;
        RECT 9.465 11.910 9.785 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 11.480 9.785 11.800 ;
      LAYER met4 ;
        RECT 9.465 11.480 9.785 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 11.050 9.785 11.370 ;
      LAYER met4 ;
        RECT 9.465 11.050 9.785 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 10.620 9.785 10.940 ;
      LAYER met4 ;
        RECT 9.465 10.620 9.785 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 10.190 9.785 10.510 ;
      LAYER met4 ;
        RECT 9.465 10.190 9.785 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 9.760 9.785 10.080 ;
      LAYER met4 ;
        RECT 9.465 9.760 9.785 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 9.330 9.785 9.650 ;
      LAYER met4 ;
        RECT 9.465 9.330 9.785 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 8.900 9.785 9.220 ;
      LAYER met4 ;
        RECT 9.465 8.900 9.785 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 13.200 9.380 13.520 ;
      LAYER met4 ;
        RECT 9.060 13.200 9.380 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 12.770 9.380 13.090 ;
      LAYER met4 ;
        RECT 9.060 12.770 9.380 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 12.340 9.380 12.660 ;
      LAYER met4 ;
        RECT 9.060 12.340 9.380 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 11.910 9.380 12.230 ;
      LAYER met4 ;
        RECT 9.060 11.910 9.380 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 11.480 9.380 11.800 ;
      LAYER met4 ;
        RECT 9.060 11.480 9.380 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 11.050 9.380 11.370 ;
      LAYER met4 ;
        RECT 9.060 11.050 9.380 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 10.620 9.380 10.940 ;
      LAYER met4 ;
        RECT 9.060 10.620 9.380 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 10.190 9.380 10.510 ;
      LAYER met4 ;
        RECT 9.060 10.190 9.380 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 9.760 9.380 10.080 ;
      LAYER met4 ;
        RECT 9.060 9.760 9.380 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 9.330 9.380 9.650 ;
      LAYER met4 ;
        RECT 9.060 9.330 9.380 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 8.900 9.380 9.220 ;
      LAYER met4 ;
        RECT 9.060 8.900 9.380 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 13.200 8.975 13.520 ;
      LAYER met4 ;
        RECT 8.655 13.200 8.975 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 12.770 8.975 13.090 ;
      LAYER met4 ;
        RECT 8.655 12.770 8.975 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 12.340 8.975 12.660 ;
      LAYER met4 ;
        RECT 8.655 12.340 8.975 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 11.910 8.975 12.230 ;
      LAYER met4 ;
        RECT 8.655 11.910 8.975 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 11.480 8.975 11.800 ;
      LAYER met4 ;
        RECT 8.655 11.480 8.975 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 11.050 8.975 11.370 ;
      LAYER met4 ;
        RECT 8.655 11.050 8.975 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 10.620 8.975 10.940 ;
      LAYER met4 ;
        RECT 8.655 10.620 8.975 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 10.190 8.975 10.510 ;
      LAYER met4 ;
        RECT 8.655 10.190 8.975 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 9.760 8.975 10.080 ;
      LAYER met4 ;
        RECT 8.655 9.760 8.975 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 9.330 8.975 9.650 ;
      LAYER met4 ;
        RECT 8.655 9.330 8.975 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 8.900 8.975 9.220 ;
      LAYER met4 ;
        RECT 8.655 8.900 8.975 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 13.200 8.570 13.520 ;
      LAYER met4 ;
        RECT 8.250 13.200 8.570 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 12.770 8.570 13.090 ;
      LAYER met4 ;
        RECT 8.250 12.770 8.570 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 12.340 8.570 12.660 ;
      LAYER met4 ;
        RECT 8.250 12.340 8.570 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 11.910 8.570 12.230 ;
      LAYER met4 ;
        RECT 8.250 11.910 8.570 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 11.480 8.570 11.800 ;
      LAYER met4 ;
        RECT 8.250 11.480 8.570 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 11.050 8.570 11.370 ;
      LAYER met4 ;
        RECT 8.250 11.050 8.570 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 10.620 8.570 10.940 ;
      LAYER met4 ;
        RECT 8.250 10.620 8.570 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 10.190 8.570 10.510 ;
      LAYER met4 ;
        RECT 8.250 10.190 8.570 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 9.760 8.570 10.080 ;
      LAYER met4 ;
        RECT 8.250 9.760 8.570 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 9.330 8.570 9.650 ;
      LAYER met4 ;
        RECT 8.250 9.330 8.570 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 8.900 8.570 9.220 ;
      LAYER met4 ;
        RECT 8.250 8.900 8.570 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 13.200 8.165 13.520 ;
      LAYER met4 ;
        RECT 7.845 13.200 8.165 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 12.770 8.165 13.090 ;
      LAYER met4 ;
        RECT 7.845 12.770 8.165 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 12.340 8.165 12.660 ;
      LAYER met4 ;
        RECT 7.845 12.340 8.165 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 11.910 8.165 12.230 ;
      LAYER met4 ;
        RECT 7.845 11.910 8.165 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 11.480 8.165 11.800 ;
      LAYER met4 ;
        RECT 7.845 11.480 8.165 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 11.050 8.165 11.370 ;
      LAYER met4 ;
        RECT 7.845 11.050 8.165 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 10.620 8.165 10.940 ;
      LAYER met4 ;
        RECT 7.845 10.620 8.165 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 10.190 8.165 10.510 ;
      LAYER met4 ;
        RECT 7.845 10.190 8.165 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 9.760 8.165 10.080 ;
      LAYER met4 ;
        RECT 7.845 9.760 8.165 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 9.330 8.165 9.650 ;
      LAYER met4 ;
        RECT 7.845 9.330 8.165 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 8.900 8.165 9.220 ;
      LAYER met4 ;
        RECT 7.845 8.900 8.165 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 13.200 7.760 13.520 ;
      LAYER met4 ;
        RECT 7.440 13.200 7.760 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 12.770 7.760 13.090 ;
      LAYER met4 ;
        RECT 7.440 12.770 7.760 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 12.340 7.760 12.660 ;
      LAYER met4 ;
        RECT 7.440 12.340 7.760 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 11.910 7.760 12.230 ;
      LAYER met4 ;
        RECT 7.440 11.910 7.760 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 11.480 7.760 11.800 ;
      LAYER met4 ;
        RECT 7.440 11.480 7.760 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 11.050 7.760 11.370 ;
      LAYER met4 ;
        RECT 7.440 11.050 7.760 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 10.620 7.760 10.940 ;
      LAYER met4 ;
        RECT 7.440 10.620 7.760 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 10.190 7.760 10.510 ;
      LAYER met4 ;
        RECT 7.440 10.190 7.760 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 9.760 7.760 10.080 ;
      LAYER met4 ;
        RECT 7.440 9.760 7.760 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 9.330 7.760 9.650 ;
      LAYER met4 ;
        RECT 7.440 9.330 7.760 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 8.900 7.760 9.220 ;
      LAYER met4 ;
        RECT 7.440 8.900 7.760 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 13.200 7.355 13.520 ;
      LAYER met4 ;
        RECT 7.035 13.200 7.355 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 12.770 7.355 13.090 ;
      LAYER met4 ;
        RECT 7.035 12.770 7.355 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 12.340 7.355 12.660 ;
      LAYER met4 ;
        RECT 7.035 12.340 7.355 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 11.910 7.355 12.230 ;
      LAYER met4 ;
        RECT 7.035 11.910 7.355 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 11.480 7.355 11.800 ;
      LAYER met4 ;
        RECT 7.035 11.480 7.355 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 11.050 7.355 11.370 ;
      LAYER met4 ;
        RECT 7.035 11.050 7.355 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 10.620 7.355 10.940 ;
      LAYER met4 ;
        RECT 7.035 10.620 7.355 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 10.190 7.355 10.510 ;
      LAYER met4 ;
        RECT 7.035 10.190 7.355 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 9.760 7.355 10.080 ;
      LAYER met4 ;
        RECT 7.035 9.760 7.355 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 9.330 7.355 9.650 ;
      LAYER met4 ;
        RECT 7.035 9.330 7.355 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 8.900 7.355 9.220 ;
      LAYER met4 ;
        RECT 7.035 8.900 7.355 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 13.200 6.950 13.520 ;
      LAYER met4 ;
        RECT 6.630 13.200 6.950 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 12.770 6.950 13.090 ;
      LAYER met4 ;
        RECT 6.630 12.770 6.950 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 12.340 6.950 12.660 ;
      LAYER met4 ;
        RECT 6.630 12.340 6.950 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 11.910 6.950 12.230 ;
      LAYER met4 ;
        RECT 6.630 11.910 6.950 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 11.480 6.950 11.800 ;
      LAYER met4 ;
        RECT 6.630 11.480 6.950 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 11.050 6.950 11.370 ;
      LAYER met4 ;
        RECT 6.630 11.050 6.950 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 10.620 6.950 10.940 ;
      LAYER met4 ;
        RECT 6.630 10.620 6.950 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 10.190 6.950 10.510 ;
      LAYER met4 ;
        RECT 6.630 10.190 6.950 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 9.760 6.950 10.080 ;
      LAYER met4 ;
        RECT 6.630 9.760 6.950 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 9.330 6.950 9.650 ;
      LAYER met4 ;
        RECT 6.630 9.330 6.950 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 8.900 6.950 9.220 ;
      LAYER met4 ;
        RECT 6.630 8.900 6.950 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 13.200 6.545 13.520 ;
      LAYER met4 ;
        RECT 6.225 13.200 6.545 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 12.770 6.545 13.090 ;
      LAYER met4 ;
        RECT 6.225 12.770 6.545 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 12.340 6.545 12.660 ;
      LAYER met4 ;
        RECT 6.225 12.340 6.545 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 11.910 6.545 12.230 ;
      LAYER met4 ;
        RECT 6.225 11.910 6.545 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 11.480 6.545 11.800 ;
      LAYER met4 ;
        RECT 6.225 11.480 6.545 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 11.050 6.545 11.370 ;
      LAYER met4 ;
        RECT 6.225 11.050 6.545 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 10.620 6.545 10.940 ;
      LAYER met4 ;
        RECT 6.225 10.620 6.545 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 10.190 6.545 10.510 ;
      LAYER met4 ;
        RECT 6.225 10.190 6.545 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 9.760 6.545 10.080 ;
      LAYER met4 ;
        RECT 6.225 9.760 6.545 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 9.330 6.545 9.650 ;
      LAYER met4 ;
        RECT 6.225 9.330 6.545 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 8.900 6.545 9.220 ;
      LAYER met4 ;
        RECT 6.225 8.900 6.545 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 13.200 6.140 13.520 ;
      LAYER met4 ;
        RECT 5.820 13.200 6.140 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 12.770 6.140 13.090 ;
      LAYER met4 ;
        RECT 5.820 12.770 6.140 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 12.340 6.140 12.660 ;
      LAYER met4 ;
        RECT 5.820 12.340 6.140 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 11.910 6.140 12.230 ;
      LAYER met4 ;
        RECT 5.820 11.910 6.140 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 11.480 6.140 11.800 ;
      LAYER met4 ;
        RECT 5.820 11.480 6.140 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 11.050 6.140 11.370 ;
      LAYER met4 ;
        RECT 5.820 11.050 6.140 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 10.620 6.140 10.940 ;
      LAYER met4 ;
        RECT 5.820 10.620 6.140 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 10.190 6.140 10.510 ;
      LAYER met4 ;
        RECT 5.820 10.190 6.140 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 9.760 6.140 10.080 ;
      LAYER met4 ;
        RECT 5.820 9.760 6.140 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 9.330 6.140 9.650 ;
      LAYER met4 ;
        RECT 5.820 9.330 6.140 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 8.900 6.140 9.220 ;
      LAYER met4 ;
        RECT 5.820 8.900 6.140 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 13.200 5.735 13.520 ;
      LAYER met4 ;
        RECT 5.415 13.200 5.735 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 12.770 5.735 13.090 ;
      LAYER met4 ;
        RECT 5.415 12.770 5.735 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 12.340 5.735 12.660 ;
      LAYER met4 ;
        RECT 5.415 12.340 5.735 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 11.910 5.735 12.230 ;
      LAYER met4 ;
        RECT 5.415 11.910 5.735 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 11.480 5.735 11.800 ;
      LAYER met4 ;
        RECT 5.415 11.480 5.735 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 11.050 5.735 11.370 ;
      LAYER met4 ;
        RECT 5.415 11.050 5.735 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 10.620 5.735 10.940 ;
      LAYER met4 ;
        RECT 5.415 10.620 5.735 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 10.190 5.735 10.510 ;
      LAYER met4 ;
        RECT 5.415 10.190 5.735 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 9.760 5.735 10.080 ;
      LAYER met4 ;
        RECT 5.415 9.760 5.735 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 9.330 5.735 9.650 ;
      LAYER met4 ;
        RECT 5.415 9.330 5.735 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 8.900 5.735 9.220 ;
      LAYER met4 ;
        RECT 5.415 8.900 5.735 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 13.200 5.330 13.520 ;
      LAYER met4 ;
        RECT 5.010 13.200 5.330 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 12.770 5.330 13.090 ;
      LAYER met4 ;
        RECT 5.010 12.770 5.330 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 12.340 5.330 12.660 ;
      LAYER met4 ;
        RECT 5.010 12.340 5.330 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 11.910 5.330 12.230 ;
      LAYER met4 ;
        RECT 5.010 11.910 5.330 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 11.480 5.330 11.800 ;
      LAYER met4 ;
        RECT 5.010 11.480 5.330 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 11.050 5.330 11.370 ;
      LAYER met4 ;
        RECT 5.010 11.050 5.330 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 10.620 5.330 10.940 ;
      LAYER met4 ;
        RECT 5.010 10.620 5.330 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 10.190 5.330 10.510 ;
      LAYER met4 ;
        RECT 5.010 10.190 5.330 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 9.760 5.330 10.080 ;
      LAYER met4 ;
        RECT 5.010 9.760 5.330 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 9.330 5.330 9.650 ;
      LAYER met4 ;
        RECT 5.010 9.330 5.330 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 8.900 5.330 9.220 ;
      LAYER met4 ;
        RECT 5.010 8.900 5.330 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 13.200 4.925 13.520 ;
      LAYER met4 ;
        RECT 4.605 13.200 4.925 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 12.770 4.925 13.090 ;
      LAYER met4 ;
        RECT 4.605 12.770 4.925 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 12.340 4.925 12.660 ;
      LAYER met4 ;
        RECT 4.605 12.340 4.925 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 11.910 4.925 12.230 ;
      LAYER met4 ;
        RECT 4.605 11.910 4.925 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 11.480 4.925 11.800 ;
      LAYER met4 ;
        RECT 4.605 11.480 4.925 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 11.050 4.925 11.370 ;
      LAYER met4 ;
        RECT 4.605 11.050 4.925 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 10.620 4.925 10.940 ;
      LAYER met4 ;
        RECT 4.605 10.620 4.925 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 10.190 4.925 10.510 ;
      LAYER met4 ;
        RECT 4.605 10.190 4.925 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 9.760 4.925 10.080 ;
      LAYER met4 ;
        RECT 4.605 9.760 4.925 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 9.330 4.925 9.650 ;
      LAYER met4 ;
        RECT 4.605 9.330 4.925 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 8.900 4.925 9.220 ;
      LAYER met4 ;
        RECT 4.605 8.900 4.925 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 13.200 4.520 13.520 ;
      LAYER met4 ;
        RECT 4.200 13.200 4.520 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 12.770 4.520 13.090 ;
      LAYER met4 ;
        RECT 4.200 12.770 4.520 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 12.340 4.520 12.660 ;
      LAYER met4 ;
        RECT 4.200 12.340 4.520 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 11.910 4.520 12.230 ;
      LAYER met4 ;
        RECT 4.200 11.910 4.520 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 11.480 4.520 11.800 ;
      LAYER met4 ;
        RECT 4.200 11.480 4.520 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 11.050 4.520 11.370 ;
      LAYER met4 ;
        RECT 4.200 11.050 4.520 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 10.620 4.520 10.940 ;
      LAYER met4 ;
        RECT 4.200 10.620 4.520 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 10.190 4.520 10.510 ;
      LAYER met4 ;
        RECT 4.200 10.190 4.520 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 9.760 4.520 10.080 ;
      LAYER met4 ;
        RECT 4.200 9.760 4.520 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 9.330 4.520 9.650 ;
      LAYER met4 ;
        RECT 4.200 9.330 4.520 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 8.900 4.520 9.220 ;
      LAYER met4 ;
        RECT 4.200 8.900 4.520 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 13.200 4.115 13.520 ;
      LAYER met4 ;
        RECT 3.795 13.200 4.115 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 12.770 4.115 13.090 ;
      LAYER met4 ;
        RECT 3.795 12.770 4.115 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 12.340 4.115 12.660 ;
      LAYER met4 ;
        RECT 3.795 12.340 4.115 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 11.910 4.115 12.230 ;
      LAYER met4 ;
        RECT 3.795 11.910 4.115 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 11.480 4.115 11.800 ;
      LAYER met4 ;
        RECT 3.795 11.480 4.115 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 11.050 4.115 11.370 ;
      LAYER met4 ;
        RECT 3.795 11.050 4.115 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 10.620 4.115 10.940 ;
      LAYER met4 ;
        RECT 3.795 10.620 4.115 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 10.190 4.115 10.510 ;
      LAYER met4 ;
        RECT 3.795 10.190 4.115 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 9.760 4.115 10.080 ;
      LAYER met4 ;
        RECT 3.795 9.760 4.115 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 9.330 4.115 9.650 ;
      LAYER met4 ;
        RECT 3.795 9.330 4.115 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 8.900 4.115 9.220 ;
      LAYER met4 ;
        RECT 3.795 8.900 4.115 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 13.200 3.710 13.520 ;
      LAYER met4 ;
        RECT 3.390 13.200 3.710 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 12.770 3.710 13.090 ;
      LAYER met4 ;
        RECT 3.390 12.770 3.710 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 12.340 3.710 12.660 ;
      LAYER met4 ;
        RECT 3.390 12.340 3.710 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 11.910 3.710 12.230 ;
      LAYER met4 ;
        RECT 3.390 11.910 3.710 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 11.480 3.710 11.800 ;
      LAYER met4 ;
        RECT 3.390 11.480 3.710 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 11.050 3.710 11.370 ;
      LAYER met4 ;
        RECT 3.390 11.050 3.710 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 10.620 3.710 10.940 ;
      LAYER met4 ;
        RECT 3.390 10.620 3.710 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 10.190 3.710 10.510 ;
      LAYER met4 ;
        RECT 3.390 10.190 3.710 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 9.760 3.710 10.080 ;
      LAYER met4 ;
        RECT 3.390 9.760 3.710 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 9.330 3.710 9.650 ;
      LAYER met4 ;
        RECT 3.390 9.330 3.710 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 8.900 3.710 9.220 ;
      LAYER met4 ;
        RECT 3.390 8.900 3.710 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 13.200 3.305 13.520 ;
      LAYER met4 ;
        RECT 2.985 13.200 3.305 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 12.770 3.305 13.090 ;
      LAYER met4 ;
        RECT 2.985 12.770 3.305 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 12.340 3.305 12.660 ;
      LAYER met4 ;
        RECT 2.985 12.340 3.305 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 11.910 3.305 12.230 ;
      LAYER met4 ;
        RECT 2.985 11.910 3.305 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 11.480 3.305 11.800 ;
      LAYER met4 ;
        RECT 2.985 11.480 3.305 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 11.050 3.305 11.370 ;
      LAYER met4 ;
        RECT 2.985 11.050 3.305 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 10.620 3.305 10.940 ;
      LAYER met4 ;
        RECT 2.985 10.620 3.305 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 10.190 3.305 10.510 ;
      LAYER met4 ;
        RECT 2.985 10.190 3.305 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 9.760 3.305 10.080 ;
      LAYER met4 ;
        RECT 2.985 9.760 3.305 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 9.330 3.305 9.650 ;
      LAYER met4 ;
        RECT 2.985 9.330 3.305 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 8.900 3.305 9.220 ;
      LAYER met4 ;
        RECT 2.985 8.900 3.305 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 13.200 2.895 13.520 ;
      LAYER met4 ;
        RECT 2.575 13.200 2.895 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 12.770 2.895 13.090 ;
      LAYER met4 ;
        RECT 2.575 12.770 2.895 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 12.340 2.895 12.660 ;
      LAYER met4 ;
        RECT 2.575 12.340 2.895 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 11.910 2.895 12.230 ;
      LAYER met4 ;
        RECT 2.575 11.910 2.895 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 11.480 2.895 11.800 ;
      LAYER met4 ;
        RECT 2.575 11.480 2.895 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 11.050 2.895 11.370 ;
      LAYER met4 ;
        RECT 2.575 11.050 2.895 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 10.620 2.895 10.940 ;
      LAYER met4 ;
        RECT 2.575 10.620 2.895 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 10.190 2.895 10.510 ;
      LAYER met4 ;
        RECT 2.575 10.190 2.895 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 9.760 2.895 10.080 ;
      LAYER met4 ;
        RECT 2.575 9.760 2.895 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 9.330 2.895 9.650 ;
      LAYER met4 ;
        RECT 2.575 9.330 2.895 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 8.900 2.895 9.220 ;
      LAYER met4 ;
        RECT 2.575 8.900 2.895 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 13.200 2.485 13.520 ;
      LAYER met4 ;
        RECT 2.165 13.200 2.485 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 12.770 2.485 13.090 ;
      LAYER met4 ;
        RECT 2.165 12.770 2.485 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 12.340 2.485 12.660 ;
      LAYER met4 ;
        RECT 2.165 12.340 2.485 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 11.910 2.485 12.230 ;
      LAYER met4 ;
        RECT 2.165 11.910 2.485 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 11.480 2.485 11.800 ;
      LAYER met4 ;
        RECT 2.165 11.480 2.485 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 11.050 2.485 11.370 ;
      LAYER met4 ;
        RECT 2.165 11.050 2.485 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 10.620 2.485 10.940 ;
      LAYER met4 ;
        RECT 2.165 10.620 2.485 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 10.190 2.485 10.510 ;
      LAYER met4 ;
        RECT 2.165 10.190 2.485 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 9.760 2.485 10.080 ;
      LAYER met4 ;
        RECT 2.165 9.760 2.485 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 9.330 2.485 9.650 ;
      LAYER met4 ;
        RECT 2.165 9.330 2.485 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 8.900 2.485 9.220 ;
      LAYER met4 ;
        RECT 2.165 8.900 2.485 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 13.200 2.075 13.520 ;
      LAYER met4 ;
        RECT 1.755 13.200 2.075 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 12.770 2.075 13.090 ;
      LAYER met4 ;
        RECT 1.755 12.770 2.075 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 12.340 2.075 12.660 ;
      LAYER met4 ;
        RECT 1.755 12.340 2.075 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 11.910 2.075 12.230 ;
      LAYER met4 ;
        RECT 1.755 11.910 2.075 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 11.480 2.075 11.800 ;
      LAYER met4 ;
        RECT 1.755 11.480 2.075 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 11.050 2.075 11.370 ;
      LAYER met4 ;
        RECT 1.755 11.050 2.075 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 10.620 2.075 10.940 ;
      LAYER met4 ;
        RECT 1.755 10.620 2.075 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 10.190 2.075 10.510 ;
      LAYER met4 ;
        RECT 1.755 10.190 2.075 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 9.760 2.075 10.080 ;
      LAYER met4 ;
        RECT 1.755 9.760 2.075 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 9.330 2.075 9.650 ;
      LAYER met4 ;
        RECT 1.755 9.330 2.075 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 8.900 2.075 9.220 ;
      LAYER met4 ;
        RECT 1.755 8.900 2.075 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 13.200 1.665 13.520 ;
      LAYER met4 ;
        RECT 1.345 13.200 1.665 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 12.770 1.665 13.090 ;
      LAYER met4 ;
        RECT 1.345 12.770 1.665 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 12.340 1.665 12.660 ;
      LAYER met4 ;
        RECT 1.345 12.340 1.665 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 11.910 1.665 12.230 ;
      LAYER met4 ;
        RECT 1.345 11.910 1.665 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 11.480 1.665 11.800 ;
      LAYER met4 ;
        RECT 1.345 11.480 1.665 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 11.050 1.665 11.370 ;
      LAYER met4 ;
        RECT 1.345 11.050 1.665 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 10.620 1.665 10.940 ;
      LAYER met4 ;
        RECT 1.345 10.620 1.665 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 10.190 1.665 10.510 ;
      LAYER met4 ;
        RECT 1.345 10.190 1.665 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 9.760 1.665 10.080 ;
      LAYER met4 ;
        RECT 1.345 9.760 1.665 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 9.330 1.665 9.650 ;
      LAYER met4 ;
        RECT 1.345 9.330 1.665 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 8.900 1.665 9.220 ;
      LAYER met4 ;
        RECT 1.345 8.900 1.665 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 13.200 1.255 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 12.770 1.255 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 12.340 1.255 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 11.910 1.255 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 11.480 1.255 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 11.050 1.255 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 10.620 1.255 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 10.190 1.255 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 9.760 1.255 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 9.330 1.255 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 8.900 1.255 9.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 13.200 0.845 13.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 12.770 0.845 13.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 12.340 0.845 12.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 11.910 0.845 12.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 11.480 0.845 11.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 11.050 0.845 11.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 10.620 0.845 10.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 10.190 0.845 10.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 9.760 0.845 10.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 9.330 0.845 9.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 8.900 0.845 9.220 ;
    END
  END VCCD
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
  END VSWITCH
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
  END VSSIO_Q
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
  END VSSD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
  END VDDA
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.495 8.890 24.395 13.530 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 96.585 75.000 174.185 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__overlay_vccd_hvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vccd_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vccd_lvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
  END VDDIO
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
  END VSSA
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
  END VCCHIB
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 6.890 74.655 11.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 11.260 74.565 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 10.830 74.565 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 10.400 74.565 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 9.970 74.565 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 9.540 74.565 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 9.110 74.565 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 8.680 74.565 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 8.250 74.565 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 7.820 74.565 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 7.390 74.565 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 6.960 74.565 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 11.260 74.160 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 10.830 74.160 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 10.400 74.160 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 9.970 74.160 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 9.540 74.160 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 9.110 74.160 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 8.680 74.160 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 8.250 74.160 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 7.820 74.160 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 7.390 74.160 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 6.960 74.160 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 11.260 73.755 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 10.830 73.755 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 10.400 73.755 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 9.970 73.755 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 9.540 73.755 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 9.110 73.755 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 8.680 73.755 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 8.250 73.755 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 7.820 73.755 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 7.390 73.755 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 6.960 73.755 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 11.260 73.350 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 10.830 73.350 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 10.400 73.350 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 9.970 73.350 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 9.540 73.350 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 9.110 73.350 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 8.680 73.350 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 8.250 73.350 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 7.820 73.350 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 7.390 73.350 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 6.960 73.350 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 11.260 72.945 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 10.830 72.945 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 10.400 72.945 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 9.970 72.945 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 9.540 72.945 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 9.110 72.945 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 8.680 72.945 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 8.250 72.945 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 7.820 72.945 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 7.390 72.945 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 6.960 72.945 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 11.260 72.540 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 10.830 72.540 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 10.400 72.540 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 9.970 72.540 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 9.540 72.540 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 9.110 72.540 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 8.680 72.540 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 8.250 72.540 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 7.820 72.540 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 7.390 72.540 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 6.960 72.540 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 11.260 72.135 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 10.830 72.135 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 10.400 72.135 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 9.970 72.135 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 9.540 72.135 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 9.110 72.135 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 8.680 72.135 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 8.250 72.135 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 7.820 72.135 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 7.390 72.135 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 6.960 72.135 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 11.260 71.730 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 10.830 71.730 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 10.400 71.730 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 9.970 71.730 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 9.540 71.730 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 9.110 71.730 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 8.680 71.730 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 8.250 71.730 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 7.820 71.730 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 7.390 71.730 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 6.960 71.730 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 11.260 71.325 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 10.830 71.325 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 10.400 71.325 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 9.970 71.325 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 9.540 71.325 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 9.110 71.325 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 8.680 71.325 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 8.250 71.325 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 7.820 71.325 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 7.390 71.325 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 6.960 71.325 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 11.260 70.920 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 10.830 70.920 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 10.400 70.920 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 9.970 70.920 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 9.540 70.920 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 9.110 70.920 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 8.680 70.920 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 8.250 70.920 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 7.820 70.920 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 7.390 70.920 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 6.960 70.920 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 11.260 70.515 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 10.830 70.515 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 10.400 70.515 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 9.970 70.515 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 9.540 70.515 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 9.110 70.515 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 8.680 70.515 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 8.250 70.515 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 7.820 70.515 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 7.390 70.515 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 6.960 70.515 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 11.260 70.110 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 10.830 70.110 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 10.400 70.110 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 9.970 70.110 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 9.540 70.110 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 9.110 70.110 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 8.680 70.110 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 8.250 70.110 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 7.820 70.110 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 7.390 70.110 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 6.960 70.110 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 11.260 69.705 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 10.830 69.705 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 10.400 69.705 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 9.970 69.705 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 9.540 69.705 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 9.110 69.705 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 8.680 69.705 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 8.250 69.705 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 7.820 69.705 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 7.390 69.705 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 6.960 69.705 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 11.260 69.300 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 10.830 69.300 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 10.400 69.300 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 9.970 69.300 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 9.540 69.300 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 9.110 69.300 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 8.680 69.300 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 8.250 69.300 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 7.820 69.300 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 7.390 69.300 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 6.960 69.300 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 11.260 68.895 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 10.830 68.895 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 10.400 68.895 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 9.970 68.895 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 9.540 68.895 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 9.110 68.895 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 8.680 68.895 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 8.250 68.895 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 7.820 68.895 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 7.390 68.895 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 6.960 68.895 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 11.260 68.490 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 10.830 68.490 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 10.400 68.490 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 9.970 68.490 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 9.540 68.490 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 9.110 68.490 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 8.680 68.490 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 8.250 68.490 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 7.820 68.490 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 7.390 68.490 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 6.960 68.490 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 11.260 68.085 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 10.830 68.085 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 10.400 68.085 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 9.970 68.085 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 9.540 68.085 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 9.110 68.085 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 8.680 68.085 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 8.250 68.085 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 7.820 68.085 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 7.390 68.085 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 6.960 68.085 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 11.260 67.680 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 10.830 67.680 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 10.400 67.680 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 9.970 67.680 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 9.540 67.680 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 9.110 67.680 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 8.680 67.680 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 8.250 67.680 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 7.820 67.680 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 7.390 67.680 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 6.960 67.680 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 11.260 67.275 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 10.830 67.275 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 10.400 67.275 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 9.970 67.275 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 9.540 67.275 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 9.110 67.275 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 8.680 67.275 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 8.250 67.275 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 7.820 67.275 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 7.390 67.275 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 6.960 67.275 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 11.260 66.870 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 10.830 66.870 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 10.400 66.870 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 9.970 66.870 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 9.540 66.870 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 9.110 66.870 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 8.680 66.870 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 8.250 66.870 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 7.820 66.870 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 7.390 66.870 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 6.960 66.870 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 11.260 66.465 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 10.830 66.465 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 10.400 66.465 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 9.970 66.465 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 9.540 66.465 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 9.110 66.465 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 8.680 66.465 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 8.250 66.465 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 7.820 66.465 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 7.390 66.465 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 6.960 66.465 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 11.260 66.060 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 10.830 66.060 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 10.400 66.060 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 9.970 66.060 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 9.540 66.060 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 9.110 66.060 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 8.680 66.060 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 8.250 66.060 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 7.820 66.060 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 7.390 66.060 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 6.960 66.060 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 11.260 65.655 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 10.830 65.655 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 10.400 65.655 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 9.970 65.655 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 9.540 65.655 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 9.110 65.655 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 8.680 65.655 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 8.250 65.655 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 7.820 65.655 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 7.390 65.655 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 6.960 65.655 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 11.260 65.250 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 10.830 65.250 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 10.400 65.250 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 9.970 65.250 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 9.540 65.250 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 9.110 65.250 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 8.680 65.250 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 8.250 65.250 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 7.820 65.250 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 7.390 65.250 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 6.960 65.250 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 11.260 64.845 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 10.830 64.845 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 10.400 64.845 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 9.970 64.845 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 9.540 64.845 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 9.110 64.845 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 8.680 64.845 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 8.250 64.845 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 7.820 64.845 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 7.390 64.845 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 6.960 64.845 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 11.260 64.440 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 10.830 64.440 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 10.400 64.440 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 9.970 64.440 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 9.540 64.440 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 9.110 64.440 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 8.680 64.440 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 8.250 64.440 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 7.820 64.440 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 7.390 64.440 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 6.960 64.440 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 11.260 64.035 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 10.830 64.035 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 10.400 64.035 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 9.970 64.035 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 9.540 64.035 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 9.110 64.035 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 8.680 64.035 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 8.250 64.035 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 7.820 64.035 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 7.390 64.035 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 6.960 64.035 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 11.260 63.630 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 10.830 63.630 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 10.400 63.630 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 9.970 63.630 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 9.540 63.630 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 9.110 63.630 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 8.680 63.630 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 8.250 63.630 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 7.820 63.630 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 7.390 63.630 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 6.960 63.630 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 11.260 63.225 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 10.830 63.225 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 10.400 63.225 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 9.970 63.225 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 9.540 63.225 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 9.110 63.225 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 8.680 63.225 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 8.250 63.225 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 7.820 63.225 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 7.390 63.225 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 6.960 63.225 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 11.260 62.820 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 10.830 62.820 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 10.400 62.820 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 9.970 62.820 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 9.540 62.820 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 9.110 62.820 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 8.680 62.820 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 8.250 62.820 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 7.820 62.820 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 7.390 62.820 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 6.960 62.820 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 11.260 62.415 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 10.830 62.415 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 10.400 62.415 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 9.970 62.415 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 9.540 62.415 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 9.110 62.415 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 8.680 62.415 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 8.250 62.415 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 7.820 62.415 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 7.390 62.415 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 6.960 62.415 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 11.260 62.010 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 10.830 62.010 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 10.400 62.010 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 9.970 62.010 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 9.540 62.010 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 9.110 62.010 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 8.680 62.010 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 8.250 62.010 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 7.820 62.010 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 7.390 62.010 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 6.960 62.010 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 11.260 61.605 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 10.830 61.605 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 10.400 61.605 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 9.970 61.605 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 9.540 61.605 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 9.110 61.605 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 8.680 61.605 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 8.250 61.605 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 7.820 61.605 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 7.390 61.605 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 6.960 61.605 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 11.260 61.200 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 10.830 61.200 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 10.400 61.200 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 9.970 61.200 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 9.540 61.200 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 9.110 61.200 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 8.680 61.200 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 8.250 61.200 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 7.820 61.200 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 7.390 61.200 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 6.960 61.200 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 11.260 60.795 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 10.830 60.795 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 10.400 60.795 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 9.970 60.795 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 9.540 60.795 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 9.110 60.795 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 8.680 60.795 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 8.250 60.795 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 7.820 60.795 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 7.390 60.795 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 6.960 60.795 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 11.260 60.390 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 10.830 60.390 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 10.400 60.390 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 9.970 60.390 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 9.540 60.390 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 9.110 60.390 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 8.680 60.390 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 8.250 60.390 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 7.820 60.390 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 7.390 60.390 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 6.960 60.390 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 11.260 59.985 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 10.830 59.985 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 10.400 59.985 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 9.970 59.985 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 9.540 59.985 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 9.110 59.985 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 8.680 59.985 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 8.250 59.985 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 7.820 59.985 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 7.390 59.985 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 6.960 59.985 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 11.260 59.580 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 10.830 59.580 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 10.400 59.580 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 9.970 59.580 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 9.540 59.580 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 9.110 59.580 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 8.680 59.580 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 8.250 59.580 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 7.820 59.580 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 7.390 59.580 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 6.960 59.580 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 11.260 59.175 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 10.830 59.175 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 10.400 59.175 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 9.970 59.175 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 9.540 59.175 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 9.110 59.175 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 8.680 59.175 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 8.250 59.175 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 7.820 59.175 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 7.390 59.175 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 6.960 59.175 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 11.260 58.770 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 10.830 58.770 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 10.400 58.770 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 9.970 58.770 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 9.540 58.770 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 9.110 58.770 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 8.680 58.770 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 8.250 58.770 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 7.820 58.770 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 7.390 58.770 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 6.960 58.770 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 11.260 58.365 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 10.830 58.365 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 10.400 58.365 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 9.970 58.365 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 9.540 58.365 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 9.110 58.365 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 8.680 58.365 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 8.250 58.365 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 7.820 58.365 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 7.390 58.365 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 6.960 58.365 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 11.260 57.960 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 10.830 57.960 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 10.400 57.960 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 9.970 57.960 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 9.540 57.960 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 9.110 57.960 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 8.680 57.960 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 8.250 57.960 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 7.820 57.960 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 7.390 57.960 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 6.960 57.960 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 11.260 57.555 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 10.830 57.555 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 10.400 57.555 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 9.970 57.555 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 9.540 57.555 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 9.110 57.555 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 8.680 57.555 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 8.250 57.555 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 7.820 57.555 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 7.390 57.555 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 6.960 57.555 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 11.260 57.150 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 10.830 57.150 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 10.400 57.150 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 9.970 57.150 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 9.540 57.150 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 9.110 57.150 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 8.680 57.150 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 8.250 57.150 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 7.820 57.150 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 7.390 57.150 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 6.960 57.150 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 11.260 56.745 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 10.830 56.745 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 10.400 56.745 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 9.970 56.745 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 9.540 56.745 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 9.110 56.745 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 8.680 56.745 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 8.250 56.745 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 7.820 56.745 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 7.390 56.745 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 6.960 56.745 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 11.260 56.340 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 10.830 56.340 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 10.400 56.340 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 9.970 56.340 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 9.540 56.340 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 9.110 56.340 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 8.680 56.340 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 8.250 56.340 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 7.820 56.340 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 7.390 56.340 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 6.960 56.340 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 11.260 55.935 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 10.830 55.935 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 10.400 55.935 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 9.970 55.935 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 9.540 55.935 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 9.110 55.935 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 8.680 55.935 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 8.250 55.935 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 7.820 55.935 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 7.390 55.935 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 6.960 55.935 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 11.260 55.530 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 10.830 55.530 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 10.400 55.530 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 9.970 55.530 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 9.540 55.530 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 9.110 55.530 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 8.680 55.530 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 8.250 55.530 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 7.820 55.530 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 7.390 55.530 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 6.960 55.530 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 11.260 55.125 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 10.830 55.125 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 10.400 55.125 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 9.970 55.125 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 9.540 55.125 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 9.110 55.125 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 8.680 55.125 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 8.250 55.125 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 7.820 55.125 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 7.390 55.125 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 6.960 55.125 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 11.260 54.720 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 10.830 54.720 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 10.400 54.720 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 9.970 54.720 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 9.540 54.720 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 9.110 54.720 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 8.680 54.720 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 8.250 54.720 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 7.820 54.720 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 7.390 54.720 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 6.960 54.720 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 11.260 54.315 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 10.830 54.315 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 10.400 54.315 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 9.970 54.315 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 9.540 54.315 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 9.110 54.315 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 8.680 54.315 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 8.250 54.315 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 7.820 54.315 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 7.390 54.315 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 6.960 54.315 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 11.260 53.910 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 10.830 53.910 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 10.400 53.910 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 9.970 53.910 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 9.540 53.910 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 9.110 53.910 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 8.680 53.910 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 8.250 53.910 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 7.820 53.910 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 7.390 53.910 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 6.960 53.910 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 11.260 53.505 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 10.830 53.505 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 10.400 53.505 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 9.970 53.505 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 9.540 53.505 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 9.110 53.505 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 8.680 53.505 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 8.250 53.505 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 7.820 53.505 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 7.390 53.505 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 6.960 53.505 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 11.260 53.095 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 10.830 53.095 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 10.400 53.095 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 9.970 53.095 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 9.540 53.095 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 9.110 53.095 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 8.680 53.095 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 8.250 53.095 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 7.820 53.095 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 7.390 53.095 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 6.960 53.095 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 11.260 52.685 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 10.830 52.685 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 10.400 52.685 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 9.970 52.685 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 9.540 52.685 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 9.110 52.685 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 8.680 52.685 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 8.250 52.685 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 7.820 52.685 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 7.390 52.685 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 6.960 52.685 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 11.260 52.275 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 10.830 52.275 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 10.400 52.275 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 9.970 52.275 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 9.540 52.275 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 9.110 52.275 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 8.680 52.275 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 8.250 52.275 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 7.820 52.275 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 7.390 52.275 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 6.960 52.275 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 11.260 51.865 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 10.830 51.865 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 10.400 51.865 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 9.970 51.865 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 9.540 51.865 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 9.110 51.865 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 8.680 51.865 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 8.250 51.865 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 7.820 51.865 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 7.390 51.865 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 6.960 51.865 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 11.260 51.455 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 10.830 51.455 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 10.400 51.455 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 9.970 51.455 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 9.540 51.455 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 9.110 51.455 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 8.680 51.455 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 8.250 51.455 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 7.820 51.455 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 7.390 51.455 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 6.960 51.455 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 11.260 51.045 11.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 10.830 51.045 11.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 10.400 51.045 10.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 9.970 51.045 10.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 9.540 51.045 9.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 9.110 51.045 9.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 8.680 51.045 8.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 8.250 51.045 8.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 7.820 51.045 8.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 7.390 51.045 7.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 6.960 51.045 7.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 11.200 24.470 11.520 ;
      LAYER met4 ;
        RECT 24.150 11.200 24.470 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 10.770 24.470 11.090 ;
      LAYER met4 ;
        RECT 24.150 10.770 24.470 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 10.340 24.470 10.660 ;
      LAYER met4 ;
        RECT 24.150 10.340 24.470 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 9.910 24.470 10.230 ;
      LAYER met4 ;
        RECT 24.150 9.910 24.470 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 9.480 24.470 9.800 ;
      LAYER met4 ;
        RECT 24.150 9.480 24.470 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 9.050 24.470 9.370 ;
      LAYER met4 ;
        RECT 24.150 9.050 24.470 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 8.620 24.470 8.940 ;
      LAYER met4 ;
        RECT 24.150 8.620 24.470 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 8.190 24.470 8.510 ;
      LAYER met4 ;
        RECT 24.150 8.190 24.470 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 7.760 24.470 8.080 ;
      LAYER met4 ;
        RECT 24.150 7.760 24.470 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 7.330 24.470 7.650 ;
      LAYER met4 ;
        RECT 24.150 7.330 24.470 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 6.900 24.470 7.220 ;
      LAYER met4 ;
        RECT 24.150 6.900 24.470 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 11.200 24.065 11.520 ;
      LAYER met4 ;
        RECT 23.745 11.200 24.065 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 10.770 24.065 11.090 ;
      LAYER met4 ;
        RECT 23.745 10.770 24.065 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 10.340 24.065 10.660 ;
      LAYER met4 ;
        RECT 23.745 10.340 24.065 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 9.910 24.065 10.230 ;
      LAYER met4 ;
        RECT 23.745 9.910 24.065 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 9.480 24.065 9.800 ;
      LAYER met4 ;
        RECT 23.745 9.480 24.065 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 9.050 24.065 9.370 ;
      LAYER met4 ;
        RECT 23.745 9.050 24.065 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 8.620 24.065 8.940 ;
      LAYER met4 ;
        RECT 23.745 8.620 24.065 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 8.190 24.065 8.510 ;
      LAYER met4 ;
        RECT 23.745 8.190 24.065 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 7.760 24.065 8.080 ;
      LAYER met4 ;
        RECT 23.745 7.760 24.065 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 7.330 24.065 7.650 ;
      LAYER met4 ;
        RECT 23.745 7.330 24.065 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 6.900 24.065 7.220 ;
      LAYER met4 ;
        RECT 23.745 6.900 24.065 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 11.200 23.660 11.520 ;
      LAYER met4 ;
        RECT 23.340 11.200 23.660 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 10.770 23.660 11.090 ;
      LAYER met4 ;
        RECT 23.340 10.770 23.660 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 10.340 23.660 10.660 ;
      LAYER met4 ;
        RECT 23.340 10.340 23.660 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 9.910 23.660 10.230 ;
      LAYER met4 ;
        RECT 23.340 9.910 23.660 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 9.480 23.660 9.800 ;
      LAYER met4 ;
        RECT 23.340 9.480 23.660 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 9.050 23.660 9.370 ;
      LAYER met4 ;
        RECT 23.340 9.050 23.660 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 8.620 23.660 8.940 ;
      LAYER met4 ;
        RECT 23.340 8.620 23.660 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 8.190 23.660 8.510 ;
      LAYER met4 ;
        RECT 23.340 8.190 23.660 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 7.760 23.660 8.080 ;
      LAYER met4 ;
        RECT 23.340 7.760 23.660 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 7.330 23.660 7.650 ;
      LAYER met4 ;
        RECT 23.340 7.330 23.660 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 6.900 23.660 7.220 ;
      LAYER met4 ;
        RECT 23.340 6.900 23.660 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 11.200 23.255 11.520 ;
      LAYER met4 ;
        RECT 22.935 11.200 23.255 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 10.770 23.255 11.090 ;
      LAYER met4 ;
        RECT 22.935 10.770 23.255 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 10.340 23.255 10.660 ;
      LAYER met4 ;
        RECT 22.935 10.340 23.255 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 9.910 23.255 10.230 ;
      LAYER met4 ;
        RECT 22.935 9.910 23.255 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 9.480 23.255 9.800 ;
      LAYER met4 ;
        RECT 22.935 9.480 23.255 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 9.050 23.255 9.370 ;
      LAYER met4 ;
        RECT 22.935 9.050 23.255 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 8.620 23.255 8.940 ;
      LAYER met4 ;
        RECT 22.935 8.620 23.255 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 8.190 23.255 8.510 ;
      LAYER met4 ;
        RECT 22.935 8.190 23.255 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 7.760 23.255 8.080 ;
      LAYER met4 ;
        RECT 22.935 7.760 23.255 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 7.330 23.255 7.650 ;
      LAYER met4 ;
        RECT 22.935 7.330 23.255 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 6.900 23.255 7.220 ;
      LAYER met4 ;
        RECT 22.935 6.900 23.255 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 11.200 22.850 11.520 ;
      LAYER met4 ;
        RECT 22.530 11.200 22.850 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 10.770 22.850 11.090 ;
      LAYER met4 ;
        RECT 22.530 10.770 22.850 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 10.340 22.850 10.660 ;
      LAYER met4 ;
        RECT 22.530 10.340 22.850 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 9.910 22.850 10.230 ;
      LAYER met4 ;
        RECT 22.530 9.910 22.850 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 9.480 22.850 9.800 ;
      LAYER met4 ;
        RECT 22.530 9.480 22.850 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 9.050 22.850 9.370 ;
      LAYER met4 ;
        RECT 22.530 9.050 22.850 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 8.620 22.850 8.940 ;
      LAYER met4 ;
        RECT 22.530 8.620 22.850 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 8.190 22.850 8.510 ;
      LAYER met4 ;
        RECT 22.530 8.190 22.850 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 7.760 22.850 8.080 ;
      LAYER met4 ;
        RECT 22.530 7.760 22.850 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 7.330 22.850 7.650 ;
      LAYER met4 ;
        RECT 22.530 7.330 22.850 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 6.900 22.850 7.220 ;
      LAYER met4 ;
        RECT 22.530 6.900 22.850 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 11.200 22.445 11.520 ;
      LAYER met4 ;
        RECT 22.125 11.200 22.445 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 10.770 22.445 11.090 ;
      LAYER met4 ;
        RECT 22.125 10.770 22.445 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 10.340 22.445 10.660 ;
      LAYER met4 ;
        RECT 22.125 10.340 22.445 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 9.910 22.445 10.230 ;
      LAYER met4 ;
        RECT 22.125 9.910 22.445 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 9.480 22.445 9.800 ;
      LAYER met4 ;
        RECT 22.125 9.480 22.445 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 9.050 22.445 9.370 ;
      LAYER met4 ;
        RECT 22.125 9.050 22.445 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 8.620 22.445 8.940 ;
      LAYER met4 ;
        RECT 22.125 8.620 22.445 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 8.190 22.445 8.510 ;
      LAYER met4 ;
        RECT 22.125 8.190 22.445 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 7.760 22.445 8.080 ;
      LAYER met4 ;
        RECT 22.125 7.760 22.445 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 7.330 22.445 7.650 ;
      LAYER met4 ;
        RECT 22.125 7.330 22.445 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 6.900 22.445 7.220 ;
      LAYER met4 ;
        RECT 22.125 6.900 22.445 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 11.200 22.040 11.520 ;
      LAYER met4 ;
        RECT 21.720 11.200 22.040 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 10.770 22.040 11.090 ;
      LAYER met4 ;
        RECT 21.720 10.770 22.040 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 10.340 22.040 10.660 ;
      LAYER met4 ;
        RECT 21.720 10.340 22.040 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 9.910 22.040 10.230 ;
      LAYER met4 ;
        RECT 21.720 9.910 22.040 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 9.480 22.040 9.800 ;
      LAYER met4 ;
        RECT 21.720 9.480 22.040 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 9.050 22.040 9.370 ;
      LAYER met4 ;
        RECT 21.720 9.050 22.040 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 8.620 22.040 8.940 ;
      LAYER met4 ;
        RECT 21.720 8.620 22.040 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 8.190 22.040 8.510 ;
      LAYER met4 ;
        RECT 21.720 8.190 22.040 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 7.760 22.040 8.080 ;
      LAYER met4 ;
        RECT 21.720 7.760 22.040 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 7.330 22.040 7.650 ;
      LAYER met4 ;
        RECT 21.720 7.330 22.040 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 6.900 22.040 7.220 ;
      LAYER met4 ;
        RECT 21.720 6.900 22.040 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 11.200 21.635 11.520 ;
      LAYER met4 ;
        RECT 21.315 11.200 21.635 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 10.770 21.635 11.090 ;
      LAYER met4 ;
        RECT 21.315 10.770 21.635 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 10.340 21.635 10.660 ;
      LAYER met4 ;
        RECT 21.315 10.340 21.635 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 9.910 21.635 10.230 ;
      LAYER met4 ;
        RECT 21.315 9.910 21.635 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 9.480 21.635 9.800 ;
      LAYER met4 ;
        RECT 21.315 9.480 21.635 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 9.050 21.635 9.370 ;
      LAYER met4 ;
        RECT 21.315 9.050 21.635 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 8.620 21.635 8.940 ;
      LAYER met4 ;
        RECT 21.315 8.620 21.635 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 8.190 21.635 8.510 ;
      LAYER met4 ;
        RECT 21.315 8.190 21.635 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 7.760 21.635 8.080 ;
      LAYER met4 ;
        RECT 21.315 7.760 21.635 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 7.330 21.635 7.650 ;
      LAYER met4 ;
        RECT 21.315 7.330 21.635 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 6.900 21.635 7.220 ;
      LAYER met4 ;
        RECT 21.315 6.900 21.635 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 11.200 21.230 11.520 ;
      LAYER met4 ;
        RECT 20.910 11.200 21.230 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 10.770 21.230 11.090 ;
      LAYER met4 ;
        RECT 20.910 10.770 21.230 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 10.340 21.230 10.660 ;
      LAYER met4 ;
        RECT 20.910 10.340 21.230 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 9.910 21.230 10.230 ;
      LAYER met4 ;
        RECT 20.910 9.910 21.230 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 9.480 21.230 9.800 ;
      LAYER met4 ;
        RECT 20.910 9.480 21.230 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 9.050 21.230 9.370 ;
      LAYER met4 ;
        RECT 20.910 9.050 21.230 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 8.620 21.230 8.940 ;
      LAYER met4 ;
        RECT 20.910 8.620 21.230 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 8.190 21.230 8.510 ;
      LAYER met4 ;
        RECT 20.910 8.190 21.230 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 7.760 21.230 8.080 ;
      LAYER met4 ;
        RECT 20.910 7.760 21.230 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 7.330 21.230 7.650 ;
      LAYER met4 ;
        RECT 20.910 7.330 21.230 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 6.900 21.230 7.220 ;
      LAYER met4 ;
        RECT 20.910 6.900 21.230 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 11.200 20.825 11.520 ;
      LAYER met4 ;
        RECT 20.505 11.200 20.825 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 10.770 20.825 11.090 ;
      LAYER met4 ;
        RECT 20.505 10.770 20.825 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 10.340 20.825 10.660 ;
      LAYER met4 ;
        RECT 20.505 10.340 20.825 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 9.910 20.825 10.230 ;
      LAYER met4 ;
        RECT 20.505 9.910 20.825 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 9.480 20.825 9.800 ;
      LAYER met4 ;
        RECT 20.505 9.480 20.825 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 9.050 20.825 9.370 ;
      LAYER met4 ;
        RECT 20.505 9.050 20.825 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 8.620 20.825 8.940 ;
      LAYER met4 ;
        RECT 20.505 8.620 20.825 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 8.190 20.825 8.510 ;
      LAYER met4 ;
        RECT 20.505 8.190 20.825 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 7.760 20.825 8.080 ;
      LAYER met4 ;
        RECT 20.505 7.760 20.825 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 7.330 20.825 7.650 ;
      LAYER met4 ;
        RECT 20.505 7.330 20.825 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 6.900 20.825 7.220 ;
      LAYER met4 ;
        RECT 20.505 6.900 20.825 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 11.200 20.420 11.520 ;
      LAYER met4 ;
        RECT 20.100 11.200 20.420 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 10.770 20.420 11.090 ;
      LAYER met4 ;
        RECT 20.100 10.770 20.420 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 10.340 20.420 10.660 ;
      LAYER met4 ;
        RECT 20.100 10.340 20.420 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 9.910 20.420 10.230 ;
      LAYER met4 ;
        RECT 20.100 9.910 20.420 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 9.480 20.420 9.800 ;
      LAYER met4 ;
        RECT 20.100 9.480 20.420 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 9.050 20.420 9.370 ;
      LAYER met4 ;
        RECT 20.100 9.050 20.420 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 8.620 20.420 8.940 ;
      LAYER met4 ;
        RECT 20.100 8.620 20.420 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 8.190 20.420 8.510 ;
      LAYER met4 ;
        RECT 20.100 8.190 20.420 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 7.760 20.420 8.080 ;
      LAYER met4 ;
        RECT 20.100 7.760 20.420 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 7.330 20.420 7.650 ;
      LAYER met4 ;
        RECT 20.100 7.330 20.420 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 6.900 20.420 7.220 ;
      LAYER met4 ;
        RECT 20.100 6.900 20.420 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 11.200 20.015 11.520 ;
      LAYER met4 ;
        RECT 19.695 11.200 20.015 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 10.770 20.015 11.090 ;
      LAYER met4 ;
        RECT 19.695 10.770 20.015 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 10.340 20.015 10.660 ;
      LAYER met4 ;
        RECT 19.695 10.340 20.015 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 9.910 20.015 10.230 ;
      LAYER met4 ;
        RECT 19.695 9.910 20.015 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 9.480 20.015 9.800 ;
      LAYER met4 ;
        RECT 19.695 9.480 20.015 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 9.050 20.015 9.370 ;
      LAYER met4 ;
        RECT 19.695 9.050 20.015 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 8.620 20.015 8.940 ;
      LAYER met4 ;
        RECT 19.695 8.620 20.015 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 8.190 20.015 8.510 ;
      LAYER met4 ;
        RECT 19.695 8.190 20.015 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 7.760 20.015 8.080 ;
      LAYER met4 ;
        RECT 19.695 7.760 20.015 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 7.330 20.015 7.650 ;
      LAYER met4 ;
        RECT 19.695 7.330 20.015 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 6.900 20.015 7.220 ;
      LAYER met4 ;
        RECT 19.695 6.900 20.015 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 11.200 19.610 11.520 ;
      LAYER met4 ;
        RECT 19.290 11.200 19.610 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 10.770 19.610 11.090 ;
      LAYER met4 ;
        RECT 19.290 10.770 19.610 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 10.340 19.610 10.660 ;
      LAYER met4 ;
        RECT 19.290 10.340 19.610 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 9.910 19.610 10.230 ;
      LAYER met4 ;
        RECT 19.290 9.910 19.610 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 9.480 19.610 9.800 ;
      LAYER met4 ;
        RECT 19.290 9.480 19.610 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 9.050 19.610 9.370 ;
      LAYER met4 ;
        RECT 19.290 9.050 19.610 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 8.620 19.610 8.940 ;
      LAYER met4 ;
        RECT 19.290 8.620 19.610 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 8.190 19.610 8.510 ;
      LAYER met4 ;
        RECT 19.290 8.190 19.610 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 7.760 19.610 8.080 ;
      LAYER met4 ;
        RECT 19.290 7.760 19.610 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 7.330 19.610 7.650 ;
      LAYER met4 ;
        RECT 19.290 7.330 19.610 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 6.900 19.610 7.220 ;
      LAYER met4 ;
        RECT 19.290 6.900 19.610 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 11.200 19.205 11.520 ;
      LAYER met4 ;
        RECT 18.885 11.200 19.205 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 10.770 19.205 11.090 ;
      LAYER met4 ;
        RECT 18.885 10.770 19.205 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 10.340 19.205 10.660 ;
      LAYER met4 ;
        RECT 18.885 10.340 19.205 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 9.910 19.205 10.230 ;
      LAYER met4 ;
        RECT 18.885 9.910 19.205 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 9.480 19.205 9.800 ;
      LAYER met4 ;
        RECT 18.885 9.480 19.205 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 9.050 19.205 9.370 ;
      LAYER met4 ;
        RECT 18.885 9.050 19.205 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 8.620 19.205 8.940 ;
      LAYER met4 ;
        RECT 18.885 8.620 19.205 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 8.190 19.205 8.510 ;
      LAYER met4 ;
        RECT 18.885 8.190 19.205 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 7.760 19.205 8.080 ;
      LAYER met4 ;
        RECT 18.885 7.760 19.205 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 7.330 19.205 7.650 ;
      LAYER met4 ;
        RECT 18.885 7.330 19.205 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 6.900 19.205 7.220 ;
      LAYER met4 ;
        RECT 18.885 6.900 19.205 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 11.200 18.800 11.520 ;
      LAYER met4 ;
        RECT 18.480 11.200 18.800 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 10.770 18.800 11.090 ;
      LAYER met4 ;
        RECT 18.480 10.770 18.800 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 10.340 18.800 10.660 ;
      LAYER met4 ;
        RECT 18.480 10.340 18.800 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 9.910 18.800 10.230 ;
      LAYER met4 ;
        RECT 18.480 9.910 18.800 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 9.480 18.800 9.800 ;
      LAYER met4 ;
        RECT 18.480 9.480 18.800 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 9.050 18.800 9.370 ;
      LAYER met4 ;
        RECT 18.480 9.050 18.800 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 8.620 18.800 8.940 ;
      LAYER met4 ;
        RECT 18.480 8.620 18.800 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 8.190 18.800 8.510 ;
      LAYER met4 ;
        RECT 18.480 8.190 18.800 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 7.760 18.800 8.080 ;
      LAYER met4 ;
        RECT 18.480 7.760 18.800 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 7.330 18.800 7.650 ;
      LAYER met4 ;
        RECT 18.480 7.330 18.800 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 6.900 18.800 7.220 ;
      LAYER met4 ;
        RECT 18.480 6.900 18.800 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 11.200 18.395 11.520 ;
      LAYER met4 ;
        RECT 18.075 11.200 18.395 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 10.770 18.395 11.090 ;
      LAYER met4 ;
        RECT 18.075 10.770 18.395 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 10.340 18.395 10.660 ;
      LAYER met4 ;
        RECT 18.075 10.340 18.395 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 9.910 18.395 10.230 ;
      LAYER met4 ;
        RECT 18.075 9.910 18.395 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 9.480 18.395 9.800 ;
      LAYER met4 ;
        RECT 18.075 9.480 18.395 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 9.050 18.395 9.370 ;
      LAYER met4 ;
        RECT 18.075 9.050 18.395 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 8.620 18.395 8.940 ;
      LAYER met4 ;
        RECT 18.075 8.620 18.395 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 8.190 18.395 8.510 ;
      LAYER met4 ;
        RECT 18.075 8.190 18.395 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 7.760 18.395 8.080 ;
      LAYER met4 ;
        RECT 18.075 7.760 18.395 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 7.330 18.395 7.650 ;
      LAYER met4 ;
        RECT 18.075 7.330 18.395 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 6.900 18.395 7.220 ;
      LAYER met4 ;
        RECT 18.075 6.900 18.395 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 11.200 17.990 11.520 ;
      LAYER met4 ;
        RECT 17.670 11.200 17.990 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 10.770 17.990 11.090 ;
      LAYER met4 ;
        RECT 17.670 10.770 17.990 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 10.340 17.990 10.660 ;
      LAYER met4 ;
        RECT 17.670 10.340 17.990 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 9.910 17.990 10.230 ;
      LAYER met4 ;
        RECT 17.670 9.910 17.990 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 9.480 17.990 9.800 ;
      LAYER met4 ;
        RECT 17.670 9.480 17.990 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 9.050 17.990 9.370 ;
      LAYER met4 ;
        RECT 17.670 9.050 17.990 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 8.620 17.990 8.940 ;
      LAYER met4 ;
        RECT 17.670 8.620 17.990 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 8.190 17.990 8.510 ;
      LAYER met4 ;
        RECT 17.670 8.190 17.990 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 7.760 17.990 8.080 ;
      LAYER met4 ;
        RECT 17.670 7.760 17.990 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 7.330 17.990 7.650 ;
      LAYER met4 ;
        RECT 17.670 7.330 17.990 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 6.900 17.990 7.220 ;
      LAYER met4 ;
        RECT 17.670 6.900 17.990 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 11.200 17.585 11.520 ;
      LAYER met4 ;
        RECT 17.265 11.200 17.585 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 10.770 17.585 11.090 ;
      LAYER met4 ;
        RECT 17.265 10.770 17.585 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 10.340 17.585 10.660 ;
      LAYER met4 ;
        RECT 17.265 10.340 17.585 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 9.910 17.585 10.230 ;
      LAYER met4 ;
        RECT 17.265 9.910 17.585 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 9.480 17.585 9.800 ;
      LAYER met4 ;
        RECT 17.265 9.480 17.585 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 9.050 17.585 9.370 ;
      LAYER met4 ;
        RECT 17.265 9.050 17.585 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 8.620 17.585 8.940 ;
      LAYER met4 ;
        RECT 17.265 8.620 17.585 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 8.190 17.585 8.510 ;
      LAYER met4 ;
        RECT 17.265 8.190 17.585 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 7.760 17.585 8.080 ;
      LAYER met4 ;
        RECT 17.265 7.760 17.585 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 7.330 17.585 7.650 ;
      LAYER met4 ;
        RECT 17.265 7.330 17.585 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 6.900 17.585 7.220 ;
      LAYER met4 ;
        RECT 17.265 6.900 17.585 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 11.200 17.180 11.520 ;
      LAYER met4 ;
        RECT 16.860 11.200 17.180 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 10.770 17.180 11.090 ;
      LAYER met4 ;
        RECT 16.860 10.770 17.180 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 10.340 17.180 10.660 ;
      LAYER met4 ;
        RECT 16.860 10.340 17.180 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 9.910 17.180 10.230 ;
      LAYER met4 ;
        RECT 16.860 9.910 17.180 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 9.480 17.180 9.800 ;
      LAYER met4 ;
        RECT 16.860 9.480 17.180 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 9.050 17.180 9.370 ;
      LAYER met4 ;
        RECT 16.860 9.050 17.180 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 8.620 17.180 8.940 ;
      LAYER met4 ;
        RECT 16.860 8.620 17.180 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 8.190 17.180 8.510 ;
      LAYER met4 ;
        RECT 16.860 8.190 17.180 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 7.760 17.180 8.080 ;
      LAYER met4 ;
        RECT 16.860 7.760 17.180 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 7.330 17.180 7.650 ;
      LAYER met4 ;
        RECT 16.860 7.330 17.180 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 6.900 17.180 7.220 ;
      LAYER met4 ;
        RECT 16.860 6.900 17.180 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 11.200 16.775 11.520 ;
      LAYER met4 ;
        RECT 16.455 11.200 16.775 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 10.770 16.775 11.090 ;
      LAYER met4 ;
        RECT 16.455 10.770 16.775 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 10.340 16.775 10.660 ;
      LAYER met4 ;
        RECT 16.455 10.340 16.775 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 9.910 16.775 10.230 ;
      LAYER met4 ;
        RECT 16.455 9.910 16.775 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 9.480 16.775 9.800 ;
      LAYER met4 ;
        RECT 16.455 9.480 16.775 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 9.050 16.775 9.370 ;
      LAYER met4 ;
        RECT 16.455 9.050 16.775 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 8.620 16.775 8.940 ;
      LAYER met4 ;
        RECT 16.455 8.620 16.775 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 8.190 16.775 8.510 ;
      LAYER met4 ;
        RECT 16.455 8.190 16.775 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 7.760 16.775 8.080 ;
      LAYER met4 ;
        RECT 16.455 7.760 16.775 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 7.330 16.775 7.650 ;
      LAYER met4 ;
        RECT 16.455 7.330 16.775 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 6.900 16.775 7.220 ;
      LAYER met4 ;
        RECT 16.455 6.900 16.775 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 11.200 16.370 11.520 ;
      LAYER met4 ;
        RECT 16.050 11.200 16.370 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 10.770 16.370 11.090 ;
      LAYER met4 ;
        RECT 16.050 10.770 16.370 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 10.340 16.370 10.660 ;
      LAYER met4 ;
        RECT 16.050 10.340 16.370 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 9.910 16.370 10.230 ;
      LAYER met4 ;
        RECT 16.050 9.910 16.370 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 9.480 16.370 9.800 ;
      LAYER met4 ;
        RECT 16.050 9.480 16.370 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 9.050 16.370 9.370 ;
      LAYER met4 ;
        RECT 16.050 9.050 16.370 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 8.620 16.370 8.940 ;
      LAYER met4 ;
        RECT 16.050 8.620 16.370 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 8.190 16.370 8.510 ;
      LAYER met4 ;
        RECT 16.050 8.190 16.370 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 7.760 16.370 8.080 ;
      LAYER met4 ;
        RECT 16.050 7.760 16.370 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 7.330 16.370 7.650 ;
      LAYER met4 ;
        RECT 16.050 7.330 16.370 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 6.900 16.370 7.220 ;
      LAYER met4 ;
        RECT 16.050 6.900 16.370 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 11.200 15.965 11.520 ;
      LAYER met4 ;
        RECT 15.645 11.200 15.965 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 10.770 15.965 11.090 ;
      LAYER met4 ;
        RECT 15.645 10.770 15.965 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 10.340 15.965 10.660 ;
      LAYER met4 ;
        RECT 15.645 10.340 15.965 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 9.910 15.965 10.230 ;
      LAYER met4 ;
        RECT 15.645 9.910 15.965 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 9.480 15.965 9.800 ;
      LAYER met4 ;
        RECT 15.645 9.480 15.965 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 9.050 15.965 9.370 ;
      LAYER met4 ;
        RECT 15.645 9.050 15.965 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 8.620 15.965 8.940 ;
      LAYER met4 ;
        RECT 15.645 8.620 15.965 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 8.190 15.965 8.510 ;
      LAYER met4 ;
        RECT 15.645 8.190 15.965 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 7.760 15.965 8.080 ;
      LAYER met4 ;
        RECT 15.645 7.760 15.965 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 7.330 15.965 7.650 ;
      LAYER met4 ;
        RECT 15.645 7.330 15.965 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 6.900 15.965 7.220 ;
      LAYER met4 ;
        RECT 15.645 6.900 15.965 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 11.200 15.560 11.520 ;
      LAYER met4 ;
        RECT 15.240 11.200 15.560 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 10.770 15.560 11.090 ;
      LAYER met4 ;
        RECT 15.240 10.770 15.560 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 10.340 15.560 10.660 ;
      LAYER met4 ;
        RECT 15.240 10.340 15.560 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 9.910 15.560 10.230 ;
      LAYER met4 ;
        RECT 15.240 9.910 15.560 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 9.480 15.560 9.800 ;
      LAYER met4 ;
        RECT 15.240 9.480 15.560 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 9.050 15.560 9.370 ;
      LAYER met4 ;
        RECT 15.240 9.050 15.560 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 8.620 15.560 8.940 ;
      LAYER met4 ;
        RECT 15.240 8.620 15.560 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 8.190 15.560 8.510 ;
      LAYER met4 ;
        RECT 15.240 8.190 15.560 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 7.760 15.560 8.080 ;
      LAYER met4 ;
        RECT 15.240 7.760 15.560 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 7.330 15.560 7.650 ;
      LAYER met4 ;
        RECT 15.240 7.330 15.560 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 6.900 15.560 7.220 ;
      LAYER met4 ;
        RECT 15.240 6.900 15.560 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 11.200 15.155 11.520 ;
      LAYER met4 ;
        RECT 14.835 11.200 15.155 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 10.770 15.155 11.090 ;
      LAYER met4 ;
        RECT 14.835 10.770 15.155 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 10.340 15.155 10.660 ;
      LAYER met4 ;
        RECT 14.835 10.340 15.155 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 9.910 15.155 10.230 ;
      LAYER met4 ;
        RECT 14.835 9.910 15.155 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 9.480 15.155 9.800 ;
      LAYER met4 ;
        RECT 14.835 9.480 15.155 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 9.050 15.155 9.370 ;
      LAYER met4 ;
        RECT 14.835 9.050 15.155 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 8.620 15.155 8.940 ;
      LAYER met4 ;
        RECT 14.835 8.620 15.155 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 8.190 15.155 8.510 ;
      LAYER met4 ;
        RECT 14.835 8.190 15.155 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 7.760 15.155 8.080 ;
      LAYER met4 ;
        RECT 14.835 7.760 15.155 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 7.330 15.155 7.650 ;
      LAYER met4 ;
        RECT 14.835 7.330 15.155 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 6.900 15.155 7.220 ;
      LAYER met4 ;
        RECT 14.835 6.900 15.155 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 11.200 14.750 11.520 ;
      LAYER met4 ;
        RECT 14.430 11.200 14.750 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 10.770 14.750 11.090 ;
      LAYER met4 ;
        RECT 14.430 10.770 14.750 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 10.340 14.750 10.660 ;
      LAYER met4 ;
        RECT 14.430 10.340 14.750 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 9.910 14.750 10.230 ;
      LAYER met4 ;
        RECT 14.430 9.910 14.750 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 9.480 14.750 9.800 ;
      LAYER met4 ;
        RECT 14.430 9.480 14.750 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 9.050 14.750 9.370 ;
      LAYER met4 ;
        RECT 14.430 9.050 14.750 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 8.620 14.750 8.940 ;
      LAYER met4 ;
        RECT 14.430 8.620 14.750 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 8.190 14.750 8.510 ;
      LAYER met4 ;
        RECT 14.430 8.190 14.750 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 7.760 14.750 8.080 ;
      LAYER met4 ;
        RECT 14.430 7.760 14.750 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 7.330 14.750 7.650 ;
      LAYER met4 ;
        RECT 14.430 7.330 14.750 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 6.900 14.750 7.220 ;
      LAYER met4 ;
        RECT 14.430 6.900 14.750 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 11.200 14.345 11.520 ;
      LAYER met4 ;
        RECT 14.025 11.200 14.345 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 10.770 14.345 11.090 ;
      LAYER met4 ;
        RECT 14.025 10.770 14.345 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 10.340 14.345 10.660 ;
      LAYER met4 ;
        RECT 14.025 10.340 14.345 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 9.910 14.345 10.230 ;
      LAYER met4 ;
        RECT 14.025 9.910 14.345 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 9.480 14.345 9.800 ;
      LAYER met4 ;
        RECT 14.025 9.480 14.345 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 9.050 14.345 9.370 ;
      LAYER met4 ;
        RECT 14.025 9.050 14.345 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 8.620 14.345 8.940 ;
      LAYER met4 ;
        RECT 14.025 8.620 14.345 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 8.190 14.345 8.510 ;
      LAYER met4 ;
        RECT 14.025 8.190 14.345 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 7.760 14.345 8.080 ;
      LAYER met4 ;
        RECT 14.025 7.760 14.345 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 7.330 14.345 7.650 ;
      LAYER met4 ;
        RECT 14.025 7.330 14.345 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 6.900 14.345 7.220 ;
      LAYER met4 ;
        RECT 14.025 6.900 14.345 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 11.200 13.940 11.520 ;
      LAYER met4 ;
        RECT 13.620 11.200 13.940 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 10.770 13.940 11.090 ;
      LAYER met4 ;
        RECT 13.620 10.770 13.940 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 10.340 13.940 10.660 ;
      LAYER met4 ;
        RECT 13.620 10.340 13.940 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 9.910 13.940 10.230 ;
      LAYER met4 ;
        RECT 13.620 9.910 13.940 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 9.480 13.940 9.800 ;
      LAYER met4 ;
        RECT 13.620 9.480 13.940 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 9.050 13.940 9.370 ;
      LAYER met4 ;
        RECT 13.620 9.050 13.940 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 8.620 13.940 8.940 ;
      LAYER met4 ;
        RECT 13.620 8.620 13.940 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 8.190 13.940 8.510 ;
      LAYER met4 ;
        RECT 13.620 8.190 13.940 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 7.760 13.940 8.080 ;
      LAYER met4 ;
        RECT 13.620 7.760 13.940 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 7.330 13.940 7.650 ;
      LAYER met4 ;
        RECT 13.620 7.330 13.940 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 6.900 13.940 7.220 ;
      LAYER met4 ;
        RECT 13.620 6.900 13.940 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 11.200 13.535 11.520 ;
      LAYER met4 ;
        RECT 13.215 11.200 13.535 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 10.770 13.535 11.090 ;
      LAYER met4 ;
        RECT 13.215 10.770 13.535 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 10.340 13.535 10.660 ;
      LAYER met4 ;
        RECT 13.215 10.340 13.535 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 9.910 13.535 10.230 ;
      LAYER met4 ;
        RECT 13.215 9.910 13.535 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 9.480 13.535 9.800 ;
      LAYER met4 ;
        RECT 13.215 9.480 13.535 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 9.050 13.535 9.370 ;
      LAYER met4 ;
        RECT 13.215 9.050 13.535 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 8.620 13.535 8.940 ;
      LAYER met4 ;
        RECT 13.215 8.620 13.535 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 8.190 13.535 8.510 ;
      LAYER met4 ;
        RECT 13.215 8.190 13.535 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 7.760 13.535 8.080 ;
      LAYER met4 ;
        RECT 13.215 7.760 13.535 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 7.330 13.535 7.650 ;
      LAYER met4 ;
        RECT 13.215 7.330 13.535 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 6.900 13.535 7.220 ;
      LAYER met4 ;
        RECT 13.215 6.900 13.535 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 11.200 13.130 11.520 ;
      LAYER met4 ;
        RECT 12.810 11.200 13.130 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 10.770 13.130 11.090 ;
      LAYER met4 ;
        RECT 12.810 10.770 13.130 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 10.340 13.130 10.660 ;
      LAYER met4 ;
        RECT 12.810 10.340 13.130 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 9.910 13.130 10.230 ;
      LAYER met4 ;
        RECT 12.810 9.910 13.130 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 9.480 13.130 9.800 ;
      LAYER met4 ;
        RECT 12.810 9.480 13.130 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 9.050 13.130 9.370 ;
      LAYER met4 ;
        RECT 12.810 9.050 13.130 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 8.620 13.130 8.940 ;
      LAYER met4 ;
        RECT 12.810 8.620 13.130 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 8.190 13.130 8.510 ;
      LAYER met4 ;
        RECT 12.810 8.190 13.130 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 7.760 13.130 8.080 ;
      LAYER met4 ;
        RECT 12.810 7.760 13.130 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 7.330 13.130 7.650 ;
      LAYER met4 ;
        RECT 12.810 7.330 13.130 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 6.900 13.130 7.220 ;
      LAYER met4 ;
        RECT 12.810 6.900 13.130 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 11.200 12.725 11.520 ;
      LAYER met4 ;
        RECT 12.405 11.200 12.725 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 10.770 12.725 11.090 ;
      LAYER met4 ;
        RECT 12.405 10.770 12.725 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 10.340 12.725 10.660 ;
      LAYER met4 ;
        RECT 12.405 10.340 12.725 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 9.910 12.725 10.230 ;
      LAYER met4 ;
        RECT 12.405 9.910 12.725 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 9.480 12.725 9.800 ;
      LAYER met4 ;
        RECT 12.405 9.480 12.725 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 9.050 12.725 9.370 ;
      LAYER met4 ;
        RECT 12.405 9.050 12.725 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 8.620 12.725 8.940 ;
      LAYER met4 ;
        RECT 12.405 8.620 12.725 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 8.190 12.725 8.510 ;
      LAYER met4 ;
        RECT 12.405 8.190 12.725 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 7.760 12.725 8.080 ;
      LAYER met4 ;
        RECT 12.405 7.760 12.725 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 7.330 12.725 7.650 ;
      LAYER met4 ;
        RECT 12.405 7.330 12.725 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 6.900 12.725 7.220 ;
      LAYER met4 ;
        RECT 12.405 6.900 12.725 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 11.200 12.320 11.520 ;
      LAYER met4 ;
        RECT 12.000 11.200 12.320 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 10.770 12.320 11.090 ;
      LAYER met4 ;
        RECT 12.000 10.770 12.320 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 10.340 12.320 10.660 ;
      LAYER met4 ;
        RECT 12.000 10.340 12.320 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 9.910 12.320 10.230 ;
      LAYER met4 ;
        RECT 12.000 9.910 12.320 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 9.480 12.320 9.800 ;
      LAYER met4 ;
        RECT 12.000 9.480 12.320 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 9.050 12.320 9.370 ;
      LAYER met4 ;
        RECT 12.000 9.050 12.320 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 8.620 12.320 8.940 ;
      LAYER met4 ;
        RECT 12.000 8.620 12.320 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 8.190 12.320 8.510 ;
      LAYER met4 ;
        RECT 12.000 8.190 12.320 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 7.760 12.320 8.080 ;
      LAYER met4 ;
        RECT 12.000 7.760 12.320 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 7.330 12.320 7.650 ;
      LAYER met4 ;
        RECT 12.000 7.330 12.320 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 6.900 12.320 7.220 ;
      LAYER met4 ;
        RECT 12.000 6.900 12.320 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 11.200 11.915 11.520 ;
      LAYER met4 ;
        RECT 11.595 11.200 11.915 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 10.770 11.915 11.090 ;
      LAYER met4 ;
        RECT 11.595 10.770 11.915 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 10.340 11.915 10.660 ;
      LAYER met4 ;
        RECT 11.595 10.340 11.915 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 9.910 11.915 10.230 ;
      LAYER met4 ;
        RECT 11.595 9.910 11.915 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 9.480 11.915 9.800 ;
      LAYER met4 ;
        RECT 11.595 9.480 11.915 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 9.050 11.915 9.370 ;
      LAYER met4 ;
        RECT 11.595 9.050 11.915 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 8.620 11.915 8.940 ;
      LAYER met4 ;
        RECT 11.595 8.620 11.915 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 8.190 11.915 8.510 ;
      LAYER met4 ;
        RECT 11.595 8.190 11.915 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 7.760 11.915 8.080 ;
      LAYER met4 ;
        RECT 11.595 7.760 11.915 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 7.330 11.915 7.650 ;
      LAYER met4 ;
        RECT 11.595 7.330 11.915 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 6.900 11.915 7.220 ;
      LAYER met4 ;
        RECT 11.595 6.900 11.915 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 11.200 11.510 11.520 ;
      LAYER met4 ;
        RECT 11.190 11.200 11.510 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 10.770 11.510 11.090 ;
      LAYER met4 ;
        RECT 11.190 10.770 11.510 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 10.340 11.510 10.660 ;
      LAYER met4 ;
        RECT 11.190 10.340 11.510 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 9.910 11.510 10.230 ;
      LAYER met4 ;
        RECT 11.190 9.910 11.510 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 9.480 11.510 9.800 ;
      LAYER met4 ;
        RECT 11.190 9.480 11.510 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 9.050 11.510 9.370 ;
      LAYER met4 ;
        RECT 11.190 9.050 11.510 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 8.620 11.510 8.940 ;
      LAYER met4 ;
        RECT 11.190 8.620 11.510 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 8.190 11.510 8.510 ;
      LAYER met4 ;
        RECT 11.190 8.190 11.510 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 7.760 11.510 8.080 ;
      LAYER met4 ;
        RECT 11.190 7.760 11.510 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 7.330 11.510 7.650 ;
      LAYER met4 ;
        RECT 11.190 7.330 11.510 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 6.900 11.510 7.220 ;
      LAYER met4 ;
        RECT 11.190 6.900 11.510 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 11.200 11.105 11.520 ;
      LAYER met4 ;
        RECT 10.785 11.200 11.105 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 10.770 11.105 11.090 ;
      LAYER met4 ;
        RECT 10.785 10.770 11.105 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 10.340 11.105 10.660 ;
      LAYER met4 ;
        RECT 10.785 10.340 11.105 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 9.910 11.105 10.230 ;
      LAYER met4 ;
        RECT 10.785 9.910 11.105 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 9.480 11.105 9.800 ;
      LAYER met4 ;
        RECT 10.785 9.480 11.105 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 9.050 11.105 9.370 ;
      LAYER met4 ;
        RECT 10.785 9.050 11.105 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 8.620 11.105 8.940 ;
      LAYER met4 ;
        RECT 10.785 8.620 11.105 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 8.190 11.105 8.510 ;
      LAYER met4 ;
        RECT 10.785 8.190 11.105 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 7.760 11.105 8.080 ;
      LAYER met4 ;
        RECT 10.785 7.760 11.105 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 7.330 11.105 7.650 ;
      LAYER met4 ;
        RECT 10.785 7.330 11.105 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 6.900 11.105 7.220 ;
      LAYER met4 ;
        RECT 10.785 6.900 11.105 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 11.200 10.700 11.520 ;
      LAYER met4 ;
        RECT 10.380 11.200 10.700 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 10.770 10.700 11.090 ;
      LAYER met4 ;
        RECT 10.380 10.770 10.700 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 10.340 10.700 10.660 ;
      LAYER met4 ;
        RECT 10.380 10.340 10.700 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 9.910 10.700 10.230 ;
      LAYER met4 ;
        RECT 10.380 9.910 10.700 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 9.480 10.700 9.800 ;
      LAYER met4 ;
        RECT 10.380 9.480 10.700 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 9.050 10.700 9.370 ;
      LAYER met4 ;
        RECT 10.380 9.050 10.700 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 8.620 10.700 8.940 ;
      LAYER met4 ;
        RECT 10.380 8.620 10.700 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 8.190 10.700 8.510 ;
      LAYER met4 ;
        RECT 10.380 8.190 10.700 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 7.760 10.700 8.080 ;
      LAYER met4 ;
        RECT 10.380 7.760 10.700 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 7.330 10.700 7.650 ;
      LAYER met4 ;
        RECT 10.380 7.330 10.700 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 6.900 10.700 7.220 ;
      LAYER met4 ;
        RECT 10.380 6.900 10.700 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 11.200 10.295 11.520 ;
      LAYER met4 ;
        RECT 9.975 11.200 10.295 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 10.770 10.295 11.090 ;
      LAYER met4 ;
        RECT 9.975 10.770 10.295 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 10.340 10.295 10.660 ;
      LAYER met4 ;
        RECT 9.975 10.340 10.295 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 9.910 10.295 10.230 ;
      LAYER met4 ;
        RECT 9.975 9.910 10.295 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 9.480 10.295 9.800 ;
      LAYER met4 ;
        RECT 9.975 9.480 10.295 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 9.050 10.295 9.370 ;
      LAYER met4 ;
        RECT 9.975 9.050 10.295 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 8.620 10.295 8.940 ;
      LAYER met4 ;
        RECT 9.975 8.620 10.295 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 8.190 10.295 8.510 ;
      LAYER met4 ;
        RECT 9.975 8.190 10.295 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 7.760 10.295 8.080 ;
      LAYER met4 ;
        RECT 9.975 7.760 10.295 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 7.330 10.295 7.650 ;
      LAYER met4 ;
        RECT 9.975 7.330 10.295 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 6.900 10.295 7.220 ;
      LAYER met4 ;
        RECT 9.975 6.900 10.295 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 11.200 9.890 11.520 ;
      LAYER met4 ;
        RECT 9.570 11.200 9.890 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 10.770 9.890 11.090 ;
      LAYER met4 ;
        RECT 9.570 10.770 9.890 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 10.340 9.890 10.660 ;
      LAYER met4 ;
        RECT 9.570 10.340 9.890 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 9.910 9.890 10.230 ;
      LAYER met4 ;
        RECT 9.570 9.910 9.890 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 9.480 9.890 9.800 ;
      LAYER met4 ;
        RECT 9.570 9.480 9.890 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 9.050 9.890 9.370 ;
      LAYER met4 ;
        RECT 9.570 9.050 9.890 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 8.620 9.890 8.940 ;
      LAYER met4 ;
        RECT 9.570 8.620 9.890 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 8.190 9.890 8.510 ;
      LAYER met4 ;
        RECT 9.570 8.190 9.890 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 7.760 9.890 8.080 ;
      LAYER met4 ;
        RECT 9.570 7.760 9.890 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 7.330 9.890 7.650 ;
      LAYER met4 ;
        RECT 9.570 7.330 9.890 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 6.900 9.890 7.220 ;
      LAYER met4 ;
        RECT 9.570 6.900 9.890 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 11.200 9.485 11.520 ;
      LAYER met4 ;
        RECT 9.165 11.200 9.485 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 10.770 9.485 11.090 ;
      LAYER met4 ;
        RECT 9.165 10.770 9.485 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 10.340 9.485 10.660 ;
      LAYER met4 ;
        RECT 9.165 10.340 9.485 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 9.910 9.485 10.230 ;
      LAYER met4 ;
        RECT 9.165 9.910 9.485 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 9.480 9.485 9.800 ;
      LAYER met4 ;
        RECT 9.165 9.480 9.485 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 9.050 9.485 9.370 ;
      LAYER met4 ;
        RECT 9.165 9.050 9.485 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 8.620 9.485 8.940 ;
      LAYER met4 ;
        RECT 9.165 8.620 9.485 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 8.190 9.485 8.510 ;
      LAYER met4 ;
        RECT 9.165 8.190 9.485 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 7.760 9.485 8.080 ;
      LAYER met4 ;
        RECT 9.165 7.760 9.485 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 7.330 9.485 7.650 ;
      LAYER met4 ;
        RECT 9.165 7.330 9.485 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 6.900 9.485 7.220 ;
      LAYER met4 ;
        RECT 9.165 6.900 9.485 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 11.200 9.080 11.520 ;
      LAYER met4 ;
        RECT 8.760 11.200 9.080 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 10.770 9.080 11.090 ;
      LAYER met4 ;
        RECT 8.760 10.770 9.080 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 10.340 9.080 10.660 ;
      LAYER met4 ;
        RECT 8.760 10.340 9.080 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 9.910 9.080 10.230 ;
      LAYER met4 ;
        RECT 8.760 9.910 9.080 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 9.480 9.080 9.800 ;
      LAYER met4 ;
        RECT 8.760 9.480 9.080 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 9.050 9.080 9.370 ;
      LAYER met4 ;
        RECT 8.760 9.050 9.080 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 8.620 9.080 8.940 ;
      LAYER met4 ;
        RECT 8.760 8.620 9.080 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 8.190 9.080 8.510 ;
      LAYER met4 ;
        RECT 8.760 8.190 9.080 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 7.760 9.080 8.080 ;
      LAYER met4 ;
        RECT 8.760 7.760 9.080 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 7.330 9.080 7.650 ;
      LAYER met4 ;
        RECT 8.760 7.330 9.080 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 6.900 9.080 7.220 ;
      LAYER met4 ;
        RECT 8.760 6.900 9.080 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 11.200 8.675 11.520 ;
      LAYER met4 ;
        RECT 8.355 11.200 8.675 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 10.770 8.675 11.090 ;
      LAYER met4 ;
        RECT 8.355 10.770 8.675 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 10.340 8.675 10.660 ;
      LAYER met4 ;
        RECT 8.355 10.340 8.675 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 9.910 8.675 10.230 ;
      LAYER met4 ;
        RECT 8.355 9.910 8.675 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 9.480 8.675 9.800 ;
      LAYER met4 ;
        RECT 8.355 9.480 8.675 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 9.050 8.675 9.370 ;
      LAYER met4 ;
        RECT 8.355 9.050 8.675 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 8.620 8.675 8.940 ;
      LAYER met4 ;
        RECT 8.355 8.620 8.675 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 8.190 8.675 8.510 ;
      LAYER met4 ;
        RECT 8.355 8.190 8.675 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 7.760 8.675 8.080 ;
      LAYER met4 ;
        RECT 8.355 7.760 8.675 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 7.330 8.675 7.650 ;
      LAYER met4 ;
        RECT 8.355 7.330 8.675 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 6.900 8.675 7.220 ;
      LAYER met4 ;
        RECT 8.355 6.900 8.675 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 11.200 8.270 11.520 ;
      LAYER met4 ;
        RECT 7.950 11.200 8.270 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 10.770 8.270 11.090 ;
      LAYER met4 ;
        RECT 7.950 10.770 8.270 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 10.340 8.270 10.660 ;
      LAYER met4 ;
        RECT 7.950 10.340 8.270 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 9.910 8.270 10.230 ;
      LAYER met4 ;
        RECT 7.950 9.910 8.270 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 9.480 8.270 9.800 ;
      LAYER met4 ;
        RECT 7.950 9.480 8.270 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 9.050 8.270 9.370 ;
      LAYER met4 ;
        RECT 7.950 9.050 8.270 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 8.620 8.270 8.940 ;
      LAYER met4 ;
        RECT 7.950 8.620 8.270 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 8.190 8.270 8.510 ;
      LAYER met4 ;
        RECT 7.950 8.190 8.270 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 7.760 8.270 8.080 ;
      LAYER met4 ;
        RECT 7.950 7.760 8.270 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 7.330 8.270 7.650 ;
      LAYER met4 ;
        RECT 7.950 7.330 8.270 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 6.900 8.270 7.220 ;
      LAYER met4 ;
        RECT 7.950 6.900 8.270 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 11.200 7.865 11.520 ;
      LAYER met4 ;
        RECT 7.545 11.200 7.865 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 10.770 7.865 11.090 ;
      LAYER met4 ;
        RECT 7.545 10.770 7.865 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 10.340 7.865 10.660 ;
      LAYER met4 ;
        RECT 7.545 10.340 7.865 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 9.910 7.865 10.230 ;
      LAYER met4 ;
        RECT 7.545 9.910 7.865 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 9.480 7.865 9.800 ;
      LAYER met4 ;
        RECT 7.545 9.480 7.865 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 9.050 7.865 9.370 ;
      LAYER met4 ;
        RECT 7.545 9.050 7.865 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 8.620 7.865 8.940 ;
      LAYER met4 ;
        RECT 7.545 8.620 7.865 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 8.190 7.865 8.510 ;
      LAYER met4 ;
        RECT 7.545 8.190 7.865 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 7.760 7.865 8.080 ;
      LAYER met4 ;
        RECT 7.545 7.760 7.865 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 7.330 7.865 7.650 ;
      LAYER met4 ;
        RECT 7.545 7.330 7.865 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 6.900 7.865 7.220 ;
      LAYER met4 ;
        RECT 7.545 6.900 7.865 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 11.200 7.460 11.520 ;
      LAYER met4 ;
        RECT 7.140 11.200 7.460 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 10.770 7.460 11.090 ;
      LAYER met4 ;
        RECT 7.140 10.770 7.460 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 10.340 7.460 10.660 ;
      LAYER met4 ;
        RECT 7.140 10.340 7.460 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 9.910 7.460 10.230 ;
      LAYER met4 ;
        RECT 7.140 9.910 7.460 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 9.480 7.460 9.800 ;
      LAYER met4 ;
        RECT 7.140 9.480 7.460 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 9.050 7.460 9.370 ;
      LAYER met4 ;
        RECT 7.140 9.050 7.460 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 8.620 7.460 8.940 ;
      LAYER met4 ;
        RECT 7.140 8.620 7.460 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 8.190 7.460 8.510 ;
      LAYER met4 ;
        RECT 7.140 8.190 7.460 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 7.760 7.460 8.080 ;
      LAYER met4 ;
        RECT 7.140 7.760 7.460 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 7.330 7.460 7.650 ;
      LAYER met4 ;
        RECT 7.140 7.330 7.460 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 6.900 7.460 7.220 ;
      LAYER met4 ;
        RECT 7.140 6.900 7.460 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 11.200 7.055 11.520 ;
      LAYER met4 ;
        RECT 6.735 11.200 7.055 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 10.770 7.055 11.090 ;
      LAYER met4 ;
        RECT 6.735 10.770 7.055 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 10.340 7.055 10.660 ;
      LAYER met4 ;
        RECT 6.735 10.340 7.055 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 9.910 7.055 10.230 ;
      LAYER met4 ;
        RECT 6.735 9.910 7.055 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 9.480 7.055 9.800 ;
      LAYER met4 ;
        RECT 6.735 9.480 7.055 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 9.050 7.055 9.370 ;
      LAYER met4 ;
        RECT 6.735 9.050 7.055 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 8.620 7.055 8.940 ;
      LAYER met4 ;
        RECT 6.735 8.620 7.055 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 8.190 7.055 8.510 ;
      LAYER met4 ;
        RECT 6.735 8.190 7.055 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 7.760 7.055 8.080 ;
      LAYER met4 ;
        RECT 6.735 7.760 7.055 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 7.330 7.055 7.650 ;
      LAYER met4 ;
        RECT 6.735 7.330 7.055 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 6.900 7.055 7.220 ;
      LAYER met4 ;
        RECT 6.735 6.900 7.055 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 11.200 6.650 11.520 ;
      LAYER met4 ;
        RECT 6.330 11.200 6.650 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 10.770 6.650 11.090 ;
      LAYER met4 ;
        RECT 6.330 10.770 6.650 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 10.340 6.650 10.660 ;
      LAYER met4 ;
        RECT 6.330 10.340 6.650 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 9.910 6.650 10.230 ;
      LAYER met4 ;
        RECT 6.330 9.910 6.650 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 9.480 6.650 9.800 ;
      LAYER met4 ;
        RECT 6.330 9.480 6.650 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 9.050 6.650 9.370 ;
      LAYER met4 ;
        RECT 6.330 9.050 6.650 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 8.620 6.650 8.940 ;
      LAYER met4 ;
        RECT 6.330 8.620 6.650 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 8.190 6.650 8.510 ;
      LAYER met4 ;
        RECT 6.330 8.190 6.650 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 7.760 6.650 8.080 ;
      LAYER met4 ;
        RECT 6.330 7.760 6.650 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 7.330 6.650 7.650 ;
      LAYER met4 ;
        RECT 6.330 7.330 6.650 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 6.900 6.650 7.220 ;
      LAYER met4 ;
        RECT 6.330 6.900 6.650 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 11.200 6.245 11.520 ;
      LAYER met4 ;
        RECT 5.925 11.200 6.245 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 10.770 6.245 11.090 ;
      LAYER met4 ;
        RECT 5.925 10.770 6.245 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 10.340 6.245 10.660 ;
      LAYER met4 ;
        RECT 5.925 10.340 6.245 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 9.910 6.245 10.230 ;
      LAYER met4 ;
        RECT 5.925 9.910 6.245 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 9.480 6.245 9.800 ;
      LAYER met4 ;
        RECT 5.925 9.480 6.245 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 9.050 6.245 9.370 ;
      LAYER met4 ;
        RECT 5.925 9.050 6.245 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 8.620 6.245 8.940 ;
      LAYER met4 ;
        RECT 5.925 8.620 6.245 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 8.190 6.245 8.510 ;
      LAYER met4 ;
        RECT 5.925 8.190 6.245 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 7.760 6.245 8.080 ;
      LAYER met4 ;
        RECT 5.925 7.760 6.245 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 7.330 6.245 7.650 ;
      LAYER met4 ;
        RECT 5.925 7.330 6.245 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 6.900 6.245 7.220 ;
      LAYER met4 ;
        RECT 5.925 6.900 6.245 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 11.200 5.840 11.520 ;
      LAYER met4 ;
        RECT 5.520 11.200 5.840 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 10.770 5.840 11.090 ;
      LAYER met4 ;
        RECT 5.520 10.770 5.840 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 10.340 5.840 10.660 ;
      LAYER met4 ;
        RECT 5.520 10.340 5.840 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 9.910 5.840 10.230 ;
      LAYER met4 ;
        RECT 5.520 9.910 5.840 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 9.480 5.840 9.800 ;
      LAYER met4 ;
        RECT 5.520 9.480 5.840 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 9.050 5.840 9.370 ;
      LAYER met4 ;
        RECT 5.520 9.050 5.840 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 8.620 5.840 8.940 ;
      LAYER met4 ;
        RECT 5.520 8.620 5.840 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 8.190 5.840 8.510 ;
      LAYER met4 ;
        RECT 5.520 8.190 5.840 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 7.760 5.840 8.080 ;
      LAYER met4 ;
        RECT 5.520 7.760 5.840 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 7.330 5.840 7.650 ;
      LAYER met4 ;
        RECT 5.520 7.330 5.840 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 6.900 5.840 7.220 ;
      LAYER met4 ;
        RECT 5.520 6.900 5.840 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 11.200 5.435 11.520 ;
      LAYER met4 ;
        RECT 5.115 11.200 5.435 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 10.770 5.435 11.090 ;
      LAYER met4 ;
        RECT 5.115 10.770 5.435 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 10.340 5.435 10.660 ;
      LAYER met4 ;
        RECT 5.115 10.340 5.435 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 9.910 5.435 10.230 ;
      LAYER met4 ;
        RECT 5.115 9.910 5.435 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 9.480 5.435 9.800 ;
      LAYER met4 ;
        RECT 5.115 9.480 5.435 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 9.050 5.435 9.370 ;
      LAYER met4 ;
        RECT 5.115 9.050 5.435 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 8.620 5.435 8.940 ;
      LAYER met4 ;
        RECT 5.115 8.620 5.435 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 8.190 5.435 8.510 ;
      LAYER met4 ;
        RECT 5.115 8.190 5.435 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 7.760 5.435 8.080 ;
      LAYER met4 ;
        RECT 5.115 7.760 5.435 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 7.330 5.435 7.650 ;
      LAYER met4 ;
        RECT 5.115 7.330 5.435 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 6.900 5.435 7.220 ;
      LAYER met4 ;
        RECT 5.115 6.900 5.435 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 11.200 5.030 11.520 ;
      LAYER met4 ;
        RECT 4.710 11.200 5.030 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 10.770 5.030 11.090 ;
      LAYER met4 ;
        RECT 4.710 10.770 5.030 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 10.340 5.030 10.660 ;
      LAYER met4 ;
        RECT 4.710 10.340 5.030 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 9.910 5.030 10.230 ;
      LAYER met4 ;
        RECT 4.710 9.910 5.030 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 9.480 5.030 9.800 ;
      LAYER met4 ;
        RECT 4.710 9.480 5.030 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 9.050 5.030 9.370 ;
      LAYER met4 ;
        RECT 4.710 9.050 5.030 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 8.620 5.030 8.940 ;
      LAYER met4 ;
        RECT 4.710 8.620 5.030 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 8.190 5.030 8.510 ;
      LAYER met4 ;
        RECT 4.710 8.190 5.030 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 7.760 5.030 8.080 ;
      LAYER met4 ;
        RECT 4.710 7.760 5.030 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 7.330 5.030 7.650 ;
      LAYER met4 ;
        RECT 4.710 7.330 5.030 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 6.900 5.030 7.220 ;
      LAYER met4 ;
        RECT 4.710 6.900 5.030 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 11.200 4.625 11.520 ;
      LAYER met4 ;
        RECT 4.305 11.200 4.625 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 10.770 4.625 11.090 ;
      LAYER met4 ;
        RECT 4.305 10.770 4.625 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 10.340 4.625 10.660 ;
      LAYER met4 ;
        RECT 4.305 10.340 4.625 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 9.910 4.625 10.230 ;
      LAYER met4 ;
        RECT 4.305 9.910 4.625 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 9.480 4.625 9.800 ;
      LAYER met4 ;
        RECT 4.305 9.480 4.625 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 9.050 4.625 9.370 ;
      LAYER met4 ;
        RECT 4.305 9.050 4.625 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 8.620 4.625 8.940 ;
      LAYER met4 ;
        RECT 4.305 8.620 4.625 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 8.190 4.625 8.510 ;
      LAYER met4 ;
        RECT 4.305 8.190 4.625 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 7.760 4.625 8.080 ;
      LAYER met4 ;
        RECT 4.305 7.760 4.625 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 7.330 4.625 7.650 ;
      LAYER met4 ;
        RECT 4.305 7.330 4.625 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 6.900 4.625 7.220 ;
      LAYER met4 ;
        RECT 4.305 6.900 4.625 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 11.200 4.220 11.520 ;
      LAYER met4 ;
        RECT 3.900 11.200 4.220 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 10.770 4.220 11.090 ;
      LAYER met4 ;
        RECT 3.900 10.770 4.220 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 10.340 4.220 10.660 ;
      LAYER met4 ;
        RECT 3.900 10.340 4.220 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 9.910 4.220 10.230 ;
      LAYER met4 ;
        RECT 3.900 9.910 4.220 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 9.480 4.220 9.800 ;
      LAYER met4 ;
        RECT 3.900 9.480 4.220 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 9.050 4.220 9.370 ;
      LAYER met4 ;
        RECT 3.900 9.050 4.220 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 8.620 4.220 8.940 ;
      LAYER met4 ;
        RECT 3.900 8.620 4.220 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 8.190 4.220 8.510 ;
      LAYER met4 ;
        RECT 3.900 8.190 4.220 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 7.760 4.220 8.080 ;
      LAYER met4 ;
        RECT 3.900 7.760 4.220 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 7.330 4.220 7.650 ;
      LAYER met4 ;
        RECT 3.900 7.330 4.220 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 6.900 4.220 7.220 ;
      LAYER met4 ;
        RECT 3.900 6.900 4.220 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 11.200 3.815 11.520 ;
      LAYER met4 ;
        RECT 3.495 11.200 3.815 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 10.770 3.815 11.090 ;
      LAYER met4 ;
        RECT 3.495 10.770 3.815 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 10.340 3.815 10.660 ;
      LAYER met4 ;
        RECT 3.495 10.340 3.815 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 9.910 3.815 10.230 ;
      LAYER met4 ;
        RECT 3.495 9.910 3.815 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 9.480 3.815 9.800 ;
      LAYER met4 ;
        RECT 3.495 9.480 3.815 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 9.050 3.815 9.370 ;
      LAYER met4 ;
        RECT 3.495 9.050 3.815 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 8.620 3.815 8.940 ;
      LAYER met4 ;
        RECT 3.495 8.620 3.815 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 8.190 3.815 8.510 ;
      LAYER met4 ;
        RECT 3.495 8.190 3.815 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 7.760 3.815 8.080 ;
      LAYER met4 ;
        RECT 3.495 7.760 3.815 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 7.330 3.815 7.650 ;
      LAYER met4 ;
        RECT 3.495 7.330 3.815 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 6.900 3.815 7.220 ;
      LAYER met4 ;
        RECT 3.495 6.900 3.815 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 11.200 3.410 11.520 ;
      LAYER met4 ;
        RECT 3.090 11.200 3.410 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 10.770 3.410 11.090 ;
      LAYER met4 ;
        RECT 3.090 10.770 3.410 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 10.340 3.410 10.660 ;
      LAYER met4 ;
        RECT 3.090 10.340 3.410 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 9.910 3.410 10.230 ;
      LAYER met4 ;
        RECT 3.090 9.910 3.410 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 9.480 3.410 9.800 ;
      LAYER met4 ;
        RECT 3.090 9.480 3.410 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 9.050 3.410 9.370 ;
      LAYER met4 ;
        RECT 3.090 9.050 3.410 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 8.620 3.410 8.940 ;
      LAYER met4 ;
        RECT 3.090 8.620 3.410 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 8.190 3.410 8.510 ;
      LAYER met4 ;
        RECT 3.090 8.190 3.410 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 7.760 3.410 8.080 ;
      LAYER met4 ;
        RECT 3.090 7.760 3.410 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 7.330 3.410 7.650 ;
      LAYER met4 ;
        RECT 3.090 7.330 3.410 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 6.900 3.410 7.220 ;
      LAYER met4 ;
        RECT 3.090 6.900 3.410 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 11.200 3.000 11.520 ;
      LAYER met4 ;
        RECT 2.680 11.200 3.000 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 10.770 3.000 11.090 ;
      LAYER met4 ;
        RECT 2.680 10.770 3.000 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 10.340 3.000 10.660 ;
      LAYER met4 ;
        RECT 2.680 10.340 3.000 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 9.910 3.000 10.230 ;
      LAYER met4 ;
        RECT 2.680 9.910 3.000 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 9.480 3.000 9.800 ;
      LAYER met4 ;
        RECT 2.680 9.480 3.000 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 9.050 3.000 9.370 ;
      LAYER met4 ;
        RECT 2.680 9.050 3.000 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 8.620 3.000 8.940 ;
      LAYER met4 ;
        RECT 2.680 8.620 3.000 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 8.190 3.000 8.510 ;
      LAYER met4 ;
        RECT 2.680 8.190 3.000 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 7.760 3.000 8.080 ;
      LAYER met4 ;
        RECT 2.680 7.760 3.000 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 7.330 3.000 7.650 ;
      LAYER met4 ;
        RECT 2.680 7.330 3.000 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 6.900 3.000 7.220 ;
      LAYER met4 ;
        RECT 2.680 6.900 3.000 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 11.200 2.590 11.520 ;
      LAYER met4 ;
        RECT 2.270 11.200 2.590 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 10.770 2.590 11.090 ;
      LAYER met4 ;
        RECT 2.270 10.770 2.590 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 10.340 2.590 10.660 ;
      LAYER met4 ;
        RECT 2.270 10.340 2.590 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 9.910 2.590 10.230 ;
      LAYER met4 ;
        RECT 2.270 9.910 2.590 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 9.480 2.590 9.800 ;
      LAYER met4 ;
        RECT 2.270 9.480 2.590 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 9.050 2.590 9.370 ;
      LAYER met4 ;
        RECT 2.270 9.050 2.590 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 8.620 2.590 8.940 ;
      LAYER met4 ;
        RECT 2.270 8.620 2.590 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 8.190 2.590 8.510 ;
      LAYER met4 ;
        RECT 2.270 8.190 2.590 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 7.760 2.590 8.080 ;
      LAYER met4 ;
        RECT 2.270 7.760 2.590 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 7.330 2.590 7.650 ;
      LAYER met4 ;
        RECT 2.270 7.330 2.590 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 6.900 2.590 7.220 ;
      LAYER met4 ;
        RECT 2.270 6.900 2.590 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 11.200 2.180 11.520 ;
      LAYER met4 ;
        RECT 1.860 11.200 2.180 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 10.770 2.180 11.090 ;
      LAYER met4 ;
        RECT 1.860 10.770 2.180 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 10.340 2.180 10.660 ;
      LAYER met4 ;
        RECT 1.860 10.340 2.180 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 9.910 2.180 10.230 ;
      LAYER met4 ;
        RECT 1.860 9.910 2.180 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 9.480 2.180 9.800 ;
      LAYER met4 ;
        RECT 1.860 9.480 2.180 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 9.050 2.180 9.370 ;
      LAYER met4 ;
        RECT 1.860 9.050 2.180 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 8.620 2.180 8.940 ;
      LAYER met4 ;
        RECT 1.860 8.620 2.180 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 8.190 2.180 8.510 ;
      LAYER met4 ;
        RECT 1.860 8.190 2.180 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 7.760 2.180 8.080 ;
      LAYER met4 ;
        RECT 1.860 7.760 2.180 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 7.330 2.180 7.650 ;
      LAYER met4 ;
        RECT 1.860 7.330 2.180 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 6.900 2.180 7.220 ;
      LAYER met4 ;
        RECT 1.860 6.900 2.180 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 11.200 1.770 11.520 ;
      LAYER met4 ;
        RECT 1.450 11.200 1.770 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 10.770 1.770 11.090 ;
      LAYER met4 ;
        RECT 1.450 10.770 1.770 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 10.340 1.770 10.660 ;
      LAYER met4 ;
        RECT 1.450 10.340 1.770 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 9.910 1.770 10.230 ;
      LAYER met4 ;
        RECT 1.450 9.910 1.770 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 9.480 1.770 9.800 ;
      LAYER met4 ;
        RECT 1.450 9.480 1.770 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 9.050 1.770 9.370 ;
      LAYER met4 ;
        RECT 1.450 9.050 1.770 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 8.620 1.770 8.940 ;
      LAYER met4 ;
        RECT 1.450 8.620 1.770 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 8.190 1.770 8.510 ;
      LAYER met4 ;
        RECT 1.450 8.190 1.770 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 7.760 1.770 8.080 ;
      LAYER met4 ;
        RECT 1.450 7.760 1.770 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 7.330 1.770 7.650 ;
      LAYER met4 ;
        RECT 1.450 7.330 1.770 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 6.900 1.770 7.220 ;
      LAYER met4 ;
        RECT 1.450 6.900 1.770 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 11.200 1.360 11.520 ;
      LAYER met4 ;
        RECT 1.270 11.200 1.360 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 10.770 1.360 11.090 ;
      LAYER met4 ;
        RECT 1.270 10.770 1.360 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 10.340 1.360 10.660 ;
      LAYER met4 ;
        RECT 1.270 10.340 1.360 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 9.910 1.360 10.230 ;
      LAYER met4 ;
        RECT 1.270 9.910 1.360 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 9.480 1.360 9.800 ;
      LAYER met4 ;
        RECT 1.270 9.480 1.360 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 9.050 1.360 9.370 ;
      LAYER met4 ;
        RECT 1.270 9.050 1.360 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 8.620 1.360 8.940 ;
      LAYER met4 ;
        RECT 1.270 8.620 1.360 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 8.190 1.360 8.510 ;
      LAYER met4 ;
        RECT 1.270 8.190 1.360 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 7.760 1.360 8.080 ;
      LAYER met4 ;
        RECT 1.270 7.760 1.360 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 7.330 1.360 7.650 ;
      LAYER met4 ;
        RECT 1.270 7.330 1.360 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 6.900 1.360 7.220 ;
      LAYER met4 ;
        RECT 1.270 6.900 1.360 7.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 11.200 0.950 11.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 10.770 0.950 11.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 10.340 0.950 10.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 9.910 0.950 10.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 9.480 0.950 9.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 9.050 0.950 9.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 8.620 0.950 8.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 8.190 0.950 8.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 7.760 0.950 8.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 7.330 0.950 7.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 6.900 0.950 7.220 ;
    END
  END VCCD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
  END VDDA
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
  END VSWITCH
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
  END VSSD
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.600 6.890 24.500 11.530 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 94.585 75.000 172.185 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__overlay_vccd_lvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vdda_hvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vdda_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
  END VSSA
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
  END VSSIO_Q
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
  END VSSD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 14.940 74.290 18.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 18.100 74.200 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 17.660 74.200 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 17.220 74.200 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 16.780 74.200 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 16.340 74.200 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 15.900 74.200 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 15.460 74.200 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 15.020 74.200 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 18.100 73.795 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 17.660 73.795 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 17.220 73.795 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 16.780 73.795 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 16.340 73.795 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 15.900 73.795 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 15.460 73.795 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 15.020 73.795 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 18.100 73.390 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 17.660 73.390 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 17.220 73.390 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 16.780 73.390 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 16.340 73.390 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 15.900 73.390 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 15.460 73.390 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 15.020 73.390 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 18.100 72.985 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 17.660 72.985 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 17.220 72.985 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 16.780 72.985 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 16.340 72.985 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 15.900 72.985 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 15.460 72.985 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 15.020 72.985 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 18.100 72.580 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 17.660 72.580 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 17.220 72.580 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 16.780 72.580 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 16.340 72.580 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 15.900 72.580 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 15.460 72.580 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 15.020 72.580 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 18.100 72.175 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 17.660 72.175 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 17.220 72.175 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 16.780 72.175 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 16.340 72.175 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 15.900 72.175 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 15.460 72.175 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 15.020 72.175 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 18.100 71.770 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 17.660 71.770 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 17.220 71.770 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 16.780 71.770 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 16.340 71.770 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 15.900 71.770 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 15.460 71.770 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 15.020 71.770 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 18.100 71.365 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 17.660 71.365 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 17.220 71.365 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 16.780 71.365 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 16.340 71.365 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 15.900 71.365 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 15.460 71.365 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 15.020 71.365 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 18.100 70.960 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 17.660 70.960 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 17.220 70.960 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 16.780 70.960 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 16.340 70.960 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 15.900 70.960 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 15.460 70.960 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 15.020 70.960 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 18.100 70.555 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 17.660 70.555 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 17.220 70.555 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 16.780 70.555 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 16.340 70.555 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 15.900 70.555 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 15.460 70.555 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 15.020 70.555 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 18.100 70.150 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 17.660 70.150 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 17.220 70.150 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 16.780 70.150 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 16.340 70.150 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 15.900 70.150 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 15.460 70.150 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 15.020 70.150 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 18.100 69.745 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 17.660 69.745 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 17.220 69.745 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 16.780 69.745 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 16.340 69.745 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 15.900 69.745 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 15.460 69.745 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 15.020 69.745 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 18.100 69.340 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 17.660 69.340 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 17.220 69.340 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 16.780 69.340 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 16.340 69.340 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 15.900 69.340 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 15.460 69.340 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 15.020 69.340 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 18.100 68.935 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 17.660 68.935 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 17.220 68.935 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 16.780 68.935 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 16.340 68.935 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 15.900 68.935 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 15.460 68.935 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 15.020 68.935 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 18.100 68.530 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 17.660 68.530 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 17.220 68.530 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 16.780 68.530 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 16.340 68.530 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 15.900 68.530 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 15.460 68.530 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 15.020 68.530 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 18.100 68.125 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 17.660 68.125 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 17.220 68.125 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 16.780 68.125 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 16.340 68.125 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 15.900 68.125 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 15.460 68.125 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 15.020 68.125 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 18.100 67.720 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 17.660 67.720 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 17.220 67.720 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 16.780 67.720 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 16.340 67.720 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 15.900 67.720 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 15.460 67.720 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 15.020 67.720 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 18.100 67.315 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 17.660 67.315 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 17.220 67.315 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 16.780 67.315 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 16.340 67.315 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 15.900 67.315 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 15.460 67.315 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 15.020 67.315 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 18.100 66.910 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 17.660 66.910 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 17.220 66.910 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 16.780 66.910 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 16.340 66.910 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 15.900 66.910 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 15.460 66.910 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 15.020 66.910 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 18.100 66.505 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 17.660 66.505 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 17.220 66.505 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 16.780 66.505 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 16.340 66.505 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 15.900 66.505 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 15.460 66.505 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 15.020 66.505 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 18.100 66.100 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 17.660 66.100 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 17.220 66.100 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 16.780 66.100 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 16.340 66.100 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 15.900 66.100 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 15.460 66.100 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 15.020 66.100 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 18.100 65.695 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 17.660 65.695 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 17.220 65.695 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 16.780 65.695 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 16.340 65.695 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 15.900 65.695 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 15.460 65.695 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 15.020 65.695 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 18.100 65.290 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 17.660 65.290 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 17.220 65.290 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 16.780 65.290 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 16.340 65.290 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 15.900 65.290 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 15.460 65.290 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 15.020 65.290 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 18.100 64.885 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 17.660 64.885 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 17.220 64.885 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 16.780 64.885 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 16.340 64.885 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 15.900 64.885 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 15.460 64.885 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 15.020 64.885 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 18.100 64.480 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 17.660 64.480 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 17.220 64.480 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 16.780 64.480 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 16.340 64.480 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 15.900 64.480 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 15.460 64.480 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 15.020 64.480 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 18.100 64.075 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 17.660 64.075 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 17.220 64.075 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 16.780 64.075 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 16.340 64.075 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 15.900 64.075 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 15.460 64.075 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 15.020 64.075 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 18.100 63.670 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 17.660 63.670 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 17.220 63.670 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 16.780 63.670 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 16.340 63.670 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 15.900 63.670 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 15.460 63.670 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 15.020 63.670 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 18.100 63.265 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 17.660 63.265 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 17.220 63.265 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 16.780 63.265 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 16.340 63.265 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 15.900 63.265 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 15.460 63.265 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 15.020 63.265 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 18.100 62.860 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 17.660 62.860 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 17.220 62.860 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 16.780 62.860 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 16.340 62.860 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 15.900 62.860 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 15.460 62.860 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 15.020 62.860 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 18.100 62.455 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 17.660 62.455 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 17.220 62.455 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 16.780 62.455 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 16.340 62.455 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 15.900 62.455 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 15.460 62.455 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 15.020 62.455 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 18.100 62.050 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 17.660 62.050 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 17.220 62.050 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 16.780 62.050 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 16.340 62.050 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 15.900 62.050 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 15.460 62.050 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 15.020 62.050 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 18.100 61.645 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 17.660 61.645 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 17.220 61.645 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 16.780 61.645 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 16.340 61.645 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 15.900 61.645 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 15.460 61.645 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 15.020 61.645 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 18.100 61.240 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 17.660 61.240 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 17.220 61.240 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 16.780 61.240 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 16.340 61.240 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 15.900 61.240 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 15.460 61.240 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 15.020 61.240 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 18.100 60.835 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 17.660 60.835 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 17.220 60.835 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 16.780 60.835 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 16.340 60.835 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 15.900 60.835 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 15.460 60.835 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 15.020 60.835 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 18.100 60.430 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 17.660 60.430 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 17.220 60.430 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 16.780 60.430 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 16.340 60.430 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 15.900 60.430 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 15.460 60.430 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 15.020 60.430 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 18.100 60.025 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 17.660 60.025 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 17.220 60.025 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 16.780 60.025 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 16.340 60.025 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 15.900 60.025 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 15.460 60.025 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 15.020 60.025 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 18.100 59.620 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 17.660 59.620 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 17.220 59.620 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 16.780 59.620 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 16.340 59.620 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 15.900 59.620 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 15.460 59.620 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 15.020 59.620 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 18.100 59.215 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 17.660 59.215 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 17.220 59.215 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 16.780 59.215 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 16.340 59.215 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 15.900 59.215 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 15.460 59.215 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 15.020 59.215 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 18.100 58.810 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 17.660 58.810 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 17.220 58.810 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 16.780 58.810 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 16.340 58.810 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 15.900 58.810 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 15.460 58.810 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 15.020 58.810 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 18.100 58.405 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 17.660 58.405 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 17.220 58.405 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 16.780 58.405 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 16.340 58.405 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 15.900 58.405 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 15.460 58.405 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 15.020 58.405 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 18.100 58.000 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 17.660 58.000 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 17.220 58.000 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 16.780 58.000 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 16.340 58.000 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 15.900 58.000 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 15.460 58.000 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 15.020 58.000 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 18.100 57.595 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 17.660 57.595 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 17.220 57.595 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 16.780 57.595 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 16.340 57.595 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 15.900 57.595 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 15.460 57.595 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 15.020 57.595 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 18.100 57.190 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 17.660 57.190 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 17.220 57.190 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 16.780 57.190 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 16.340 57.190 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 15.900 57.190 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 15.460 57.190 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 15.020 57.190 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 18.100 56.785 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 17.660 56.785 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 17.220 56.785 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 16.780 56.785 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 16.340 56.785 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 15.900 56.785 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 15.460 56.785 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 15.020 56.785 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 18.100 56.380 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 17.660 56.380 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 17.220 56.380 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 16.780 56.380 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 16.340 56.380 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 15.900 56.380 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 15.460 56.380 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 15.020 56.380 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 18.100 55.975 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 17.660 55.975 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 17.220 55.975 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 16.780 55.975 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 16.340 55.975 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 15.900 55.975 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 15.460 55.975 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 15.020 55.975 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 18.100 55.570 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 17.660 55.570 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 17.220 55.570 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 16.780 55.570 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 16.340 55.570 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 15.900 55.570 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 15.460 55.570 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 15.020 55.570 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 18.100 55.165 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 17.660 55.165 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 17.220 55.165 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 16.780 55.165 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 16.340 55.165 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 15.900 55.165 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 15.460 55.165 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 15.020 55.165 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 18.100 54.760 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 17.660 54.760 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 17.220 54.760 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 16.780 54.760 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 16.340 54.760 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 15.900 54.760 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 15.460 54.760 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 15.020 54.760 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 18.100 54.355 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 17.660 54.355 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 17.220 54.355 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 16.780 54.355 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 16.340 54.355 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 15.900 54.355 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 15.460 54.355 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 15.020 54.355 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 18.100 53.950 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 17.660 53.950 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 17.220 53.950 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 16.780 53.950 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 16.340 53.950 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 15.900 53.950 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 15.460 53.950 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 15.020 53.950 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 18.100 53.545 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 17.660 53.545 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 17.220 53.545 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 16.780 53.545 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 16.340 53.545 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 15.900 53.545 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 15.460 53.545 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 15.020 53.545 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 18.100 53.140 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 17.660 53.140 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 17.220 53.140 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 16.780 53.140 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 16.340 53.140 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 15.900 53.140 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 15.460 53.140 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 15.020 53.140 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 18.100 52.730 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 17.660 52.730 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 17.220 52.730 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 16.780 52.730 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 16.340 52.730 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 15.900 52.730 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 15.460 52.730 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 15.020 52.730 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 18.100 52.320 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 17.660 52.320 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 17.220 52.320 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 16.780 52.320 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 16.340 52.320 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 15.900 52.320 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 15.460 52.320 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 15.020 52.320 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 18.100 51.910 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 17.660 51.910 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 17.220 51.910 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 16.780 51.910 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 16.340 51.910 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 15.900 51.910 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 15.460 51.910 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 15.020 51.910 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 18.100 51.500 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 17.660 51.500 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 17.220 51.500 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 16.780 51.500 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 16.340 51.500 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 15.900 51.500 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 15.460 51.500 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 15.020 51.500 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 18.100 51.090 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 17.660 51.090 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 17.220 51.090 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 16.780 51.090 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 16.340 51.090 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 15.900 51.090 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 15.460 51.090 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 15.020 51.090 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 18.100 50.680 18.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 17.660 50.680 17.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 17.220 50.680 17.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 16.780 50.680 16.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 16.340 50.680 16.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 15.900 50.680 16.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 15.460 50.680 15.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 15.020 50.680 15.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 18.040 24.365 18.360 ;
      LAYER met4 ;
        RECT 24.045 18.040 24.365 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 17.600 24.365 17.920 ;
      LAYER met4 ;
        RECT 24.045 17.600 24.365 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 17.160 24.365 17.480 ;
      LAYER met4 ;
        RECT 24.045 17.160 24.365 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 16.720 24.365 17.040 ;
      LAYER met4 ;
        RECT 24.045 16.720 24.365 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 16.280 24.365 16.600 ;
      LAYER met4 ;
        RECT 24.045 16.280 24.365 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 15.840 24.365 16.160 ;
      LAYER met4 ;
        RECT 24.045 15.840 24.365 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 15.400 24.365 15.720 ;
      LAYER met4 ;
        RECT 24.045 15.400 24.365 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 14.960 24.365 15.280 ;
      LAYER met4 ;
        RECT 24.045 14.960 24.365 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 18.040 23.960 18.360 ;
      LAYER met4 ;
        RECT 23.640 18.040 23.960 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 17.600 23.960 17.920 ;
      LAYER met4 ;
        RECT 23.640 17.600 23.960 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 17.160 23.960 17.480 ;
      LAYER met4 ;
        RECT 23.640 17.160 23.960 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 16.720 23.960 17.040 ;
      LAYER met4 ;
        RECT 23.640 16.720 23.960 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 16.280 23.960 16.600 ;
      LAYER met4 ;
        RECT 23.640 16.280 23.960 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 15.840 23.960 16.160 ;
      LAYER met4 ;
        RECT 23.640 15.840 23.960 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 15.400 23.960 15.720 ;
      LAYER met4 ;
        RECT 23.640 15.400 23.960 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 14.960 23.960 15.280 ;
      LAYER met4 ;
        RECT 23.640 14.960 23.960 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 18.040 23.555 18.360 ;
      LAYER met4 ;
        RECT 23.235 18.040 23.555 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 17.600 23.555 17.920 ;
      LAYER met4 ;
        RECT 23.235 17.600 23.555 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 17.160 23.555 17.480 ;
      LAYER met4 ;
        RECT 23.235 17.160 23.555 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 16.720 23.555 17.040 ;
      LAYER met4 ;
        RECT 23.235 16.720 23.555 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 16.280 23.555 16.600 ;
      LAYER met4 ;
        RECT 23.235 16.280 23.555 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 15.840 23.555 16.160 ;
      LAYER met4 ;
        RECT 23.235 15.840 23.555 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 15.400 23.555 15.720 ;
      LAYER met4 ;
        RECT 23.235 15.400 23.555 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 14.960 23.555 15.280 ;
      LAYER met4 ;
        RECT 23.235 14.960 23.555 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 18.040 23.150 18.360 ;
      LAYER met4 ;
        RECT 22.830 18.040 23.150 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 17.600 23.150 17.920 ;
      LAYER met4 ;
        RECT 22.830 17.600 23.150 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 17.160 23.150 17.480 ;
      LAYER met4 ;
        RECT 22.830 17.160 23.150 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 16.720 23.150 17.040 ;
      LAYER met4 ;
        RECT 22.830 16.720 23.150 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 16.280 23.150 16.600 ;
      LAYER met4 ;
        RECT 22.830 16.280 23.150 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 15.840 23.150 16.160 ;
      LAYER met4 ;
        RECT 22.830 15.840 23.150 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 15.400 23.150 15.720 ;
      LAYER met4 ;
        RECT 22.830 15.400 23.150 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 14.960 23.150 15.280 ;
      LAYER met4 ;
        RECT 22.830 14.960 23.150 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 18.040 22.745 18.360 ;
      LAYER met4 ;
        RECT 22.425 18.040 22.745 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 17.600 22.745 17.920 ;
      LAYER met4 ;
        RECT 22.425 17.600 22.745 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 17.160 22.745 17.480 ;
      LAYER met4 ;
        RECT 22.425 17.160 22.745 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 16.720 22.745 17.040 ;
      LAYER met4 ;
        RECT 22.425 16.720 22.745 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 16.280 22.745 16.600 ;
      LAYER met4 ;
        RECT 22.425 16.280 22.745 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 15.840 22.745 16.160 ;
      LAYER met4 ;
        RECT 22.425 15.840 22.745 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 15.400 22.745 15.720 ;
      LAYER met4 ;
        RECT 22.425 15.400 22.745 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 14.960 22.745 15.280 ;
      LAYER met4 ;
        RECT 22.425 14.960 22.745 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 18.040 22.340 18.360 ;
      LAYER met4 ;
        RECT 22.020 18.040 22.340 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 17.600 22.340 17.920 ;
      LAYER met4 ;
        RECT 22.020 17.600 22.340 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 17.160 22.340 17.480 ;
      LAYER met4 ;
        RECT 22.020 17.160 22.340 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 16.720 22.340 17.040 ;
      LAYER met4 ;
        RECT 22.020 16.720 22.340 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 16.280 22.340 16.600 ;
      LAYER met4 ;
        RECT 22.020 16.280 22.340 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 15.840 22.340 16.160 ;
      LAYER met4 ;
        RECT 22.020 15.840 22.340 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 15.400 22.340 15.720 ;
      LAYER met4 ;
        RECT 22.020 15.400 22.340 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 14.960 22.340 15.280 ;
      LAYER met4 ;
        RECT 22.020 14.960 22.340 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 18.040 21.935 18.360 ;
      LAYER met4 ;
        RECT 21.615 18.040 21.935 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 17.600 21.935 17.920 ;
      LAYER met4 ;
        RECT 21.615 17.600 21.935 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 17.160 21.935 17.480 ;
      LAYER met4 ;
        RECT 21.615 17.160 21.935 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 16.720 21.935 17.040 ;
      LAYER met4 ;
        RECT 21.615 16.720 21.935 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 16.280 21.935 16.600 ;
      LAYER met4 ;
        RECT 21.615 16.280 21.935 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 15.840 21.935 16.160 ;
      LAYER met4 ;
        RECT 21.615 15.840 21.935 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 15.400 21.935 15.720 ;
      LAYER met4 ;
        RECT 21.615 15.400 21.935 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 14.960 21.935 15.280 ;
      LAYER met4 ;
        RECT 21.615 14.960 21.935 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 18.040 21.530 18.360 ;
      LAYER met4 ;
        RECT 21.210 18.040 21.530 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 17.600 21.530 17.920 ;
      LAYER met4 ;
        RECT 21.210 17.600 21.530 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 17.160 21.530 17.480 ;
      LAYER met4 ;
        RECT 21.210 17.160 21.530 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 16.720 21.530 17.040 ;
      LAYER met4 ;
        RECT 21.210 16.720 21.530 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 16.280 21.530 16.600 ;
      LAYER met4 ;
        RECT 21.210 16.280 21.530 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 15.840 21.530 16.160 ;
      LAYER met4 ;
        RECT 21.210 15.840 21.530 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 15.400 21.530 15.720 ;
      LAYER met4 ;
        RECT 21.210 15.400 21.530 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 14.960 21.530 15.280 ;
      LAYER met4 ;
        RECT 21.210 14.960 21.530 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 18.040 21.125 18.360 ;
      LAYER met4 ;
        RECT 20.805 18.040 21.125 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 17.600 21.125 17.920 ;
      LAYER met4 ;
        RECT 20.805 17.600 21.125 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 17.160 21.125 17.480 ;
      LAYER met4 ;
        RECT 20.805 17.160 21.125 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 16.720 21.125 17.040 ;
      LAYER met4 ;
        RECT 20.805 16.720 21.125 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 16.280 21.125 16.600 ;
      LAYER met4 ;
        RECT 20.805 16.280 21.125 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 15.840 21.125 16.160 ;
      LAYER met4 ;
        RECT 20.805 15.840 21.125 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 15.400 21.125 15.720 ;
      LAYER met4 ;
        RECT 20.805 15.400 21.125 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 14.960 21.125 15.280 ;
      LAYER met4 ;
        RECT 20.805 14.960 21.125 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 18.040 20.720 18.360 ;
      LAYER met4 ;
        RECT 20.400 18.040 20.720 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 17.600 20.720 17.920 ;
      LAYER met4 ;
        RECT 20.400 17.600 20.720 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 17.160 20.720 17.480 ;
      LAYER met4 ;
        RECT 20.400 17.160 20.720 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 16.720 20.720 17.040 ;
      LAYER met4 ;
        RECT 20.400 16.720 20.720 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 16.280 20.720 16.600 ;
      LAYER met4 ;
        RECT 20.400 16.280 20.720 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 15.840 20.720 16.160 ;
      LAYER met4 ;
        RECT 20.400 15.840 20.720 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 15.400 20.720 15.720 ;
      LAYER met4 ;
        RECT 20.400 15.400 20.720 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 14.960 20.720 15.280 ;
      LAYER met4 ;
        RECT 20.400 14.960 20.720 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 18.040 20.315 18.360 ;
      LAYER met4 ;
        RECT 19.995 18.040 20.315 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 17.600 20.315 17.920 ;
      LAYER met4 ;
        RECT 19.995 17.600 20.315 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 17.160 20.315 17.480 ;
      LAYER met4 ;
        RECT 19.995 17.160 20.315 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 16.720 20.315 17.040 ;
      LAYER met4 ;
        RECT 19.995 16.720 20.315 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 16.280 20.315 16.600 ;
      LAYER met4 ;
        RECT 19.995 16.280 20.315 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 15.840 20.315 16.160 ;
      LAYER met4 ;
        RECT 19.995 15.840 20.315 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 15.400 20.315 15.720 ;
      LAYER met4 ;
        RECT 19.995 15.400 20.315 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 14.960 20.315 15.280 ;
      LAYER met4 ;
        RECT 19.995 14.960 20.315 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 18.040 19.910 18.360 ;
      LAYER met4 ;
        RECT 19.590 18.040 19.910 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 17.600 19.910 17.920 ;
      LAYER met4 ;
        RECT 19.590 17.600 19.910 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 17.160 19.910 17.480 ;
      LAYER met4 ;
        RECT 19.590 17.160 19.910 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 16.720 19.910 17.040 ;
      LAYER met4 ;
        RECT 19.590 16.720 19.910 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 16.280 19.910 16.600 ;
      LAYER met4 ;
        RECT 19.590 16.280 19.910 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 15.840 19.910 16.160 ;
      LAYER met4 ;
        RECT 19.590 15.840 19.910 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 15.400 19.910 15.720 ;
      LAYER met4 ;
        RECT 19.590 15.400 19.910 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 14.960 19.910 15.280 ;
      LAYER met4 ;
        RECT 19.590 14.960 19.910 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 18.040 19.505 18.360 ;
      LAYER met4 ;
        RECT 19.185 18.040 19.505 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 17.600 19.505 17.920 ;
      LAYER met4 ;
        RECT 19.185 17.600 19.505 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 17.160 19.505 17.480 ;
      LAYER met4 ;
        RECT 19.185 17.160 19.505 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 16.720 19.505 17.040 ;
      LAYER met4 ;
        RECT 19.185 16.720 19.505 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 16.280 19.505 16.600 ;
      LAYER met4 ;
        RECT 19.185 16.280 19.505 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 15.840 19.505 16.160 ;
      LAYER met4 ;
        RECT 19.185 15.840 19.505 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 15.400 19.505 15.720 ;
      LAYER met4 ;
        RECT 19.185 15.400 19.505 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 14.960 19.505 15.280 ;
      LAYER met4 ;
        RECT 19.185 14.960 19.505 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 18.040 19.100 18.360 ;
      LAYER met4 ;
        RECT 18.780 18.040 19.100 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 17.600 19.100 17.920 ;
      LAYER met4 ;
        RECT 18.780 17.600 19.100 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 17.160 19.100 17.480 ;
      LAYER met4 ;
        RECT 18.780 17.160 19.100 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 16.720 19.100 17.040 ;
      LAYER met4 ;
        RECT 18.780 16.720 19.100 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 16.280 19.100 16.600 ;
      LAYER met4 ;
        RECT 18.780 16.280 19.100 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 15.840 19.100 16.160 ;
      LAYER met4 ;
        RECT 18.780 15.840 19.100 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 15.400 19.100 15.720 ;
      LAYER met4 ;
        RECT 18.780 15.400 19.100 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 14.960 19.100 15.280 ;
      LAYER met4 ;
        RECT 18.780 14.960 19.100 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 18.040 18.695 18.360 ;
      LAYER met4 ;
        RECT 18.375 18.040 18.695 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 17.600 18.695 17.920 ;
      LAYER met4 ;
        RECT 18.375 17.600 18.695 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 17.160 18.695 17.480 ;
      LAYER met4 ;
        RECT 18.375 17.160 18.695 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 16.720 18.695 17.040 ;
      LAYER met4 ;
        RECT 18.375 16.720 18.695 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 16.280 18.695 16.600 ;
      LAYER met4 ;
        RECT 18.375 16.280 18.695 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 15.840 18.695 16.160 ;
      LAYER met4 ;
        RECT 18.375 15.840 18.695 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 15.400 18.695 15.720 ;
      LAYER met4 ;
        RECT 18.375 15.400 18.695 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 14.960 18.695 15.280 ;
      LAYER met4 ;
        RECT 18.375 14.960 18.695 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 18.040 18.290 18.360 ;
      LAYER met4 ;
        RECT 17.970 18.040 18.290 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 17.600 18.290 17.920 ;
      LAYER met4 ;
        RECT 17.970 17.600 18.290 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 17.160 18.290 17.480 ;
      LAYER met4 ;
        RECT 17.970 17.160 18.290 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 16.720 18.290 17.040 ;
      LAYER met4 ;
        RECT 17.970 16.720 18.290 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 16.280 18.290 16.600 ;
      LAYER met4 ;
        RECT 17.970 16.280 18.290 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 15.840 18.290 16.160 ;
      LAYER met4 ;
        RECT 17.970 15.840 18.290 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 15.400 18.290 15.720 ;
      LAYER met4 ;
        RECT 17.970 15.400 18.290 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 14.960 18.290 15.280 ;
      LAYER met4 ;
        RECT 17.970 14.960 18.290 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 18.040 17.885 18.360 ;
      LAYER met4 ;
        RECT 17.565 18.040 17.885 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 17.600 17.885 17.920 ;
      LAYER met4 ;
        RECT 17.565 17.600 17.885 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 17.160 17.885 17.480 ;
      LAYER met4 ;
        RECT 17.565 17.160 17.885 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 16.720 17.885 17.040 ;
      LAYER met4 ;
        RECT 17.565 16.720 17.885 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 16.280 17.885 16.600 ;
      LAYER met4 ;
        RECT 17.565 16.280 17.885 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 15.840 17.885 16.160 ;
      LAYER met4 ;
        RECT 17.565 15.840 17.885 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 15.400 17.885 15.720 ;
      LAYER met4 ;
        RECT 17.565 15.400 17.885 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 14.960 17.885 15.280 ;
      LAYER met4 ;
        RECT 17.565 14.960 17.885 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 18.040 17.480 18.360 ;
      LAYER met4 ;
        RECT 17.160 18.040 17.480 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 17.600 17.480 17.920 ;
      LAYER met4 ;
        RECT 17.160 17.600 17.480 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 17.160 17.480 17.480 ;
      LAYER met4 ;
        RECT 17.160 17.160 17.480 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 16.720 17.480 17.040 ;
      LAYER met4 ;
        RECT 17.160 16.720 17.480 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 16.280 17.480 16.600 ;
      LAYER met4 ;
        RECT 17.160 16.280 17.480 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 15.840 17.480 16.160 ;
      LAYER met4 ;
        RECT 17.160 15.840 17.480 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 15.400 17.480 15.720 ;
      LAYER met4 ;
        RECT 17.160 15.400 17.480 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 14.960 17.480 15.280 ;
      LAYER met4 ;
        RECT 17.160 14.960 17.480 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 18.040 17.075 18.360 ;
      LAYER met4 ;
        RECT 16.755 18.040 17.075 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 17.600 17.075 17.920 ;
      LAYER met4 ;
        RECT 16.755 17.600 17.075 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 17.160 17.075 17.480 ;
      LAYER met4 ;
        RECT 16.755 17.160 17.075 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 16.720 17.075 17.040 ;
      LAYER met4 ;
        RECT 16.755 16.720 17.075 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 16.280 17.075 16.600 ;
      LAYER met4 ;
        RECT 16.755 16.280 17.075 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 15.840 17.075 16.160 ;
      LAYER met4 ;
        RECT 16.755 15.840 17.075 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 15.400 17.075 15.720 ;
      LAYER met4 ;
        RECT 16.755 15.400 17.075 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 14.960 17.075 15.280 ;
      LAYER met4 ;
        RECT 16.755 14.960 17.075 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 18.040 16.670 18.360 ;
      LAYER met4 ;
        RECT 16.350 18.040 16.670 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 17.600 16.670 17.920 ;
      LAYER met4 ;
        RECT 16.350 17.600 16.670 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 17.160 16.670 17.480 ;
      LAYER met4 ;
        RECT 16.350 17.160 16.670 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 16.720 16.670 17.040 ;
      LAYER met4 ;
        RECT 16.350 16.720 16.670 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 16.280 16.670 16.600 ;
      LAYER met4 ;
        RECT 16.350 16.280 16.670 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 15.840 16.670 16.160 ;
      LAYER met4 ;
        RECT 16.350 15.840 16.670 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 15.400 16.670 15.720 ;
      LAYER met4 ;
        RECT 16.350 15.400 16.670 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 14.960 16.670 15.280 ;
      LAYER met4 ;
        RECT 16.350 14.960 16.670 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 18.040 16.265 18.360 ;
      LAYER met4 ;
        RECT 15.945 18.040 16.265 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 17.600 16.265 17.920 ;
      LAYER met4 ;
        RECT 15.945 17.600 16.265 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 17.160 16.265 17.480 ;
      LAYER met4 ;
        RECT 15.945 17.160 16.265 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 16.720 16.265 17.040 ;
      LAYER met4 ;
        RECT 15.945 16.720 16.265 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 16.280 16.265 16.600 ;
      LAYER met4 ;
        RECT 15.945 16.280 16.265 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 15.840 16.265 16.160 ;
      LAYER met4 ;
        RECT 15.945 15.840 16.265 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 15.400 16.265 15.720 ;
      LAYER met4 ;
        RECT 15.945 15.400 16.265 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 14.960 16.265 15.280 ;
      LAYER met4 ;
        RECT 15.945 14.960 16.265 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 18.040 15.860 18.360 ;
      LAYER met4 ;
        RECT 15.540 18.040 15.860 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 17.600 15.860 17.920 ;
      LAYER met4 ;
        RECT 15.540 17.600 15.860 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 17.160 15.860 17.480 ;
      LAYER met4 ;
        RECT 15.540 17.160 15.860 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 16.720 15.860 17.040 ;
      LAYER met4 ;
        RECT 15.540 16.720 15.860 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 16.280 15.860 16.600 ;
      LAYER met4 ;
        RECT 15.540 16.280 15.860 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 15.840 15.860 16.160 ;
      LAYER met4 ;
        RECT 15.540 15.840 15.860 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 15.400 15.860 15.720 ;
      LAYER met4 ;
        RECT 15.540 15.400 15.860 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 14.960 15.860 15.280 ;
      LAYER met4 ;
        RECT 15.540 14.960 15.860 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 18.040 15.455 18.360 ;
      LAYER met4 ;
        RECT 15.135 18.040 15.455 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 17.600 15.455 17.920 ;
      LAYER met4 ;
        RECT 15.135 17.600 15.455 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 17.160 15.455 17.480 ;
      LAYER met4 ;
        RECT 15.135 17.160 15.455 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 16.720 15.455 17.040 ;
      LAYER met4 ;
        RECT 15.135 16.720 15.455 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 16.280 15.455 16.600 ;
      LAYER met4 ;
        RECT 15.135 16.280 15.455 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 15.840 15.455 16.160 ;
      LAYER met4 ;
        RECT 15.135 15.840 15.455 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 15.400 15.455 15.720 ;
      LAYER met4 ;
        RECT 15.135 15.400 15.455 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 14.960 15.455 15.280 ;
      LAYER met4 ;
        RECT 15.135 14.960 15.455 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 18.040 15.050 18.360 ;
      LAYER met4 ;
        RECT 14.730 18.040 15.050 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 17.600 15.050 17.920 ;
      LAYER met4 ;
        RECT 14.730 17.600 15.050 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 17.160 15.050 17.480 ;
      LAYER met4 ;
        RECT 14.730 17.160 15.050 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 16.720 15.050 17.040 ;
      LAYER met4 ;
        RECT 14.730 16.720 15.050 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 16.280 15.050 16.600 ;
      LAYER met4 ;
        RECT 14.730 16.280 15.050 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 15.840 15.050 16.160 ;
      LAYER met4 ;
        RECT 14.730 15.840 15.050 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 15.400 15.050 15.720 ;
      LAYER met4 ;
        RECT 14.730 15.400 15.050 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 14.960 15.050 15.280 ;
      LAYER met4 ;
        RECT 14.730 14.960 15.050 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 18.040 14.645 18.360 ;
      LAYER met4 ;
        RECT 14.325 18.040 14.645 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 17.600 14.645 17.920 ;
      LAYER met4 ;
        RECT 14.325 17.600 14.645 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 17.160 14.645 17.480 ;
      LAYER met4 ;
        RECT 14.325 17.160 14.645 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 16.720 14.645 17.040 ;
      LAYER met4 ;
        RECT 14.325 16.720 14.645 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 16.280 14.645 16.600 ;
      LAYER met4 ;
        RECT 14.325 16.280 14.645 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 15.840 14.645 16.160 ;
      LAYER met4 ;
        RECT 14.325 15.840 14.645 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 15.400 14.645 15.720 ;
      LAYER met4 ;
        RECT 14.325 15.400 14.645 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 14.960 14.645 15.280 ;
      LAYER met4 ;
        RECT 14.325 14.960 14.645 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 18.040 14.240 18.360 ;
      LAYER met4 ;
        RECT 13.920 18.040 14.240 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 17.600 14.240 17.920 ;
      LAYER met4 ;
        RECT 13.920 17.600 14.240 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 17.160 14.240 17.480 ;
      LAYER met4 ;
        RECT 13.920 17.160 14.240 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 16.720 14.240 17.040 ;
      LAYER met4 ;
        RECT 13.920 16.720 14.240 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 16.280 14.240 16.600 ;
      LAYER met4 ;
        RECT 13.920 16.280 14.240 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 15.840 14.240 16.160 ;
      LAYER met4 ;
        RECT 13.920 15.840 14.240 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 15.400 14.240 15.720 ;
      LAYER met4 ;
        RECT 13.920 15.400 14.240 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 14.960 14.240 15.280 ;
      LAYER met4 ;
        RECT 13.920 14.960 14.240 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 18.040 13.835 18.360 ;
      LAYER met4 ;
        RECT 13.515 18.040 13.835 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 17.600 13.835 17.920 ;
      LAYER met4 ;
        RECT 13.515 17.600 13.835 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 17.160 13.835 17.480 ;
      LAYER met4 ;
        RECT 13.515 17.160 13.835 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 16.720 13.835 17.040 ;
      LAYER met4 ;
        RECT 13.515 16.720 13.835 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 16.280 13.835 16.600 ;
      LAYER met4 ;
        RECT 13.515 16.280 13.835 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 15.840 13.835 16.160 ;
      LAYER met4 ;
        RECT 13.515 15.840 13.835 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 15.400 13.835 15.720 ;
      LAYER met4 ;
        RECT 13.515 15.400 13.835 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 14.960 13.835 15.280 ;
      LAYER met4 ;
        RECT 13.515 14.960 13.835 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 18.040 13.430 18.360 ;
      LAYER met4 ;
        RECT 13.110 18.040 13.430 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 17.600 13.430 17.920 ;
      LAYER met4 ;
        RECT 13.110 17.600 13.430 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 17.160 13.430 17.480 ;
      LAYER met4 ;
        RECT 13.110 17.160 13.430 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 16.720 13.430 17.040 ;
      LAYER met4 ;
        RECT 13.110 16.720 13.430 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 16.280 13.430 16.600 ;
      LAYER met4 ;
        RECT 13.110 16.280 13.430 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 15.840 13.430 16.160 ;
      LAYER met4 ;
        RECT 13.110 15.840 13.430 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 15.400 13.430 15.720 ;
      LAYER met4 ;
        RECT 13.110 15.400 13.430 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 14.960 13.430 15.280 ;
      LAYER met4 ;
        RECT 13.110 14.960 13.430 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 18.040 13.025 18.360 ;
      LAYER met4 ;
        RECT 12.705 18.040 13.025 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 17.600 13.025 17.920 ;
      LAYER met4 ;
        RECT 12.705 17.600 13.025 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 17.160 13.025 17.480 ;
      LAYER met4 ;
        RECT 12.705 17.160 13.025 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 16.720 13.025 17.040 ;
      LAYER met4 ;
        RECT 12.705 16.720 13.025 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 16.280 13.025 16.600 ;
      LAYER met4 ;
        RECT 12.705 16.280 13.025 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 15.840 13.025 16.160 ;
      LAYER met4 ;
        RECT 12.705 15.840 13.025 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 15.400 13.025 15.720 ;
      LAYER met4 ;
        RECT 12.705 15.400 13.025 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 14.960 13.025 15.280 ;
      LAYER met4 ;
        RECT 12.705 14.960 13.025 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 18.040 12.620 18.360 ;
      LAYER met4 ;
        RECT 12.300 18.040 12.620 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 17.600 12.620 17.920 ;
      LAYER met4 ;
        RECT 12.300 17.600 12.620 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 17.160 12.620 17.480 ;
      LAYER met4 ;
        RECT 12.300 17.160 12.620 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 16.720 12.620 17.040 ;
      LAYER met4 ;
        RECT 12.300 16.720 12.620 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 16.280 12.620 16.600 ;
      LAYER met4 ;
        RECT 12.300 16.280 12.620 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 15.840 12.620 16.160 ;
      LAYER met4 ;
        RECT 12.300 15.840 12.620 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 15.400 12.620 15.720 ;
      LAYER met4 ;
        RECT 12.300 15.400 12.620 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 14.960 12.620 15.280 ;
      LAYER met4 ;
        RECT 12.300 14.960 12.620 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 18.040 12.215 18.360 ;
      LAYER met4 ;
        RECT 11.895 18.040 12.215 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 17.600 12.215 17.920 ;
      LAYER met4 ;
        RECT 11.895 17.600 12.215 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 17.160 12.215 17.480 ;
      LAYER met4 ;
        RECT 11.895 17.160 12.215 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 16.720 12.215 17.040 ;
      LAYER met4 ;
        RECT 11.895 16.720 12.215 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 16.280 12.215 16.600 ;
      LAYER met4 ;
        RECT 11.895 16.280 12.215 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 15.840 12.215 16.160 ;
      LAYER met4 ;
        RECT 11.895 15.840 12.215 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 15.400 12.215 15.720 ;
      LAYER met4 ;
        RECT 11.895 15.400 12.215 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 14.960 12.215 15.280 ;
      LAYER met4 ;
        RECT 11.895 14.960 12.215 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 18.040 11.810 18.360 ;
      LAYER met4 ;
        RECT 11.490 18.040 11.810 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 17.600 11.810 17.920 ;
      LAYER met4 ;
        RECT 11.490 17.600 11.810 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 17.160 11.810 17.480 ;
      LAYER met4 ;
        RECT 11.490 17.160 11.810 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 16.720 11.810 17.040 ;
      LAYER met4 ;
        RECT 11.490 16.720 11.810 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 16.280 11.810 16.600 ;
      LAYER met4 ;
        RECT 11.490 16.280 11.810 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 15.840 11.810 16.160 ;
      LAYER met4 ;
        RECT 11.490 15.840 11.810 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 15.400 11.810 15.720 ;
      LAYER met4 ;
        RECT 11.490 15.400 11.810 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 14.960 11.810 15.280 ;
      LAYER met4 ;
        RECT 11.490 14.960 11.810 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 18.040 11.405 18.360 ;
      LAYER met4 ;
        RECT 11.085 18.040 11.405 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 17.600 11.405 17.920 ;
      LAYER met4 ;
        RECT 11.085 17.600 11.405 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 17.160 11.405 17.480 ;
      LAYER met4 ;
        RECT 11.085 17.160 11.405 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 16.720 11.405 17.040 ;
      LAYER met4 ;
        RECT 11.085 16.720 11.405 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 16.280 11.405 16.600 ;
      LAYER met4 ;
        RECT 11.085 16.280 11.405 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 15.840 11.405 16.160 ;
      LAYER met4 ;
        RECT 11.085 15.840 11.405 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 15.400 11.405 15.720 ;
      LAYER met4 ;
        RECT 11.085 15.400 11.405 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 14.960 11.405 15.280 ;
      LAYER met4 ;
        RECT 11.085 14.960 11.405 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 18.040 11.000 18.360 ;
      LAYER met4 ;
        RECT 10.680 18.040 11.000 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 17.600 11.000 17.920 ;
      LAYER met4 ;
        RECT 10.680 17.600 11.000 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 17.160 11.000 17.480 ;
      LAYER met4 ;
        RECT 10.680 17.160 11.000 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 16.720 11.000 17.040 ;
      LAYER met4 ;
        RECT 10.680 16.720 11.000 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 16.280 11.000 16.600 ;
      LAYER met4 ;
        RECT 10.680 16.280 11.000 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 15.840 11.000 16.160 ;
      LAYER met4 ;
        RECT 10.680 15.840 11.000 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 15.400 11.000 15.720 ;
      LAYER met4 ;
        RECT 10.680 15.400 11.000 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 14.960 11.000 15.280 ;
      LAYER met4 ;
        RECT 10.680 14.960 11.000 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 18.040 10.595 18.360 ;
      LAYER met4 ;
        RECT 10.275 18.040 10.595 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 17.600 10.595 17.920 ;
      LAYER met4 ;
        RECT 10.275 17.600 10.595 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 17.160 10.595 17.480 ;
      LAYER met4 ;
        RECT 10.275 17.160 10.595 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 16.720 10.595 17.040 ;
      LAYER met4 ;
        RECT 10.275 16.720 10.595 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 16.280 10.595 16.600 ;
      LAYER met4 ;
        RECT 10.275 16.280 10.595 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 15.840 10.595 16.160 ;
      LAYER met4 ;
        RECT 10.275 15.840 10.595 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 15.400 10.595 15.720 ;
      LAYER met4 ;
        RECT 10.275 15.400 10.595 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 14.960 10.595 15.280 ;
      LAYER met4 ;
        RECT 10.275 14.960 10.595 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 18.040 10.190 18.360 ;
      LAYER met4 ;
        RECT 9.870 18.040 10.190 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 17.600 10.190 17.920 ;
      LAYER met4 ;
        RECT 9.870 17.600 10.190 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 17.160 10.190 17.480 ;
      LAYER met4 ;
        RECT 9.870 17.160 10.190 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 16.720 10.190 17.040 ;
      LAYER met4 ;
        RECT 9.870 16.720 10.190 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 16.280 10.190 16.600 ;
      LAYER met4 ;
        RECT 9.870 16.280 10.190 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 15.840 10.190 16.160 ;
      LAYER met4 ;
        RECT 9.870 15.840 10.190 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 15.400 10.190 15.720 ;
      LAYER met4 ;
        RECT 9.870 15.400 10.190 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 14.960 10.190 15.280 ;
      LAYER met4 ;
        RECT 9.870 14.960 10.190 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 18.040 9.785 18.360 ;
      LAYER met4 ;
        RECT 9.465 18.040 9.785 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 17.600 9.785 17.920 ;
      LAYER met4 ;
        RECT 9.465 17.600 9.785 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 17.160 9.785 17.480 ;
      LAYER met4 ;
        RECT 9.465 17.160 9.785 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 16.720 9.785 17.040 ;
      LAYER met4 ;
        RECT 9.465 16.720 9.785 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 16.280 9.785 16.600 ;
      LAYER met4 ;
        RECT 9.465 16.280 9.785 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 15.840 9.785 16.160 ;
      LAYER met4 ;
        RECT 9.465 15.840 9.785 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 15.400 9.785 15.720 ;
      LAYER met4 ;
        RECT 9.465 15.400 9.785 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 14.960 9.785 15.280 ;
      LAYER met4 ;
        RECT 9.465 14.960 9.785 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 18.040 9.380 18.360 ;
      LAYER met4 ;
        RECT 9.060 18.040 9.380 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 17.600 9.380 17.920 ;
      LAYER met4 ;
        RECT 9.060 17.600 9.380 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 17.160 9.380 17.480 ;
      LAYER met4 ;
        RECT 9.060 17.160 9.380 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 16.720 9.380 17.040 ;
      LAYER met4 ;
        RECT 9.060 16.720 9.380 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 16.280 9.380 16.600 ;
      LAYER met4 ;
        RECT 9.060 16.280 9.380 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 15.840 9.380 16.160 ;
      LAYER met4 ;
        RECT 9.060 15.840 9.380 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 15.400 9.380 15.720 ;
      LAYER met4 ;
        RECT 9.060 15.400 9.380 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 14.960 9.380 15.280 ;
      LAYER met4 ;
        RECT 9.060 14.960 9.380 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 18.040 8.975 18.360 ;
      LAYER met4 ;
        RECT 8.655 18.040 8.975 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 17.600 8.975 17.920 ;
      LAYER met4 ;
        RECT 8.655 17.600 8.975 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 17.160 8.975 17.480 ;
      LAYER met4 ;
        RECT 8.655 17.160 8.975 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 16.720 8.975 17.040 ;
      LAYER met4 ;
        RECT 8.655 16.720 8.975 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 16.280 8.975 16.600 ;
      LAYER met4 ;
        RECT 8.655 16.280 8.975 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 15.840 8.975 16.160 ;
      LAYER met4 ;
        RECT 8.655 15.840 8.975 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 15.400 8.975 15.720 ;
      LAYER met4 ;
        RECT 8.655 15.400 8.975 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 14.960 8.975 15.280 ;
      LAYER met4 ;
        RECT 8.655 14.960 8.975 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 18.040 8.570 18.360 ;
      LAYER met4 ;
        RECT 8.250 18.040 8.570 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 17.600 8.570 17.920 ;
      LAYER met4 ;
        RECT 8.250 17.600 8.570 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 17.160 8.570 17.480 ;
      LAYER met4 ;
        RECT 8.250 17.160 8.570 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 16.720 8.570 17.040 ;
      LAYER met4 ;
        RECT 8.250 16.720 8.570 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 16.280 8.570 16.600 ;
      LAYER met4 ;
        RECT 8.250 16.280 8.570 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 15.840 8.570 16.160 ;
      LAYER met4 ;
        RECT 8.250 15.840 8.570 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 15.400 8.570 15.720 ;
      LAYER met4 ;
        RECT 8.250 15.400 8.570 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 14.960 8.570 15.280 ;
      LAYER met4 ;
        RECT 8.250 14.960 8.570 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 18.040 8.165 18.360 ;
      LAYER met4 ;
        RECT 7.845 18.040 8.165 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 17.600 8.165 17.920 ;
      LAYER met4 ;
        RECT 7.845 17.600 8.165 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 17.160 8.165 17.480 ;
      LAYER met4 ;
        RECT 7.845 17.160 8.165 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 16.720 8.165 17.040 ;
      LAYER met4 ;
        RECT 7.845 16.720 8.165 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 16.280 8.165 16.600 ;
      LAYER met4 ;
        RECT 7.845 16.280 8.165 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 15.840 8.165 16.160 ;
      LAYER met4 ;
        RECT 7.845 15.840 8.165 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 15.400 8.165 15.720 ;
      LAYER met4 ;
        RECT 7.845 15.400 8.165 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 14.960 8.165 15.280 ;
      LAYER met4 ;
        RECT 7.845 14.960 8.165 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 18.040 7.760 18.360 ;
      LAYER met4 ;
        RECT 7.440 18.040 7.760 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 17.600 7.760 17.920 ;
      LAYER met4 ;
        RECT 7.440 17.600 7.760 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 17.160 7.760 17.480 ;
      LAYER met4 ;
        RECT 7.440 17.160 7.760 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 16.720 7.760 17.040 ;
      LAYER met4 ;
        RECT 7.440 16.720 7.760 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 16.280 7.760 16.600 ;
      LAYER met4 ;
        RECT 7.440 16.280 7.760 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 15.840 7.760 16.160 ;
      LAYER met4 ;
        RECT 7.440 15.840 7.760 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 15.400 7.760 15.720 ;
      LAYER met4 ;
        RECT 7.440 15.400 7.760 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 14.960 7.760 15.280 ;
      LAYER met4 ;
        RECT 7.440 14.960 7.760 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 18.040 7.355 18.360 ;
      LAYER met4 ;
        RECT 7.035 18.040 7.355 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 17.600 7.355 17.920 ;
      LAYER met4 ;
        RECT 7.035 17.600 7.355 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 17.160 7.355 17.480 ;
      LAYER met4 ;
        RECT 7.035 17.160 7.355 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 16.720 7.355 17.040 ;
      LAYER met4 ;
        RECT 7.035 16.720 7.355 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 16.280 7.355 16.600 ;
      LAYER met4 ;
        RECT 7.035 16.280 7.355 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 15.840 7.355 16.160 ;
      LAYER met4 ;
        RECT 7.035 15.840 7.355 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 15.400 7.355 15.720 ;
      LAYER met4 ;
        RECT 7.035 15.400 7.355 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 14.960 7.355 15.280 ;
      LAYER met4 ;
        RECT 7.035 14.960 7.355 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 18.040 6.950 18.360 ;
      LAYER met4 ;
        RECT 6.630 18.040 6.950 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 17.600 6.950 17.920 ;
      LAYER met4 ;
        RECT 6.630 17.600 6.950 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 17.160 6.950 17.480 ;
      LAYER met4 ;
        RECT 6.630 17.160 6.950 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 16.720 6.950 17.040 ;
      LAYER met4 ;
        RECT 6.630 16.720 6.950 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 16.280 6.950 16.600 ;
      LAYER met4 ;
        RECT 6.630 16.280 6.950 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 15.840 6.950 16.160 ;
      LAYER met4 ;
        RECT 6.630 15.840 6.950 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 15.400 6.950 15.720 ;
      LAYER met4 ;
        RECT 6.630 15.400 6.950 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 14.960 6.950 15.280 ;
      LAYER met4 ;
        RECT 6.630 14.960 6.950 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 18.040 6.545 18.360 ;
      LAYER met4 ;
        RECT 6.225 18.040 6.545 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 17.600 6.545 17.920 ;
      LAYER met4 ;
        RECT 6.225 17.600 6.545 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 17.160 6.545 17.480 ;
      LAYER met4 ;
        RECT 6.225 17.160 6.545 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 16.720 6.545 17.040 ;
      LAYER met4 ;
        RECT 6.225 16.720 6.545 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 16.280 6.545 16.600 ;
      LAYER met4 ;
        RECT 6.225 16.280 6.545 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 15.840 6.545 16.160 ;
      LAYER met4 ;
        RECT 6.225 15.840 6.545 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 15.400 6.545 15.720 ;
      LAYER met4 ;
        RECT 6.225 15.400 6.545 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 14.960 6.545 15.280 ;
      LAYER met4 ;
        RECT 6.225 14.960 6.545 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 18.040 6.140 18.360 ;
      LAYER met4 ;
        RECT 5.820 18.040 6.140 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 17.600 6.140 17.920 ;
      LAYER met4 ;
        RECT 5.820 17.600 6.140 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 17.160 6.140 17.480 ;
      LAYER met4 ;
        RECT 5.820 17.160 6.140 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 16.720 6.140 17.040 ;
      LAYER met4 ;
        RECT 5.820 16.720 6.140 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 16.280 6.140 16.600 ;
      LAYER met4 ;
        RECT 5.820 16.280 6.140 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 15.840 6.140 16.160 ;
      LAYER met4 ;
        RECT 5.820 15.840 6.140 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 15.400 6.140 15.720 ;
      LAYER met4 ;
        RECT 5.820 15.400 6.140 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 14.960 6.140 15.280 ;
      LAYER met4 ;
        RECT 5.820 14.960 6.140 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 18.040 5.735 18.360 ;
      LAYER met4 ;
        RECT 5.415 18.040 5.735 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 17.600 5.735 17.920 ;
      LAYER met4 ;
        RECT 5.415 17.600 5.735 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 17.160 5.735 17.480 ;
      LAYER met4 ;
        RECT 5.415 17.160 5.735 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 16.720 5.735 17.040 ;
      LAYER met4 ;
        RECT 5.415 16.720 5.735 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 16.280 5.735 16.600 ;
      LAYER met4 ;
        RECT 5.415 16.280 5.735 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 15.840 5.735 16.160 ;
      LAYER met4 ;
        RECT 5.415 15.840 5.735 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 15.400 5.735 15.720 ;
      LAYER met4 ;
        RECT 5.415 15.400 5.735 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 14.960 5.735 15.280 ;
      LAYER met4 ;
        RECT 5.415 14.960 5.735 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 18.040 5.330 18.360 ;
      LAYER met4 ;
        RECT 5.010 18.040 5.330 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 17.600 5.330 17.920 ;
      LAYER met4 ;
        RECT 5.010 17.600 5.330 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 17.160 5.330 17.480 ;
      LAYER met4 ;
        RECT 5.010 17.160 5.330 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 16.720 5.330 17.040 ;
      LAYER met4 ;
        RECT 5.010 16.720 5.330 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 16.280 5.330 16.600 ;
      LAYER met4 ;
        RECT 5.010 16.280 5.330 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 15.840 5.330 16.160 ;
      LAYER met4 ;
        RECT 5.010 15.840 5.330 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 15.400 5.330 15.720 ;
      LAYER met4 ;
        RECT 5.010 15.400 5.330 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 14.960 5.330 15.280 ;
      LAYER met4 ;
        RECT 5.010 14.960 5.330 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 18.040 4.925 18.360 ;
      LAYER met4 ;
        RECT 4.605 18.040 4.925 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 17.600 4.925 17.920 ;
      LAYER met4 ;
        RECT 4.605 17.600 4.925 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 17.160 4.925 17.480 ;
      LAYER met4 ;
        RECT 4.605 17.160 4.925 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 16.720 4.925 17.040 ;
      LAYER met4 ;
        RECT 4.605 16.720 4.925 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 16.280 4.925 16.600 ;
      LAYER met4 ;
        RECT 4.605 16.280 4.925 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 15.840 4.925 16.160 ;
      LAYER met4 ;
        RECT 4.605 15.840 4.925 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 15.400 4.925 15.720 ;
      LAYER met4 ;
        RECT 4.605 15.400 4.925 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 14.960 4.925 15.280 ;
      LAYER met4 ;
        RECT 4.605 14.960 4.925 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 18.040 4.520 18.360 ;
      LAYER met4 ;
        RECT 4.200 18.040 4.520 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 17.600 4.520 17.920 ;
      LAYER met4 ;
        RECT 4.200 17.600 4.520 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 17.160 4.520 17.480 ;
      LAYER met4 ;
        RECT 4.200 17.160 4.520 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 16.720 4.520 17.040 ;
      LAYER met4 ;
        RECT 4.200 16.720 4.520 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 16.280 4.520 16.600 ;
      LAYER met4 ;
        RECT 4.200 16.280 4.520 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 15.840 4.520 16.160 ;
      LAYER met4 ;
        RECT 4.200 15.840 4.520 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 15.400 4.520 15.720 ;
      LAYER met4 ;
        RECT 4.200 15.400 4.520 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 14.960 4.520 15.280 ;
      LAYER met4 ;
        RECT 4.200 14.960 4.520 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 18.040 4.115 18.360 ;
      LAYER met4 ;
        RECT 3.795 18.040 4.115 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 17.600 4.115 17.920 ;
      LAYER met4 ;
        RECT 3.795 17.600 4.115 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 17.160 4.115 17.480 ;
      LAYER met4 ;
        RECT 3.795 17.160 4.115 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 16.720 4.115 17.040 ;
      LAYER met4 ;
        RECT 3.795 16.720 4.115 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 16.280 4.115 16.600 ;
      LAYER met4 ;
        RECT 3.795 16.280 4.115 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 15.840 4.115 16.160 ;
      LAYER met4 ;
        RECT 3.795 15.840 4.115 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 15.400 4.115 15.720 ;
      LAYER met4 ;
        RECT 3.795 15.400 4.115 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 14.960 4.115 15.280 ;
      LAYER met4 ;
        RECT 3.795 14.960 4.115 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 18.040 3.710 18.360 ;
      LAYER met4 ;
        RECT 3.390 18.040 3.710 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 17.600 3.710 17.920 ;
      LAYER met4 ;
        RECT 3.390 17.600 3.710 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 17.160 3.710 17.480 ;
      LAYER met4 ;
        RECT 3.390 17.160 3.710 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 16.720 3.710 17.040 ;
      LAYER met4 ;
        RECT 3.390 16.720 3.710 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 16.280 3.710 16.600 ;
      LAYER met4 ;
        RECT 3.390 16.280 3.710 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 15.840 3.710 16.160 ;
      LAYER met4 ;
        RECT 3.390 15.840 3.710 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 15.400 3.710 15.720 ;
      LAYER met4 ;
        RECT 3.390 15.400 3.710 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 14.960 3.710 15.280 ;
      LAYER met4 ;
        RECT 3.390 14.960 3.710 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 18.040 3.305 18.360 ;
      LAYER met4 ;
        RECT 2.985 18.040 3.305 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 17.600 3.305 17.920 ;
      LAYER met4 ;
        RECT 2.985 17.600 3.305 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 17.160 3.305 17.480 ;
      LAYER met4 ;
        RECT 2.985 17.160 3.305 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 16.720 3.305 17.040 ;
      LAYER met4 ;
        RECT 2.985 16.720 3.305 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 16.280 3.305 16.600 ;
      LAYER met4 ;
        RECT 2.985 16.280 3.305 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 15.840 3.305 16.160 ;
      LAYER met4 ;
        RECT 2.985 15.840 3.305 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 15.400 3.305 15.720 ;
      LAYER met4 ;
        RECT 2.985 15.400 3.305 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 14.960 3.305 15.280 ;
      LAYER met4 ;
        RECT 2.985 14.960 3.305 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 18.040 2.895 18.360 ;
      LAYER met4 ;
        RECT 2.575 18.040 2.895 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 17.600 2.895 17.920 ;
      LAYER met4 ;
        RECT 2.575 17.600 2.895 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 17.160 2.895 17.480 ;
      LAYER met4 ;
        RECT 2.575 17.160 2.895 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 16.720 2.895 17.040 ;
      LAYER met4 ;
        RECT 2.575 16.720 2.895 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 16.280 2.895 16.600 ;
      LAYER met4 ;
        RECT 2.575 16.280 2.895 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 15.840 2.895 16.160 ;
      LAYER met4 ;
        RECT 2.575 15.840 2.895 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 15.400 2.895 15.720 ;
      LAYER met4 ;
        RECT 2.575 15.400 2.895 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 14.960 2.895 15.280 ;
      LAYER met4 ;
        RECT 2.575 14.960 2.895 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 18.040 2.485 18.360 ;
      LAYER met4 ;
        RECT 2.165 18.040 2.485 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 17.600 2.485 17.920 ;
      LAYER met4 ;
        RECT 2.165 17.600 2.485 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 17.160 2.485 17.480 ;
      LAYER met4 ;
        RECT 2.165 17.160 2.485 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 16.720 2.485 17.040 ;
      LAYER met4 ;
        RECT 2.165 16.720 2.485 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 16.280 2.485 16.600 ;
      LAYER met4 ;
        RECT 2.165 16.280 2.485 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 15.840 2.485 16.160 ;
      LAYER met4 ;
        RECT 2.165 15.840 2.485 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 15.400 2.485 15.720 ;
      LAYER met4 ;
        RECT 2.165 15.400 2.485 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 14.960 2.485 15.280 ;
      LAYER met4 ;
        RECT 2.165 14.960 2.485 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 18.040 2.075 18.360 ;
      LAYER met4 ;
        RECT 1.755 18.040 2.075 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 17.600 2.075 17.920 ;
      LAYER met4 ;
        RECT 1.755 17.600 2.075 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 17.160 2.075 17.480 ;
      LAYER met4 ;
        RECT 1.755 17.160 2.075 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 16.720 2.075 17.040 ;
      LAYER met4 ;
        RECT 1.755 16.720 2.075 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 16.280 2.075 16.600 ;
      LAYER met4 ;
        RECT 1.755 16.280 2.075 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 15.840 2.075 16.160 ;
      LAYER met4 ;
        RECT 1.755 15.840 2.075 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 15.400 2.075 15.720 ;
      LAYER met4 ;
        RECT 1.755 15.400 2.075 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 14.960 2.075 15.280 ;
      LAYER met4 ;
        RECT 1.755 14.960 2.075 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 18.040 1.665 18.360 ;
      LAYER met4 ;
        RECT 1.345 18.040 1.665 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 17.600 1.665 17.920 ;
      LAYER met4 ;
        RECT 1.345 17.600 1.665 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 17.160 1.665 17.480 ;
      LAYER met4 ;
        RECT 1.345 17.160 1.665 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 16.720 1.665 17.040 ;
      LAYER met4 ;
        RECT 1.345 16.720 1.665 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 16.280 1.665 16.600 ;
      LAYER met4 ;
        RECT 1.345 16.280 1.665 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 15.840 1.665 16.160 ;
      LAYER met4 ;
        RECT 1.345 15.840 1.665 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 15.400 1.665 15.720 ;
      LAYER met4 ;
        RECT 1.345 15.400 1.665 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 14.960 1.665 15.280 ;
      LAYER met4 ;
        RECT 1.345 14.960 1.665 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 18.040 1.255 18.360 ;
      LAYER met4 ;
        RECT 0.965 18.040 1.255 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 17.600 1.255 17.920 ;
      LAYER met4 ;
        RECT 0.965 17.600 1.255 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 17.160 1.255 17.480 ;
      LAYER met4 ;
        RECT 0.965 17.160 1.255 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 16.720 1.255 17.040 ;
      LAYER met4 ;
        RECT 0.965 16.720 1.255 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 16.280 1.255 16.600 ;
      LAYER met4 ;
        RECT 0.965 16.280 1.255 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 15.840 1.255 16.160 ;
      LAYER met4 ;
        RECT 0.965 15.840 1.255 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 15.400 1.255 15.720 ;
      LAYER met4 ;
        RECT 0.965 15.400 1.255 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 14.960 1.255 15.280 ;
      LAYER met4 ;
        RECT 0.965 14.960 1.255 15.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 18.040 0.845 18.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 17.600 0.845 17.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 17.160 0.845 17.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 16.720 0.845 17.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 16.280 0.845 16.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 15.840 0.845 16.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 15.400 0.845 15.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 14.960 0.845 15.280 ;
    END
  END VDDA
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
  END VSSIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
  END VCCHIB
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
  END VSWITCH
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.495 14.940 24.395 18.380 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 96.585 75.000 174.185 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__overlay_vdda_hvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vdda_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vdda_lvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
  END VSWITCH
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 12.940 74.655 16.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 16.100 74.565 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 15.660 74.565 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 15.220 74.565 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 14.780 74.565 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 14.340 74.565 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 13.900 74.565 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 13.460 74.565 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 13.020 74.565 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 16.100 74.160 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 15.660 74.160 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 15.220 74.160 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 14.780 74.160 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 14.340 74.160 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 13.900 74.160 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 13.460 74.160 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 13.020 74.160 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 16.100 73.755 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 15.660 73.755 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 15.220 73.755 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 14.780 73.755 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 14.340 73.755 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 13.900 73.755 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 13.460 73.755 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 13.020 73.755 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 16.100 73.350 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 15.660 73.350 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 15.220 73.350 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 14.780 73.350 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 14.340 73.350 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 13.900 73.350 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 13.460 73.350 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 13.020 73.350 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 16.100 72.945 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 15.660 72.945 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 15.220 72.945 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 14.780 72.945 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 14.340 72.945 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 13.900 72.945 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 13.460 72.945 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 13.020 72.945 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 16.100 72.540 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 15.660 72.540 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 15.220 72.540 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 14.780 72.540 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 14.340 72.540 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 13.900 72.540 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 13.460 72.540 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 13.020 72.540 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 16.100 72.135 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 15.660 72.135 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 15.220 72.135 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 14.780 72.135 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 14.340 72.135 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 13.900 72.135 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 13.460 72.135 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 13.020 72.135 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 16.100 71.730 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 15.660 71.730 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 15.220 71.730 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 14.780 71.730 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 14.340 71.730 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 13.900 71.730 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 13.460 71.730 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 13.020 71.730 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 16.100 71.325 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 15.660 71.325 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 15.220 71.325 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 14.780 71.325 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 14.340 71.325 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 13.900 71.325 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 13.460 71.325 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 13.020 71.325 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 16.100 70.920 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 15.660 70.920 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 15.220 70.920 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 14.780 70.920 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 14.340 70.920 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 13.900 70.920 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 13.460 70.920 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 13.020 70.920 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 16.100 70.515 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 15.660 70.515 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 15.220 70.515 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 14.780 70.515 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 14.340 70.515 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 13.900 70.515 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 13.460 70.515 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 13.020 70.515 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 16.100 70.110 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 15.660 70.110 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 15.220 70.110 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 14.780 70.110 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 14.340 70.110 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 13.900 70.110 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 13.460 70.110 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 13.020 70.110 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 16.100 69.705 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 15.660 69.705 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 15.220 69.705 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 14.780 69.705 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 14.340 69.705 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 13.900 69.705 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 13.460 69.705 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 13.020 69.705 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 16.100 69.300 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 15.660 69.300 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 15.220 69.300 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 14.780 69.300 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 14.340 69.300 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 13.900 69.300 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 13.460 69.300 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 13.020 69.300 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 16.100 68.895 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 15.660 68.895 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 15.220 68.895 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 14.780 68.895 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 14.340 68.895 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 13.900 68.895 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 13.460 68.895 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 13.020 68.895 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 16.100 68.490 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 15.660 68.490 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 15.220 68.490 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 14.780 68.490 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 14.340 68.490 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 13.900 68.490 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 13.460 68.490 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 13.020 68.490 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 16.100 68.085 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 15.660 68.085 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 15.220 68.085 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 14.780 68.085 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 14.340 68.085 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 13.900 68.085 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 13.460 68.085 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 13.020 68.085 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 16.100 67.680 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 15.660 67.680 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 15.220 67.680 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 14.780 67.680 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 14.340 67.680 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 13.900 67.680 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 13.460 67.680 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 13.020 67.680 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 16.100 67.275 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 15.660 67.275 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 15.220 67.275 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 14.780 67.275 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 14.340 67.275 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 13.900 67.275 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 13.460 67.275 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 13.020 67.275 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 16.100 66.870 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 15.660 66.870 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 15.220 66.870 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 14.780 66.870 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 14.340 66.870 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 13.900 66.870 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 13.460 66.870 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 13.020 66.870 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 16.100 66.465 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 15.660 66.465 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 15.220 66.465 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 14.780 66.465 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 14.340 66.465 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 13.900 66.465 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 13.460 66.465 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 13.020 66.465 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 16.100 66.060 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 15.660 66.060 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 15.220 66.060 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 14.780 66.060 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 14.340 66.060 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 13.900 66.060 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 13.460 66.060 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 13.020 66.060 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 16.100 65.655 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 15.660 65.655 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 15.220 65.655 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 14.780 65.655 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 14.340 65.655 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 13.900 65.655 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 13.460 65.655 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 13.020 65.655 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 16.100 65.250 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 15.660 65.250 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 15.220 65.250 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 14.780 65.250 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 14.340 65.250 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 13.900 65.250 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 13.460 65.250 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 13.020 65.250 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 16.100 64.845 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 15.660 64.845 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 15.220 64.845 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 14.780 64.845 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 14.340 64.845 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 13.900 64.845 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 13.460 64.845 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 13.020 64.845 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 16.100 64.440 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 15.660 64.440 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 15.220 64.440 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 14.780 64.440 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 14.340 64.440 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 13.900 64.440 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 13.460 64.440 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 13.020 64.440 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 16.100 64.035 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 15.660 64.035 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 15.220 64.035 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 14.780 64.035 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 14.340 64.035 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 13.900 64.035 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 13.460 64.035 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 13.020 64.035 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 16.100 63.630 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 15.660 63.630 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 15.220 63.630 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 14.780 63.630 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 14.340 63.630 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 13.900 63.630 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 13.460 63.630 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 13.020 63.630 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 16.100 63.225 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 15.660 63.225 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 15.220 63.225 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 14.780 63.225 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 14.340 63.225 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 13.900 63.225 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 13.460 63.225 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 13.020 63.225 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 16.100 62.820 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 15.660 62.820 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 15.220 62.820 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 14.780 62.820 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 14.340 62.820 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 13.900 62.820 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 13.460 62.820 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 13.020 62.820 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 16.100 62.415 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 15.660 62.415 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 15.220 62.415 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 14.780 62.415 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 14.340 62.415 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 13.900 62.415 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 13.460 62.415 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 13.020 62.415 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 16.100 62.010 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 15.660 62.010 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 15.220 62.010 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 14.780 62.010 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 14.340 62.010 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 13.900 62.010 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 13.460 62.010 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 13.020 62.010 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 16.100 61.605 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 15.660 61.605 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 15.220 61.605 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 14.780 61.605 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 14.340 61.605 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 13.900 61.605 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 13.460 61.605 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 13.020 61.605 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 16.100 61.200 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 15.660 61.200 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 15.220 61.200 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 14.780 61.200 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 14.340 61.200 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 13.900 61.200 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 13.460 61.200 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 13.020 61.200 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 16.100 60.795 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 15.660 60.795 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 15.220 60.795 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 14.780 60.795 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 14.340 60.795 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 13.900 60.795 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 13.460 60.795 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 13.020 60.795 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 16.100 60.390 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 15.660 60.390 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 15.220 60.390 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 14.780 60.390 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 14.340 60.390 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 13.900 60.390 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 13.460 60.390 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 13.020 60.390 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 16.100 59.985 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 15.660 59.985 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 15.220 59.985 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 14.780 59.985 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 14.340 59.985 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 13.900 59.985 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 13.460 59.985 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 13.020 59.985 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 16.100 59.580 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 15.660 59.580 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 15.220 59.580 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 14.780 59.580 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 14.340 59.580 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 13.900 59.580 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 13.460 59.580 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 13.020 59.580 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 16.100 59.175 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 15.660 59.175 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 15.220 59.175 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 14.780 59.175 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 14.340 59.175 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 13.900 59.175 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 13.460 59.175 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 13.020 59.175 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 16.100 58.770 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 15.660 58.770 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 15.220 58.770 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 14.780 58.770 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 14.340 58.770 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 13.900 58.770 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 13.460 58.770 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 13.020 58.770 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 16.100 58.365 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 15.660 58.365 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 15.220 58.365 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 14.780 58.365 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 14.340 58.365 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 13.900 58.365 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 13.460 58.365 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 13.020 58.365 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 16.100 57.960 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 15.660 57.960 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 15.220 57.960 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 14.780 57.960 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 14.340 57.960 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 13.900 57.960 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 13.460 57.960 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 13.020 57.960 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 16.100 57.555 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 15.660 57.555 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 15.220 57.555 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 14.780 57.555 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 14.340 57.555 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 13.900 57.555 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 13.460 57.555 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 13.020 57.555 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 16.100 57.150 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 15.660 57.150 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 15.220 57.150 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 14.780 57.150 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 14.340 57.150 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 13.900 57.150 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 13.460 57.150 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 13.020 57.150 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 16.100 56.745 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 15.660 56.745 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 15.220 56.745 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 14.780 56.745 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 14.340 56.745 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 13.900 56.745 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 13.460 56.745 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 13.020 56.745 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 16.100 56.340 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 15.660 56.340 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 15.220 56.340 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 14.780 56.340 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 14.340 56.340 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 13.900 56.340 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 13.460 56.340 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 13.020 56.340 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 16.100 55.935 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 15.660 55.935 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 15.220 55.935 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 14.780 55.935 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 14.340 55.935 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 13.900 55.935 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 13.460 55.935 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 13.020 55.935 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 16.100 55.530 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 15.660 55.530 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 15.220 55.530 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 14.780 55.530 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 14.340 55.530 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 13.900 55.530 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 13.460 55.530 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 13.020 55.530 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 16.100 55.125 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 15.660 55.125 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 15.220 55.125 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 14.780 55.125 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 14.340 55.125 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 13.900 55.125 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 13.460 55.125 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 13.020 55.125 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 16.100 54.720 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 15.660 54.720 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 15.220 54.720 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 14.780 54.720 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 14.340 54.720 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 13.900 54.720 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 13.460 54.720 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 13.020 54.720 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 16.100 54.315 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 15.660 54.315 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 15.220 54.315 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 14.780 54.315 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 14.340 54.315 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 13.900 54.315 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 13.460 54.315 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 13.020 54.315 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 16.100 53.910 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 15.660 53.910 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 15.220 53.910 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 14.780 53.910 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 14.340 53.910 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 13.900 53.910 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 13.460 53.910 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 13.020 53.910 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 16.100 53.505 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 15.660 53.505 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 15.220 53.505 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 14.780 53.505 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 14.340 53.505 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 13.900 53.505 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 13.460 53.505 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 13.020 53.505 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 16.100 53.095 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 15.660 53.095 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 15.220 53.095 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 14.780 53.095 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 14.340 53.095 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 13.900 53.095 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 13.460 53.095 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 13.020 53.095 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 16.100 52.685 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 15.660 52.685 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 15.220 52.685 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 14.780 52.685 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 14.340 52.685 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 13.900 52.685 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 13.460 52.685 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 13.020 52.685 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 16.100 52.275 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 15.660 52.275 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 15.220 52.275 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 14.780 52.275 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 14.340 52.275 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 13.900 52.275 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 13.460 52.275 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 13.020 52.275 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 16.100 51.865 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 15.660 51.865 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 15.220 51.865 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 14.780 51.865 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 14.340 51.865 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 13.900 51.865 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 13.460 51.865 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 13.020 51.865 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 16.100 51.455 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 15.660 51.455 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 15.220 51.455 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 14.780 51.455 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 14.340 51.455 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 13.900 51.455 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 13.460 51.455 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 13.020 51.455 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 16.100 51.045 16.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 15.660 51.045 15.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 15.220 51.045 15.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 14.780 51.045 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 14.340 51.045 14.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 13.900 51.045 14.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 13.460 51.045 13.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 13.020 51.045 13.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 16.040 24.470 16.360 ;
      LAYER met4 ;
        RECT 24.150 16.040 24.470 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 15.600 24.470 15.920 ;
      LAYER met4 ;
        RECT 24.150 15.600 24.470 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 15.160 24.470 15.480 ;
      LAYER met4 ;
        RECT 24.150 15.160 24.470 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 14.720 24.470 15.040 ;
      LAYER met4 ;
        RECT 24.150 14.720 24.470 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 14.280 24.470 14.600 ;
      LAYER met4 ;
        RECT 24.150 14.280 24.470 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 13.840 24.470 14.160 ;
      LAYER met4 ;
        RECT 24.150 13.840 24.470 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 13.400 24.470 13.720 ;
      LAYER met4 ;
        RECT 24.150 13.400 24.470 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 12.960 24.470 13.280 ;
      LAYER met4 ;
        RECT 24.150 12.960 24.470 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 16.040 24.065 16.360 ;
      LAYER met4 ;
        RECT 23.745 16.040 24.065 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 15.600 24.065 15.920 ;
      LAYER met4 ;
        RECT 23.745 15.600 24.065 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 15.160 24.065 15.480 ;
      LAYER met4 ;
        RECT 23.745 15.160 24.065 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 14.720 24.065 15.040 ;
      LAYER met4 ;
        RECT 23.745 14.720 24.065 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 14.280 24.065 14.600 ;
      LAYER met4 ;
        RECT 23.745 14.280 24.065 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 13.840 24.065 14.160 ;
      LAYER met4 ;
        RECT 23.745 13.840 24.065 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 13.400 24.065 13.720 ;
      LAYER met4 ;
        RECT 23.745 13.400 24.065 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 12.960 24.065 13.280 ;
      LAYER met4 ;
        RECT 23.745 12.960 24.065 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 16.040 23.660 16.360 ;
      LAYER met4 ;
        RECT 23.340 16.040 23.660 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 15.600 23.660 15.920 ;
      LAYER met4 ;
        RECT 23.340 15.600 23.660 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 15.160 23.660 15.480 ;
      LAYER met4 ;
        RECT 23.340 15.160 23.660 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 14.720 23.660 15.040 ;
      LAYER met4 ;
        RECT 23.340 14.720 23.660 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 14.280 23.660 14.600 ;
      LAYER met4 ;
        RECT 23.340 14.280 23.660 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 13.840 23.660 14.160 ;
      LAYER met4 ;
        RECT 23.340 13.840 23.660 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 13.400 23.660 13.720 ;
      LAYER met4 ;
        RECT 23.340 13.400 23.660 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.340 12.960 23.660 13.280 ;
      LAYER met4 ;
        RECT 23.340 12.960 23.660 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 16.040 23.255 16.360 ;
      LAYER met4 ;
        RECT 22.935 16.040 23.255 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 15.600 23.255 15.920 ;
      LAYER met4 ;
        RECT 22.935 15.600 23.255 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 15.160 23.255 15.480 ;
      LAYER met4 ;
        RECT 22.935 15.160 23.255 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 14.720 23.255 15.040 ;
      LAYER met4 ;
        RECT 22.935 14.720 23.255 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 14.280 23.255 14.600 ;
      LAYER met4 ;
        RECT 22.935 14.280 23.255 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 13.840 23.255 14.160 ;
      LAYER met4 ;
        RECT 22.935 13.840 23.255 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 13.400 23.255 13.720 ;
      LAYER met4 ;
        RECT 22.935 13.400 23.255 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.935 12.960 23.255 13.280 ;
      LAYER met4 ;
        RECT 22.935 12.960 23.255 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 16.040 22.850 16.360 ;
      LAYER met4 ;
        RECT 22.530 16.040 22.850 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 15.600 22.850 15.920 ;
      LAYER met4 ;
        RECT 22.530 15.600 22.850 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 15.160 22.850 15.480 ;
      LAYER met4 ;
        RECT 22.530 15.160 22.850 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 14.720 22.850 15.040 ;
      LAYER met4 ;
        RECT 22.530 14.720 22.850 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 14.280 22.850 14.600 ;
      LAYER met4 ;
        RECT 22.530 14.280 22.850 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 13.840 22.850 14.160 ;
      LAYER met4 ;
        RECT 22.530 13.840 22.850 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 13.400 22.850 13.720 ;
      LAYER met4 ;
        RECT 22.530 13.400 22.850 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.530 12.960 22.850 13.280 ;
      LAYER met4 ;
        RECT 22.530 12.960 22.850 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 16.040 22.445 16.360 ;
      LAYER met4 ;
        RECT 22.125 16.040 22.445 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 15.600 22.445 15.920 ;
      LAYER met4 ;
        RECT 22.125 15.600 22.445 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 15.160 22.445 15.480 ;
      LAYER met4 ;
        RECT 22.125 15.160 22.445 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 14.720 22.445 15.040 ;
      LAYER met4 ;
        RECT 22.125 14.720 22.445 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 14.280 22.445 14.600 ;
      LAYER met4 ;
        RECT 22.125 14.280 22.445 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 13.840 22.445 14.160 ;
      LAYER met4 ;
        RECT 22.125 13.840 22.445 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 13.400 22.445 13.720 ;
      LAYER met4 ;
        RECT 22.125 13.400 22.445 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.125 12.960 22.445 13.280 ;
      LAYER met4 ;
        RECT 22.125 12.960 22.445 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 16.040 22.040 16.360 ;
      LAYER met4 ;
        RECT 21.720 16.040 22.040 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 15.600 22.040 15.920 ;
      LAYER met4 ;
        RECT 21.720 15.600 22.040 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 15.160 22.040 15.480 ;
      LAYER met4 ;
        RECT 21.720 15.160 22.040 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 14.720 22.040 15.040 ;
      LAYER met4 ;
        RECT 21.720 14.720 22.040 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 14.280 22.040 14.600 ;
      LAYER met4 ;
        RECT 21.720 14.280 22.040 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 13.840 22.040 14.160 ;
      LAYER met4 ;
        RECT 21.720 13.840 22.040 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 13.400 22.040 13.720 ;
      LAYER met4 ;
        RECT 21.720 13.400 22.040 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.720 12.960 22.040 13.280 ;
      LAYER met4 ;
        RECT 21.720 12.960 22.040 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 16.040 21.635 16.360 ;
      LAYER met4 ;
        RECT 21.315 16.040 21.635 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 15.600 21.635 15.920 ;
      LAYER met4 ;
        RECT 21.315 15.600 21.635 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 15.160 21.635 15.480 ;
      LAYER met4 ;
        RECT 21.315 15.160 21.635 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 14.720 21.635 15.040 ;
      LAYER met4 ;
        RECT 21.315 14.720 21.635 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 14.280 21.635 14.600 ;
      LAYER met4 ;
        RECT 21.315 14.280 21.635 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 13.840 21.635 14.160 ;
      LAYER met4 ;
        RECT 21.315 13.840 21.635 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 13.400 21.635 13.720 ;
      LAYER met4 ;
        RECT 21.315 13.400 21.635 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.315 12.960 21.635 13.280 ;
      LAYER met4 ;
        RECT 21.315 12.960 21.635 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 16.040 21.230 16.360 ;
      LAYER met4 ;
        RECT 20.910 16.040 21.230 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 15.600 21.230 15.920 ;
      LAYER met4 ;
        RECT 20.910 15.600 21.230 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 15.160 21.230 15.480 ;
      LAYER met4 ;
        RECT 20.910 15.160 21.230 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 14.720 21.230 15.040 ;
      LAYER met4 ;
        RECT 20.910 14.720 21.230 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 14.280 21.230 14.600 ;
      LAYER met4 ;
        RECT 20.910 14.280 21.230 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 13.840 21.230 14.160 ;
      LAYER met4 ;
        RECT 20.910 13.840 21.230 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 13.400 21.230 13.720 ;
      LAYER met4 ;
        RECT 20.910 13.400 21.230 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.910 12.960 21.230 13.280 ;
      LAYER met4 ;
        RECT 20.910 12.960 21.230 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 16.040 20.825 16.360 ;
      LAYER met4 ;
        RECT 20.505 16.040 20.825 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 15.600 20.825 15.920 ;
      LAYER met4 ;
        RECT 20.505 15.600 20.825 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 15.160 20.825 15.480 ;
      LAYER met4 ;
        RECT 20.505 15.160 20.825 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 14.720 20.825 15.040 ;
      LAYER met4 ;
        RECT 20.505 14.720 20.825 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 14.280 20.825 14.600 ;
      LAYER met4 ;
        RECT 20.505 14.280 20.825 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 13.840 20.825 14.160 ;
      LAYER met4 ;
        RECT 20.505 13.840 20.825 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 13.400 20.825 13.720 ;
      LAYER met4 ;
        RECT 20.505 13.400 20.825 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.505 12.960 20.825 13.280 ;
      LAYER met4 ;
        RECT 20.505 12.960 20.825 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 16.040 20.420 16.360 ;
      LAYER met4 ;
        RECT 20.100 16.040 20.420 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 15.600 20.420 15.920 ;
      LAYER met4 ;
        RECT 20.100 15.600 20.420 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 15.160 20.420 15.480 ;
      LAYER met4 ;
        RECT 20.100 15.160 20.420 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 14.720 20.420 15.040 ;
      LAYER met4 ;
        RECT 20.100 14.720 20.420 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 14.280 20.420 14.600 ;
      LAYER met4 ;
        RECT 20.100 14.280 20.420 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 13.840 20.420 14.160 ;
      LAYER met4 ;
        RECT 20.100 13.840 20.420 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 13.400 20.420 13.720 ;
      LAYER met4 ;
        RECT 20.100 13.400 20.420 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.100 12.960 20.420 13.280 ;
      LAYER met4 ;
        RECT 20.100 12.960 20.420 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 16.040 20.015 16.360 ;
      LAYER met4 ;
        RECT 19.695 16.040 20.015 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 15.600 20.015 15.920 ;
      LAYER met4 ;
        RECT 19.695 15.600 20.015 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 15.160 20.015 15.480 ;
      LAYER met4 ;
        RECT 19.695 15.160 20.015 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 14.720 20.015 15.040 ;
      LAYER met4 ;
        RECT 19.695 14.720 20.015 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 14.280 20.015 14.600 ;
      LAYER met4 ;
        RECT 19.695 14.280 20.015 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 13.840 20.015 14.160 ;
      LAYER met4 ;
        RECT 19.695 13.840 20.015 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 13.400 20.015 13.720 ;
      LAYER met4 ;
        RECT 19.695 13.400 20.015 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 12.960 20.015 13.280 ;
      LAYER met4 ;
        RECT 19.695 12.960 20.015 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 16.040 19.610 16.360 ;
      LAYER met4 ;
        RECT 19.290 16.040 19.610 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 15.600 19.610 15.920 ;
      LAYER met4 ;
        RECT 19.290 15.600 19.610 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 15.160 19.610 15.480 ;
      LAYER met4 ;
        RECT 19.290 15.160 19.610 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 14.720 19.610 15.040 ;
      LAYER met4 ;
        RECT 19.290 14.720 19.610 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 14.280 19.610 14.600 ;
      LAYER met4 ;
        RECT 19.290 14.280 19.610 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 13.840 19.610 14.160 ;
      LAYER met4 ;
        RECT 19.290 13.840 19.610 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 13.400 19.610 13.720 ;
      LAYER met4 ;
        RECT 19.290 13.400 19.610 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.290 12.960 19.610 13.280 ;
      LAYER met4 ;
        RECT 19.290 12.960 19.610 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 16.040 19.205 16.360 ;
      LAYER met4 ;
        RECT 18.885 16.040 19.205 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 15.600 19.205 15.920 ;
      LAYER met4 ;
        RECT 18.885 15.600 19.205 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 15.160 19.205 15.480 ;
      LAYER met4 ;
        RECT 18.885 15.160 19.205 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 14.720 19.205 15.040 ;
      LAYER met4 ;
        RECT 18.885 14.720 19.205 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 14.280 19.205 14.600 ;
      LAYER met4 ;
        RECT 18.885 14.280 19.205 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 13.840 19.205 14.160 ;
      LAYER met4 ;
        RECT 18.885 13.840 19.205 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 13.400 19.205 13.720 ;
      LAYER met4 ;
        RECT 18.885 13.400 19.205 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.885 12.960 19.205 13.280 ;
      LAYER met4 ;
        RECT 18.885 12.960 19.205 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 16.040 18.800 16.360 ;
      LAYER met4 ;
        RECT 18.480 16.040 18.800 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 15.600 18.800 15.920 ;
      LAYER met4 ;
        RECT 18.480 15.600 18.800 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 15.160 18.800 15.480 ;
      LAYER met4 ;
        RECT 18.480 15.160 18.800 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 14.720 18.800 15.040 ;
      LAYER met4 ;
        RECT 18.480 14.720 18.800 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 14.280 18.800 14.600 ;
      LAYER met4 ;
        RECT 18.480 14.280 18.800 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 13.840 18.800 14.160 ;
      LAYER met4 ;
        RECT 18.480 13.840 18.800 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 13.400 18.800 13.720 ;
      LAYER met4 ;
        RECT 18.480 13.400 18.800 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.480 12.960 18.800 13.280 ;
      LAYER met4 ;
        RECT 18.480 12.960 18.800 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 16.040 18.395 16.360 ;
      LAYER met4 ;
        RECT 18.075 16.040 18.395 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 15.600 18.395 15.920 ;
      LAYER met4 ;
        RECT 18.075 15.600 18.395 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 15.160 18.395 15.480 ;
      LAYER met4 ;
        RECT 18.075 15.160 18.395 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 14.720 18.395 15.040 ;
      LAYER met4 ;
        RECT 18.075 14.720 18.395 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 14.280 18.395 14.600 ;
      LAYER met4 ;
        RECT 18.075 14.280 18.395 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 13.840 18.395 14.160 ;
      LAYER met4 ;
        RECT 18.075 13.840 18.395 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 13.400 18.395 13.720 ;
      LAYER met4 ;
        RECT 18.075 13.400 18.395 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.075 12.960 18.395 13.280 ;
      LAYER met4 ;
        RECT 18.075 12.960 18.395 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 16.040 17.990 16.360 ;
      LAYER met4 ;
        RECT 17.670 16.040 17.990 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 15.600 17.990 15.920 ;
      LAYER met4 ;
        RECT 17.670 15.600 17.990 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 15.160 17.990 15.480 ;
      LAYER met4 ;
        RECT 17.670 15.160 17.990 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 14.720 17.990 15.040 ;
      LAYER met4 ;
        RECT 17.670 14.720 17.990 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 14.280 17.990 14.600 ;
      LAYER met4 ;
        RECT 17.670 14.280 17.990 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 13.840 17.990 14.160 ;
      LAYER met4 ;
        RECT 17.670 13.840 17.990 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 13.400 17.990 13.720 ;
      LAYER met4 ;
        RECT 17.670 13.400 17.990 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.670 12.960 17.990 13.280 ;
      LAYER met4 ;
        RECT 17.670 12.960 17.990 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 16.040 17.585 16.360 ;
      LAYER met4 ;
        RECT 17.265 16.040 17.585 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 15.600 17.585 15.920 ;
      LAYER met4 ;
        RECT 17.265 15.600 17.585 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 15.160 17.585 15.480 ;
      LAYER met4 ;
        RECT 17.265 15.160 17.585 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 14.720 17.585 15.040 ;
      LAYER met4 ;
        RECT 17.265 14.720 17.585 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 14.280 17.585 14.600 ;
      LAYER met4 ;
        RECT 17.265 14.280 17.585 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 13.840 17.585 14.160 ;
      LAYER met4 ;
        RECT 17.265 13.840 17.585 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 13.400 17.585 13.720 ;
      LAYER met4 ;
        RECT 17.265 13.400 17.585 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.265 12.960 17.585 13.280 ;
      LAYER met4 ;
        RECT 17.265 12.960 17.585 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 16.040 17.180 16.360 ;
      LAYER met4 ;
        RECT 16.860 16.040 17.180 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 15.600 17.180 15.920 ;
      LAYER met4 ;
        RECT 16.860 15.600 17.180 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 15.160 17.180 15.480 ;
      LAYER met4 ;
        RECT 16.860 15.160 17.180 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 14.720 17.180 15.040 ;
      LAYER met4 ;
        RECT 16.860 14.720 17.180 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 14.280 17.180 14.600 ;
      LAYER met4 ;
        RECT 16.860 14.280 17.180 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 13.840 17.180 14.160 ;
      LAYER met4 ;
        RECT 16.860 13.840 17.180 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 13.400 17.180 13.720 ;
      LAYER met4 ;
        RECT 16.860 13.400 17.180 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.860 12.960 17.180 13.280 ;
      LAYER met4 ;
        RECT 16.860 12.960 17.180 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 16.040 16.775 16.360 ;
      LAYER met4 ;
        RECT 16.455 16.040 16.775 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 15.600 16.775 15.920 ;
      LAYER met4 ;
        RECT 16.455 15.600 16.775 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 15.160 16.775 15.480 ;
      LAYER met4 ;
        RECT 16.455 15.160 16.775 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 14.720 16.775 15.040 ;
      LAYER met4 ;
        RECT 16.455 14.720 16.775 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 14.280 16.775 14.600 ;
      LAYER met4 ;
        RECT 16.455 14.280 16.775 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 13.840 16.775 14.160 ;
      LAYER met4 ;
        RECT 16.455 13.840 16.775 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 13.400 16.775 13.720 ;
      LAYER met4 ;
        RECT 16.455 13.400 16.775 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 12.960 16.775 13.280 ;
      LAYER met4 ;
        RECT 16.455 12.960 16.775 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 16.040 16.370 16.360 ;
      LAYER met4 ;
        RECT 16.050 16.040 16.370 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 15.600 16.370 15.920 ;
      LAYER met4 ;
        RECT 16.050 15.600 16.370 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 15.160 16.370 15.480 ;
      LAYER met4 ;
        RECT 16.050 15.160 16.370 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 14.720 16.370 15.040 ;
      LAYER met4 ;
        RECT 16.050 14.720 16.370 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 14.280 16.370 14.600 ;
      LAYER met4 ;
        RECT 16.050 14.280 16.370 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 13.840 16.370 14.160 ;
      LAYER met4 ;
        RECT 16.050 13.840 16.370 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 13.400 16.370 13.720 ;
      LAYER met4 ;
        RECT 16.050 13.400 16.370 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.050 12.960 16.370 13.280 ;
      LAYER met4 ;
        RECT 16.050 12.960 16.370 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 16.040 15.965 16.360 ;
      LAYER met4 ;
        RECT 15.645 16.040 15.965 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 15.600 15.965 15.920 ;
      LAYER met4 ;
        RECT 15.645 15.600 15.965 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 15.160 15.965 15.480 ;
      LAYER met4 ;
        RECT 15.645 15.160 15.965 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 14.720 15.965 15.040 ;
      LAYER met4 ;
        RECT 15.645 14.720 15.965 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 14.280 15.965 14.600 ;
      LAYER met4 ;
        RECT 15.645 14.280 15.965 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 13.840 15.965 14.160 ;
      LAYER met4 ;
        RECT 15.645 13.840 15.965 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 13.400 15.965 13.720 ;
      LAYER met4 ;
        RECT 15.645 13.400 15.965 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 12.960 15.965 13.280 ;
      LAYER met4 ;
        RECT 15.645 12.960 15.965 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 16.040 15.560 16.360 ;
      LAYER met4 ;
        RECT 15.240 16.040 15.560 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 15.600 15.560 15.920 ;
      LAYER met4 ;
        RECT 15.240 15.600 15.560 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 15.160 15.560 15.480 ;
      LAYER met4 ;
        RECT 15.240 15.160 15.560 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 14.720 15.560 15.040 ;
      LAYER met4 ;
        RECT 15.240 14.720 15.560 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 14.280 15.560 14.600 ;
      LAYER met4 ;
        RECT 15.240 14.280 15.560 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 13.840 15.560 14.160 ;
      LAYER met4 ;
        RECT 15.240 13.840 15.560 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 13.400 15.560 13.720 ;
      LAYER met4 ;
        RECT 15.240 13.400 15.560 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.240 12.960 15.560 13.280 ;
      LAYER met4 ;
        RECT 15.240 12.960 15.560 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 16.040 15.155 16.360 ;
      LAYER met4 ;
        RECT 14.835 16.040 15.155 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 15.600 15.155 15.920 ;
      LAYER met4 ;
        RECT 14.835 15.600 15.155 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 15.160 15.155 15.480 ;
      LAYER met4 ;
        RECT 14.835 15.160 15.155 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 14.720 15.155 15.040 ;
      LAYER met4 ;
        RECT 14.835 14.720 15.155 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 14.280 15.155 14.600 ;
      LAYER met4 ;
        RECT 14.835 14.280 15.155 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 13.840 15.155 14.160 ;
      LAYER met4 ;
        RECT 14.835 13.840 15.155 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 13.400 15.155 13.720 ;
      LAYER met4 ;
        RECT 14.835 13.400 15.155 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.835 12.960 15.155 13.280 ;
      LAYER met4 ;
        RECT 14.835 12.960 15.155 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 16.040 14.750 16.360 ;
      LAYER met4 ;
        RECT 14.430 16.040 14.750 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 15.600 14.750 15.920 ;
      LAYER met4 ;
        RECT 14.430 15.600 14.750 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 15.160 14.750 15.480 ;
      LAYER met4 ;
        RECT 14.430 15.160 14.750 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 14.720 14.750 15.040 ;
      LAYER met4 ;
        RECT 14.430 14.720 14.750 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 14.280 14.750 14.600 ;
      LAYER met4 ;
        RECT 14.430 14.280 14.750 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 13.840 14.750 14.160 ;
      LAYER met4 ;
        RECT 14.430 13.840 14.750 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 13.400 14.750 13.720 ;
      LAYER met4 ;
        RECT 14.430 13.400 14.750 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.430 12.960 14.750 13.280 ;
      LAYER met4 ;
        RECT 14.430 12.960 14.750 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 16.040 14.345 16.360 ;
      LAYER met4 ;
        RECT 14.025 16.040 14.345 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 15.600 14.345 15.920 ;
      LAYER met4 ;
        RECT 14.025 15.600 14.345 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 15.160 14.345 15.480 ;
      LAYER met4 ;
        RECT 14.025 15.160 14.345 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 14.720 14.345 15.040 ;
      LAYER met4 ;
        RECT 14.025 14.720 14.345 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 14.280 14.345 14.600 ;
      LAYER met4 ;
        RECT 14.025 14.280 14.345 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 13.840 14.345 14.160 ;
      LAYER met4 ;
        RECT 14.025 13.840 14.345 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 13.400 14.345 13.720 ;
      LAYER met4 ;
        RECT 14.025 13.400 14.345 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.025 12.960 14.345 13.280 ;
      LAYER met4 ;
        RECT 14.025 12.960 14.345 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 16.040 13.940 16.360 ;
      LAYER met4 ;
        RECT 13.620 16.040 13.940 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 15.600 13.940 15.920 ;
      LAYER met4 ;
        RECT 13.620 15.600 13.940 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 15.160 13.940 15.480 ;
      LAYER met4 ;
        RECT 13.620 15.160 13.940 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 14.720 13.940 15.040 ;
      LAYER met4 ;
        RECT 13.620 14.720 13.940 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 14.280 13.940 14.600 ;
      LAYER met4 ;
        RECT 13.620 14.280 13.940 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 13.840 13.940 14.160 ;
      LAYER met4 ;
        RECT 13.620 13.840 13.940 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 13.400 13.940 13.720 ;
      LAYER met4 ;
        RECT 13.620 13.400 13.940 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.620 12.960 13.940 13.280 ;
      LAYER met4 ;
        RECT 13.620 12.960 13.940 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 16.040 13.535 16.360 ;
      LAYER met4 ;
        RECT 13.215 16.040 13.535 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 15.600 13.535 15.920 ;
      LAYER met4 ;
        RECT 13.215 15.600 13.535 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 15.160 13.535 15.480 ;
      LAYER met4 ;
        RECT 13.215 15.160 13.535 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 14.720 13.535 15.040 ;
      LAYER met4 ;
        RECT 13.215 14.720 13.535 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 14.280 13.535 14.600 ;
      LAYER met4 ;
        RECT 13.215 14.280 13.535 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 13.840 13.535 14.160 ;
      LAYER met4 ;
        RECT 13.215 13.840 13.535 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 13.400 13.535 13.720 ;
      LAYER met4 ;
        RECT 13.215 13.400 13.535 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.215 12.960 13.535 13.280 ;
      LAYER met4 ;
        RECT 13.215 12.960 13.535 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 16.040 13.130 16.360 ;
      LAYER met4 ;
        RECT 12.810 16.040 13.130 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 15.600 13.130 15.920 ;
      LAYER met4 ;
        RECT 12.810 15.600 13.130 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 15.160 13.130 15.480 ;
      LAYER met4 ;
        RECT 12.810 15.160 13.130 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 14.720 13.130 15.040 ;
      LAYER met4 ;
        RECT 12.810 14.720 13.130 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 14.280 13.130 14.600 ;
      LAYER met4 ;
        RECT 12.810 14.280 13.130 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 13.840 13.130 14.160 ;
      LAYER met4 ;
        RECT 12.810 13.840 13.130 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 13.400 13.130 13.720 ;
      LAYER met4 ;
        RECT 12.810 13.400 13.130 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.810 12.960 13.130 13.280 ;
      LAYER met4 ;
        RECT 12.810 12.960 13.130 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 16.040 12.725 16.360 ;
      LAYER met4 ;
        RECT 12.405 16.040 12.725 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 15.600 12.725 15.920 ;
      LAYER met4 ;
        RECT 12.405 15.600 12.725 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 15.160 12.725 15.480 ;
      LAYER met4 ;
        RECT 12.405 15.160 12.725 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 14.720 12.725 15.040 ;
      LAYER met4 ;
        RECT 12.405 14.720 12.725 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 14.280 12.725 14.600 ;
      LAYER met4 ;
        RECT 12.405 14.280 12.725 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 13.840 12.725 14.160 ;
      LAYER met4 ;
        RECT 12.405 13.840 12.725 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 13.400 12.725 13.720 ;
      LAYER met4 ;
        RECT 12.405 13.400 12.725 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.405 12.960 12.725 13.280 ;
      LAYER met4 ;
        RECT 12.405 12.960 12.725 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 16.040 12.320 16.360 ;
      LAYER met4 ;
        RECT 12.000 16.040 12.320 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 15.600 12.320 15.920 ;
      LAYER met4 ;
        RECT 12.000 15.600 12.320 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 15.160 12.320 15.480 ;
      LAYER met4 ;
        RECT 12.000 15.160 12.320 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 14.720 12.320 15.040 ;
      LAYER met4 ;
        RECT 12.000 14.720 12.320 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 14.280 12.320 14.600 ;
      LAYER met4 ;
        RECT 12.000 14.280 12.320 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 13.840 12.320 14.160 ;
      LAYER met4 ;
        RECT 12.000 13.840 12.320 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 13.400 12.320 13.720 ;
      LAYER met4 ;
        RECT 12.000 13.400 12.320 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.000 12.960 12.320 13.280 ;
      LAYER met4 ;
        RECT 12.000 12.960 12.320 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 16.040 11.915 16.360 ;
      LAYER met4 ;
        RECT 11.595 16.040 11.915 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 15.600 11.915 15.920 ;
      LAYER met4 ;
        RECT 11.595 15.600 11.915 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 15.160 11.915 15.480 ;
      LAYER met4 ;
        RECT 11.595 15.160 11.915 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 14.720 11.915 15.040 ;
      LAYER met4 ;
        RECT 11.595 14.720 11.915 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 14.280 11.915 14.600 ;
      LAYER met4 ;
        RECT 11.595 14.280 11.915 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 13.840 11.915 14.160 ;
      LAYER met4 ;
        RECT 11.595 13.840 11.915 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 13.400 11.915 13.720 ;
      LAYER met4 ;
        RECT 11.595 13.400 11.915 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.595 12.960 11.915 13.280 ;
      LAYER met4 ;
        RECT 11.595 12.960 11.915 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 16.040 11.510 16.360 ;
      LAYER met4 ;
        RECT 11.190 16.040 11.510 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 15.600 11.510 15.920 ;
      LAYER met4 ;
        RECT 11.190 15.600 11.510 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 15.160 11.510 15.480 ;
      LAYER met4 ;
        RECT 11.190 15.160 11.510 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 14.720 11.510 15.040 ;
      LAYER met4 ;
        RECT 11.190 14.720 11.510 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 14.280 11.510 14.600 ;
      LAYER met4 ;
        RECT 11.190 14.280 11.510 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 13.840 11.510 14.160 ;
      LAYER met4 ;
        RECT 11.190 13.840 11.510 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 13.400 11.510 13.720 ;
      LAYER met4 ;
        RECT 11.190 13.400 11.510 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.190 12.960 11.510 13.280 ;
      LAYER met4 ;
        RECT 11.190 12.960 11.510 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 16.040 11.105 16.360 ;
      LAYER met4 ;
        RECT 10.785 16.040 11.105 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 15.600 11.105 15.920 ;
      LAYER met4 ;
        RECT 10.785 15.600 11.105 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 15.160 11.105 15.480 ;
      LAYER met4 ;
        RECT 10.785 15.160 11.105 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 14.720 11.105 15.040 ;
      LAYER met4 ;
        RECT 10.785 14.720 11.105 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 14.280 11.105 14.600 ;
      LAYER met4 ;
        RECT 10.785 14.280 11.105 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 13.840 11.105 14.160 ;
      LAYER met4 ;
        RECT 10.785 13.840 11.105 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 13.400 11.105 13.720 ;
      LAYER met4 ;
        RECT 10.785 13.400 11.105 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 12.960 11.105 13.280 ;
      LAYER met4 ;
        RECT 10.785 12.960 11.105 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 16.040 10.700 16.360 ;
      LAYER met4 ;
        RECT 10.380 16.040 10.700 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 15.600 10.700 15.920 ;
      LAYER met4 ;
        RECT 10.380 15.600 10.700 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 15.160 10.700 15.480 ;
      LAYER met4 ;
        RECT 10.380 15.160 10.700 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 14.720 10.700 15.040 ;
      LAYER met4 ;
        RECT 10.380 14.720 10.700 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 14.280 10.700 14.600 ;
      LAYER met4 ;
        RECT 10.380 14.280 10.700 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 13.840 10.700 14.160 ;
      LAYER met4 ;
        RECT 10.380 13.840 10.700 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 13.400 10.700 13.720 ;
      LAYER met4 ;
        RECT 10.380 13.400 10.700 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.380 12.960 10.700 13.280 ;
      LAYER met4 ;
        RECT 10.380 12.960 10.700 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 16.040 10.295 16.360 ;
      LAYER met4 ;
        RECT 9.975 16.040 10.295 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 15.600 10.295 15.920 ;
      LAYER met4 ;
        RECT 9.975 15.600 10.295 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 15.160 10.295 15.480 ;
      LAYER met4 ;
        RECT 9.975 15.160 10.295 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 14.720 10.295 15.040 ;
      LAYER met4 ;
        RECT 9.975 14.720 10.295 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 14.280 10.295 14.600 ;
      LAYER met4 ;
        RECT 9.975 14.280 10.295 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 13.840 10.295 14.160 ;
      LAYER met4 ;
        RECT 9.975 13.840 10.295 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 13.400 10.295 13.720 ;
      LAYER met4 ;
        RECT 9.975 13.400 10.295 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.975 12.960 10.295 13.280 ;
      LAYER met4 ;
        RECT 9.975 12.960 10.295 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 16.040 9.890 16.360 ;
      LAYER met4 ;
        RECT 9.570 16.040 9.890 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 15.600 9.890 15.920 ;
      LAYER met4 ;
        RECT 9.570 15.600 9.890 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 15.160 9.890 15.480 ;
      LAYER met4 ;
        RECT 9.570 15.160 9.890 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 14.720 9.890 15.040 ;
      LAYER met4 ;
        RECT 9.570 14.720 9.890 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 14.280 9.890 14.600 ;
      LAYER met4 ;
        RECT 9.570 14.280 9.890 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 13.840 9.890 14.160 ;
      LAYER met4 ;
        RECT 9.570 13.840 9.890 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 13.400 9.890 13.720 ;
      LAYER met4 ;
        RECT 9.570 13.400 9.890 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.570 12.960 9.890 13.280 ;
      LAYER met4 ;
        RECT 9.570 12.960 9.890 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 16.040 9.485 16.360 ;
      LAYER met4 ;
        RECT 9.165 16.040 9.485 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 15.600 9.485 15.920 ;
      LAYER met4 ;
        RECT 9.165 15.600 9.485 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 15.160 9.485 15.480 ;
      LAYER met4 ;
        RECT 9.165 15.160 9.485 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 14.720 9.485 15.040 ;
      LAYER met4 ;
        RECT 9.165 14.720 9.485 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 14.280 9.485 14.600 ;
      LAYER met4 ;
        RECT 9.165 14.280 9.485 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 13.840 9.485 14.160 ;
      LAYER met4 ;
        RECT 9.165 13.840 9.485 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 13.400 9.485 13.720 ;
      LAYER met4 ;
        RECT 9.165 13.400 9.485 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.165 12.960 9.485 13.280 ;
      LAYER met4 ;
        RECT 9.165 12.960 9.485 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 16.040 9.080 16.360 ;
      LAYER met4 ;
        RECT 8.760 16.040 9.080 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 15.600 9.080 15.920 ;
      LAYER met4 ;
        RECT 8.760 15.600 9.080 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 15.160 9.080 15.480 ;
      LAYER met4 ;
        RECT 8.760 15.160 9.080 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 14.720 9.080 15.040 ;
      LAYER met4 ;
        RECT 8.760 14.720 9.080 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 14.280 9.080 14.600 ;
      LAYER met4 ;
        RECT 8.760 14.280 9.080 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 13.840 9.080 14.160 ;
      LAYER met4 ;
        RECT 8.760 13.840 9.080 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 13.400 9.080 13.720 ;
      LAYER met4 ;
        RECT 8.760 13.400 9.080 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.760 12.960 9.080 13.280 ;
      LAYER met4 ;
        RECT 8.760 12.960 9.080 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 16.040 8.675 16.360 ;
      LAYER met4 ;
        RECT 8.355 16.040 8.675 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 15.600 8.675 15.920 ;
      LAYER met4 ;
        RECT 8.355 15.600 8.675 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 15.160 8.675 15.480 ;
      LAYER met4 ;
        RECT 8.355 15.160 8.675 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 14.720 8.675 15.040 ;
      LAYER met4 ;
        RECT 8.355 14.720 8.675 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 14.280 8.675 14.600 ;
      LAYER met4 ;
        RECT 8.355 14.280 8.675 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 13.840 8.675 14.160 ;
      LAYER met4 ;
        RECT 8.355 13.840 8.675 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 13.400 8.675 13.720 ;
      LAYER met4 ;
        RECT 8.355 13.400 8.675 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.355 12.960 8.675 13.280 ;
      LAYER met4 ;
        RECT 8.355 12.960 8.675 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 16.040 8.270 16.360 ;
      LAYER met4 ;
        RECT 7.950 16.040 8.270 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 15.600 8.270 15.920 ;
      LAYER met4 ;
        RECT 7.950 15.600 8.270 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 15.160 8.270 15.480 ;
      LAYER met4 ;
        RECT 7.950 15.160 8.270 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 14.720 8.270 15.040 ;
      LAYER met4 ;
        RECT 7.950 14.720 8.270 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 14.280 8.270 14.600 ;
      LAYER met4 ;
        RECT 7.950 14.280 8.270 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 13.840 8.270 14.160 ;
      LAYER met4 ;
        RECT 7.950 13.840 8.270 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 13.400 8.270 13.720 ;
      LAYER met4 ;
        RECT 7.950 13.400 8.270 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.950 12.960 8.270 13.280 ;
      LAYER met4 ;
        RECT 7.950 12.960 8.270 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 16.040 7.865 16.360 ;
      LAYER met4 ;
        RECT 7.545 16.040 7.865 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 15.600 7.865 15.920 ;
      LAYER met4 ;
        RECT 7.545 15.600 7.865 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 15.160 7.865 15.480 ;
      LAYER met4 ;
        RECT 7.545 15.160 7.865 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 14.720 7.865 15.040 ;
      LAYER met4 ;
        RECT 7.545 14.720 7.865 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 14.280 7.865 14.600 ;
      LAYER met4 ;
        RECT 7.545 14.280 7.865 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 13.840 7.865 14.160 ;
      LAYER met4 ;
        RECT 7.545 13.840 7.865 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 13.400 7.865 13.720 ;
      LAYER met4 ;
        RECT 7.545 13.400 7.865 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.545 12.960 7.865 13.280 ;
      LAYER met4 ;
        RECT 7.545 12.960 7.865 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 16.040 7.460 16.360 ;
      LAYER met4 ;
        RECT 7.140 16.040 7.460 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 15.600 7.460 15.920 ;
      LAYER met4 ;
        RECT 7.140 15.600 7.460 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 15.160 7.460 15.480 ;
      LAYER met4 ;
        RECT 7.140 15.160 7.460 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 14.720 7.460 15.040 ;
      LAYER met4 ;
        RECT 7.140 14.720 7.460 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 14.280 7.460 14.600 ;
      LAYER met4 ;
        RECT 7.140 14.280 7.460 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 13.840 7.460 14.160 ;
      LAYER met4 ;
        RECT 7.140 13.840 7.460 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 13.400 7.460 13.720 ;
      LAYER met4 ;
        RECT 7.140 13.400 7.460 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.140 12.960 7.460 13.280 ;
      LAYER met4 ;
        RECT 7.140 12.960 7.460 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 16.040 7.055 16.360 ;
      LAYER met4 ;
        RECT 6.735 16.040 7.055 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 15.600 7.055 15.920 ;
      LAYER met4 ;
        RECT 6.735 15.600 7.055 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 15.160 7.055 15.480 ;
      LAYER met4 ;
        RECT 6.735 15.160 7.055 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 14.720 7.055 15.040 ;
      LAYER met4 ;
        RECT 6.735 14.720 7.055 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 14.280 7.055 14.600 ;
      LAYER met4 ;
        RECT 6.735 14.280 7.055 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 13.840 7.055 14.160 ;
      LAYER met4 ;
        RECT 6.735 13.840 7.055 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 13.400 7.055 13.720 ;
      LAYER met4 ;
        RECT 6.735 13.400 7.055 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.735 12.960 7.055 13.280 ;
      LAYER met4 ;
        RECT 6.735 12.960 7.055 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 16.040 6.650 16.360 ;
      LAYER met4 ;
        RECT 6.330 16.040 6.650 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 15.600 6.650 15.920 ;
      LAYER met4 ;
        RECT 6.330 15.600 6.650 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 15.160 6.650 15.480 ;
      LAYER met4 ;
        RECT 6.330 15.160 6.650 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 14.720 6.650 15.040 ;
      LAYER met4 ;
        RECT 6.330 14.720 6.650 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 14.280 6.650 14.600 ;
      LAYER met4 ;
        RECT 6.330 14.280 6.650 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 13.840 6.650 14.160 ;
      LAYER met4 ;
        RECT 6.330 13.840 6.650 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 13.400 6.650 13.720 ;
      LAYER met4 ;
        RECT 6.330 13.400 6.650 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.330 12.960 6.650 13.280 ;
      LAYER met4 ;
        RECT 6.330 12.960 6.650 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 16.040 6.245 16.360 ;
      LAYER met4 ;
        RECT 5.925 16.040 6.245 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 15.600 6.245 15.920 ;
      LAYER met4 ;
        RECT 5.925 15.600 6.245 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 15.160 6.245 15.480 ;
      LAYER met4 ;
        RECT 5.925 15.160 6.245 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 14.720 6.245 15.040 ;
      LAYER met4 ;
        RECT 5.925 14.720 6.245 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 14.280 6.245 14.600 ;
      LAYER met4 ;
        RECT 5.925 14.280 6.245 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 13.840 6.245 14.160 ;
      LAYER met4 ;
        RECT 5.925 13.840 6.245 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 13.400 6.245 13.720 ;
      LAYER met4 ;
        RECT 5.925 13.400 6.245 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.925 12.960 6.245 13.280 ;
      LAYER met4 ;
        RECT 5.925 12.960 6.245 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 16.040 5.840 16.360 ;
      LAYER met4 ;
        RECT 5.520 16.040 5.840 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 15.600 5.840 15.920 ;
      LAYER met4 ;
        RECT 5.520 15.600 5.840 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 15.160 5.840 15.480 ;
      LAYER met4 ;
        RECT 5.520 15.160 5.840 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 14.720 5.840 15.040 ;
      LAYER met4 ;
        RECT 5.520 14.720 5.840 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 14.280 5.840 14.600 ;
      LAYER met4 ;
        RECT 5.520 14.280 5.840 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 13.840 5.840 14.160 ;
      LAYER met4 ;
        RECT 5.520 13.840 5.840 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 13.400 5.840 13.720 ;
      LAYER met4 ;
        RECT 5.520 13.400 5.840 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 12.960 5.840 13.280 ;
      LAYER met4 ;
        RECT 5.520 12.960 5.840 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 16.040 5.435 16.360 ;
      LAYER met4 ;
        RECT 5.115 16.040 5.435 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 15.600 5.435 15.920 ;
      LAYER met4 ;
        RECT 5.115 15.600 5.435 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 15.160 5.435 15.480 ;
      LAYER met4 ;
        RECT 5.115 15.160 5.435 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 14.720 5.435 15.040 ;
      LAYER met4 ;
        RECT 5.115 14.720 5.435 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 14.280 5.435 14.600 ;
      LAYER met4 ;
        RECT 5.115 14.280 5.435 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 13.840 5.435 14.160 ;
      LAYER met4 ;
        RECT 5.115 13.840 5.435 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 13.400 5.435 13.720 ;
      LAYER met4 ;
        RECT 5.115 13.400 5.435 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.115 12.960 5.435 13.280 ;
      LAYER met4 ;
        RECT 5.115 12.960 5.435 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 16.040 5.030 16.360 ;
      LAYER met4 ;
        RECT 4.710 16.040 5.030 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 15.600 5.030 15.920 ;
      LAYER met4 ;
        RECT 4.710 15.600 5.030 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 15.160 5.030 15.480 ;
      LAYER met4 ;
        RECT 4.710 15.160 5.030 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 14.720 5.030 15.040 ;
      LAYER met4 ;
        RECT 4.710 14.720 5.030 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 14.280 5.030 14.600 ;
      LAYER met4 ;
        RECT 4.710 14.280 5.030 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 13.840 5.030 14.160 ;
      LAYER met4 ;
        RECT 4.710 13.840 5.030 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 13.400 5.030 13.720 ;
      LAYER met4 ;
        RECT 4.710 13.400 5.030 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.710 12.960 5.030 13.280 ;
      LAYER met4 ;
        RECT 4.710 12.960 5.030 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 16.040 4.625 16.360 ;
      LAYER met4 ;
        RECT 4.305 16.040 4.625 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 15.600 4.625 15.920 ;
      LAYER met4 ;
        RECT 4.305 15.600 4.625 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 15.160 4.625 15.480 ;
      LAYER met4 ;
        RECT 4.305 15.160 4.625 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 14.720 4.625 15.040 ;
      LAYER met4 ;
        RECT 4.305 14.720 4.625 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 14.280 4.625 14.600 ;
      LAYER met4 ;
        RECT 4.305 14.280 4.625 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 13.840 4.625 14.160 ;
      LAYER met4 ;
        RECT 4.305 13.840 4.625 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 13.400 4.625 13.720 ;
      LAYER met4 ;
        RECT 4.305 13.400 4.625 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.305 12.960 4.625 13.280 ;
      LAYER met4 ;
        RECT 4.305 12.960 4.625 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 16.040 4.220 16.360 ;
      LAYER met4 ;
        RECT 3.900 16.040 4.220 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 15.600 4.220 15.920 ;
      LAYER met4 ;
        RECT 3.900 15.600 4.220 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 15.160 4.220 15.480 ;
      LAYER met4 ;
        RECT 3.900 15.160 4.220 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 14.720 4.220 15.040 ;
      LAYER met4 ;
        RECT 3.900 14.720 4.220 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 14.280 4.220 14.600 ;
      LAYER met4 ;
        RECT 3.900 14.280 4.220 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 13.840 4.220 14.160 ;
      LAYER met4 ;
        RECT 3.900 13.840 4.220 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 13.400 4.220 13.720 ;
      LAYER met4 ;
        RECT 3.900 13.400 4.220 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.900 12.960 4.220 13.280 ;
      LAYER met4 ;
        RECT 3.900 12.960 4.220 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 16.040 3.815 16.360 ;
      LAYER met4 ;
        RECT 3.495 16.040 3.815 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 15.600 3.815 15.920 ;
      LAYER met4 ;
        RECT 3.495 15.600 3.815 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 15.160 3.815 15.480 ;
      LAYER met4 ;
        RECT 3.495 15.160 3.815 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 14.720 3.815 15.040 ;
      LAYER met4 ;
        RECT 3.495 14.720 3.815 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 14.280 3.815 14.600 ;
      LAYER met4 ;
        RECT 3.495 14.280 3.815 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 13.840 3.815 14.160 ;
      LAYER met4 ;
        RECT 3.495 13.840 3.815 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 13.400 3.815 13.720 ;
      LAYER met4 ;
        RECT 3.495 13.400 3.815 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.495 12.960 3.815 13.280 ;
      LAYER met4 ;
        RECT 3.495 12.960 3.815 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 16.040 3.410 16.360 ;
      LAYER met4 ;
        RECT 3.090 16.040 3.410 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 15.600 3.410 15.920 ;
      LAYER met4 ;
        RECT 3.090 15.600 3.410 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 15.160 3.410 15.480 ;
      LAYER met4 ;
        RECT 3.090 15.160 3.410 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 14.720 3.410 15.040 ;
      LAYER met4 ;
        RECT 3.090 14.720 3.410 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 14.280 3.410 14.600 ;
      LAYER met4 ;
        RECT 3.090 14.280 3.410 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 13.840 3.410 14.160 ;
      LAYER met4 ;
        RECT 3.090 13.840 3.410 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 13.400 3.410 13.720 ;
      LAYER met4 ;
        RECT 3.090 13.400 3.410 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.090 12.960 3.410 13.280 ;
      LAYER met4 ;
        RECT 3.090 12.960 3.410 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 16.040 3.000 16.360 ;
      LAYER met4 ;
        RECT 2.680 16.040 3.000 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 15.600 3.000 15.920 ;
      LAYER met4 ;
        RECT 2.680 15.600 3.000 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 15.160 3.000 15.480 ;
      LAYER met4 ;
        RECT 2.680 15.160 3.000 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 14.720 3.000 15.040 ;
      LAYER met4 ;
        RECT 2.680 14.720 3.000 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 14.280 3.000 14.600 ;
      LAYER met4 ;
        RECT 2.680 14.280 3.000 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 13.840 3.000 14.160 ;
      LAYER met4 ;
        RECT 2.680 13.840 3.000 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 13.400 3.000 13.720 ;
      LAYER met4 ;
        RECT 2.680 13.400 3.000 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 12.960 3.000 13.280 ;
      LAYER met4 ;
        RECT 2.680 12.960 3.000 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 16.040 2.590 16.360 ;
      LAYER met4 ;
        RECT 2.270 16.040 2.590 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 15.600 2.590 15.920 ;
      LAYER met4 ;
        RECT 2.270 15.600 2.590 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 15.160 2.590 15.480 ;
      LAYER met4 ;
        RECT 2.270 15.160 2.590 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 14.720 2.590 15.040 ;
      LAYER met4 ;
        RECT 2.270 14.720 2.590 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 14.280 2.590 14.600 ;
      LAYER met4 ;
        RECT 2.270 14.280 2.590 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 13.840 2.590 14.160 ;
      LAYER met4 ;
        RECT 2.270 13.840 2.590 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 13.400 2.590 13.720 ;
      LAYER met4 ;
        RECT 2.270 13.400 2.590 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.270 12.960 2.590 13.280 ;
      LAYER met4 ;
        RECT 2.270 12.960 2.590 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 16.040 2.180 16.360 ;
      LAYER met4 ;
        RECT 1.860 16.040 2.180 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 15.600 2.180 15.920 ;
      LAYER met4 ;
        RECT 1.860 15.600 2.180 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 15.160 2.180 15.480 ;
      LAYER met4 ;
        RECT 1.860 15.160 2.180 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 14.720 2.180 15.040 ;
      LAYER met4 ;
        RECT 1.860 14.720 2.180 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 14.280 2.180 14.600 ;
      LAYER met4 ;
        RECT 1.860 14.280 2.180 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 13.840 2.180 14.160 ;
      LAYER met4 ;
        RECT 1.860 13.840 2.180 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 13.400 2.180 13.720 ;
      LAYER met4 ;
        RECT 1.860 13.400 2.180 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.860 12.960 2.180 13.280 ;
      LAYER met4 ;
        RECT 1.860 12.960 2.180 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 16.040 1.770 16.360 ;
      LAYER met4 ;
        RECT 1.450 16.040 1.770 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 15.600 1.770 15.920 ;
      LAYER met4 ;
        RECT 1.450 15.600 1.770 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 15.160 1.770 15.480 ;
      LAYER met4 ;
        RECT 1.450 15.160 1.770 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 14.720 1.770 15.040 ;
      LAYER met4 ;
        RECT 1.450 14.720 1.770 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 14.280 1.770 14.600 ;
      LAYER met4 ;
        RECT 1.450 14.280 1.770 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 13.840 1.770 14.160 ;
      LAYER met4 ;
        RECT 1.450 13.840 1.770 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 13.400 1.770 13.720 ;
      LAYER met4 ;
        RECT 1.450 13.400 1.770 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.450 12.960 1.770 13.280 ;
      LAYER met4 ;
        RECT 1.450 12.960 1.770 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 16.040 1.360 16.360 ;
      LAYER met4 ;
        RECT 1.040 16.040 1.360 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 15.600 1.360 15.920 ;
      LAYER met4 ;
        RECT 1.040 15.600 1.360 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 15.160 1.360 15.480 ;
      LAYER met4 ;
        RECT 1.040 15.160 1.360 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 14.720 1.360 15.040 ;
      LAYER met4 ;
        RECT 1.040 14.720 1.360 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 14.280 1.360 14.600 ;
      LAYER met4 ;
        RECT 1.040 14.280 1.360 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 13.840 1.360 14.160 ;
      LAYER met4 ;
        RECT 1.040 13.840 1.360 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 13.400 1.360 13.720 ;
      LAYER met4 ;
        RECT 1.040 13.400 1.360 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.040 12.960 1.360 13.280 ;
      LAYER met4 ;
        RECT 1.040 12.960 1.360 13.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 16.040 0.950 16.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 15.600 0.950 15.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 15.160 0.950 15.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 14.720 0.950 15.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 14.280 0.950 14.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 13.840 0.950 14.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 13.400 0.950 13.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 12.960 0.950 13.280 ;
    END
  END VDDA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
  END VSSD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
  END VSSA
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
  END VSSIO_Q
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  OBS
      LAYER met3 ;
        RECT 0.600 12.940 24.500 16.380 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 94.585 75.000 172.185 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__overlay_vdda_lvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vddio_hvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vddio_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSIO
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
  END VSSIO
  PIN VSSA
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
  END VSSA
  PIN VDDIO
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN VCCHIB
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
  END VCCHIB
  PIN VDDA
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
  END VDDA
  PIN VCCD
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
  END VCCD
  PIN VSSIO_Q
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
  END VSWITCH
  PIN VSSD
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
  END VSSD
  PIN AMUXBUS_A
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.495 19.790 74.290 94.765 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 96.585 75.000 174.185 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__overlay_vddio_hvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vddio_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vddio_lvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 62.090 74.655 66.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 66.260 74.565 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 65.850 74.565 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 65.440 74.565 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 65.030 74.565 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 64.620 74.565 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 64.210 74.565 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 63.800 74.565 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 63.390 74.565 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 62.980 74.565 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 62.570 74.565 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 62.160 74.565 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 66.260 74.155 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 65.850 74.155 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 65.440 74.155 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 65.030 74.155 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 64.620 74.155 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 64.210 74.155 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 63.800 74.155 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 63.390 74.155 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 62.980 74.155 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 62.570 74.155 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 62.160 74.155 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 66.260 73.745 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 65.850 73.745 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 65.440 73.745 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 65.030 73.745 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 64.620 73.745 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 64.210 73.745 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 63.800 73.745 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 63.390 73.745 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 62.980 73.745 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 62.570 73.745 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 62.160 73.745 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 66.260 73.335 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 65.850 73.335 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 65.440 73.335 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 65.030 73.335 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 64.620 73.335 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 64.210 73.335 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 63.800 73.335 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 63.390 73.335 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 62.980 73.335 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 62.570 73.335 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 62.160 73.335 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 66.260 72.925 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 65.850 72.925 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 65.440 72.925 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 65.030 72.925 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 64.620 72.925 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 64.210 72.925 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 63.800 72.925 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 63.390 72.925 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 62.980 72.925 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 62.570 72.925 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 62.160 72.925 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 66.260 72.515 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 65.850 72.515 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 65.440 72.515 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 65.030 72.515 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 64.620 72.515 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 64.210 72.515 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 63.800 72.515 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 63.390 72.515 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 62.980 72.515 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 62.570 72.515 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 62.160 72.515 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 66.260 72.105 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 65.850 72.105 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 65.440 72.105 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 65.030 72.105 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 64.620 72.105 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 64.210 72.105 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 63.800 72.105 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 63.390 72.105 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 62.980 72.105 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 62.570 72.105 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 62.160 72.105 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 66.260 71.700 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 65.850 71.700 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 65.440 71.700 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 65.030 71.700 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 64.620 71.700 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 64.210 71.700 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 63.800 71.700 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 63.390 71.700 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 62.980 71.700 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 62.570 71.700 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 62.160 71.700 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 66.260 71.295 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 65.850 71.295 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 65.440 71.295 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 65.030 71.295 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 64.620 71.295 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 64.210 71.295 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 63.800 71.295 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 63.390 71.295 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 62.980 71.295 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 62.570 71.295 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 62.160 71.295 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 66.260 70.890 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 65.850 70.890 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 65.440 70.890 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 65.030 70.890 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 64.620 70.890 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 64.210 70.890 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 63.800 70.890 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 63.390 70.890 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 62.980 70.890 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 62.570 70.890 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 62.160 70.890 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 66.260 70.485 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 65.850 70.485 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 65.440 70.485 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 65.030 70.485 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 64.620 70.485 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 64.210 70.485 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 63.800 70.485 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 63.390 70.485 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 62.980 70.485 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 62.570 70.485 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 62.160 70.485 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 66.260 70.080 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 65.850 70.080 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 65.440 70.080 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 65.030 70.080 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 64.620 70.080 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 64.210 70.080 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 63.800 70.080 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 63.390 70.080 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 62.980 70.080 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 62.570 70.080 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 62.160 70.080 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 66.260 69.675 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 65.850 69.675 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 65.440 69.675 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 65.030 69.675 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 64.620 69.675 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 64.210 69.675 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 63.800 69.675 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 63.390 69.675 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 62.980 69.675 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 62.570 69.675 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 62.160 69.675 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 66.260 69.270 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 65.850 69.270 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 65.440 69.270 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 65.030 69.270 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 64.620 69.270 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 64.210 69.270 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 63.800 69.270 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 63.390 69.270 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 62.980 69.270 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 62.570 69.270 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 62.160 69.270 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 66.260 68.865 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 65.850 68.865 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 65.440 68.865 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 65.030 68.865 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 64.620 68.865 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 64.210 68.865 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 63.800 68.865 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 63.390 68.865 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 62.980 68.865 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 62.570 68.865 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 62.160 68.865 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 66.260 68.460 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 65.850 68.460 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 65.440 68.460 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 65.030 68.460 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 64.620 68.460 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 64.210 68.460 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 63.800 68.460 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 63.390 68.460 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 62.980 68.460 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 62.570 68.460 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 62.160 68.460 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 66.260 68.055 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 65.850 68.055 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 65.440 68.055 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 65.030 68.055 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 64.620 68.055 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 64.210 68.055 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 63.800 68.055 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 63.390 68.055 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 62.980 68.055 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 62.570 68.055 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 62.160 68.055 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 66.260 67.650 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 65.850 67.650 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 65.440 67.650 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 65.030 67.650 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 64.620 67.650 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 64.210 67.650 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 63.800 67.650 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 63.390 67.650 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 62.980 67.650 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 62.570 67.650 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 62.160 67.650 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 66.260 67.245 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 65.850 67.245 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 65.440 67.245 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 65.030 67.245 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 64.620 67.245 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 64.210 67.245 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 63.800 67.245 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 63.390 67.245 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 62.980 67.245 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 62.570 67.245 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 62.160 67.245 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 66.260 66.840 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 65.850 66.840 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 65.440 66.840 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 65.030 66.840 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 64.620 66.840 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 64.210 66.840 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 63.800 66.840 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 63.390 66.840 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 62.980 66.840 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 62.570 66.840 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 62.160 66.840 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 66.260 66.435 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 65.850 66.435 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 65.440 66.435 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 65.030 66.435 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 64.620 66.435 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 64.210 66.435 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 63.800 66.435 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 63.390 66.435 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 62.980 66.435 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 62.570 66.435 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 62.160 66.435 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 66.260 66.030 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 65.850 66.030 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 65.440 66.030 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 65.030 66.030 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 64.620 66.030 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 64.210 66.030 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 63.800 66.030 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 63.390 66.030 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 62.980 66.030 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 62.570 66.030 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 62.160 66.030 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 66.260 65.625 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 65.850 65.625 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 65.440 65.625 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 65.030 65.625 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 64.620 65.625 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 64.210 65.625 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 63.800 65.625 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 63.390 65.625 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 62.980 65.625 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 62.570 65.625 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 62.160 65.625 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 66.260 65.220 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 65.850 65.220 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 65.440 65.220 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 65.030 65.220 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 64.620 65.220 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 64.210 65.220 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 63.800 65.220 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 63.390 65.220 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 62.980 65.220 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 62.570 65.220 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 62.160 65.220 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 66.260 64.815 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 65.850 64.815 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 65.440 64.815 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 65.030 64.815 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 64.620 64.815 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 64.210 64.815 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 63.800 64.815 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 63.390 64.815 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 62.980 64.815 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 62.570 64.815 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 62.160 64.815 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 66.260 64.410 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 65.850 64.410 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 65.440 64.410 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 65.030 64.410 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 64.620 64.410 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 64.210 64.410 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 63.800 64.410 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 63.390 64.410 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 62.980 64.410 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 62.570 64.410 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 62.160 64.410 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 66.260 64.005 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 65.850 64.005 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 65.440 64.005 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 65.030 64.005 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 64.620 64.005 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 64.210 64.005 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 63.800 64.005 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 63.390 64.005 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 62.980 64.005 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 62.570 64.005 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 62.160 64.005 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 66.260 63.600 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 65.850 63.600 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 65.440 63.600 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 65.030 63.600 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 64.620 63.600 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 64.210 63.600 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 63.800 63.600 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 63.390 63.600 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 62.980 63.600 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 62.570 63.600 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 62.160 63.600 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 66.260 63.195 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 65.850 63.195 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 65.440 63.195 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 65.030 63.195 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 64.620 63.195 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 64.210 63.195 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 63.800 63.195 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 63.390 63.195 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 62.980 63.195 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 62.570 63.195 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 62.160 63.195 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 66.260 62.790 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 65.850 62.790 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 65.440 62.790 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 65.030 62.790 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 64.620 62.790 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 64.210 62.790 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 63.800 62.790 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 63.390 62.790 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 62.980 62.790 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 62.570 62.790 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 62.160 62.790 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 66.260 62.385 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 65.850 62.385 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 65.440 62.385 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 65.030 62.385 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 64.620 62.385 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 64.210 62.385 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 63.800 62.385 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 63.390 62.385 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 62.980 62.385 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 62.570 62.385 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 62.160 62.385 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 66.260 61.980 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 65.850 61.980 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 65.440 61.980 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 65.030 61.980 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 64.620 61.980 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 64.210 61.980 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 63.800 61.980 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 63.390 61.980 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 62.980 61.980 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 62.570 61.980 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 62.160 61.980 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 66.260 61.575 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 65.850 61.575 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 65.440 61.575 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 65.030 61.575 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 64.620 61.575 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 64.210 61.575 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 63.800 61.575 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 63.390 61.575 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 62.980 61.575 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 62.570 61.575 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 62.160 61.575 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 66.260 61.170 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 65.850 61.170 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 65.440 61.170 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 65.030 61.170 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 64.620 61.170 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 64.210 61.170 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 63.800 61.170 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 63.390 61.170 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 62.980 61.170 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 62.570 61.170 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 62.160 61.170 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 66.260 60.765 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 65.850 60.765 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 65.440 60.765 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 65.030 60.765 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 64.620 60.765 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 64.210 60.765 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 63.800 60.765 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 63.390 60.765 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 62.980 60.765 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 62.570 60.765 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 62.160 60.765 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 66.260 60.360 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 65.850 60.360 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 65.440 60.360 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 65.030 60.360 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 64.620 60.360 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 64.210 60.360 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 63.800 60.360 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 63.390 60.360 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 62.980 60.360 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 62.570 60.360 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 62.160 60.360 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 66.260 59.955 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 65.850 59.955 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 65.440 59.955 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 65.030 59.955 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 64.620 59.955 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 64.210 59.955 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 63.800 59.955 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 63.390 59.955 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 62.980 59.955 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 62.570 59.955 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 62.160 59.955 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 66.260 59.550 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 65.850 59.550 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 65.440 59.550 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 65.030 59.550 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 64.620 59.550 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 64.210 59.550 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 63.800 59.550 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 63.390 59.550 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 62.980 59.550 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 62.570 59.550 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 62.160 59.550 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 66.260 59.145 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 65.850 59.145 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 65.440 59.145 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 65.030 59.145 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 64.620 59.145 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 64.210 59.145 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 63.800 59.145 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 63.390 59.145 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 62.980 59.145 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 62.570 59.145 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 62.160 59.145 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 66.260 58.740 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 65.850 58.740 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 65.440 58.740 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 65.030 58.740 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 64.620 58.740 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 64.210 58.740 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 63.800 58.740 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 63.390 58.740 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 62.980 58.740 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 62.570 58.740 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 62.160 58.740 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 66.260 58.335 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 65.850 58.335 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 65.440 58.335 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 65.030 58.335 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 64.620 58.335 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 64.210 58.335 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 63.800 58.335 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 63.390 58.335 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 62.980 58.335 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 62.570 58.335 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 62.160 58.335 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 66.260 57.930 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 65.850 57.930 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 65.440 57.930 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 65.030 57.930 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 64.620 57.930 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 64.210 57.930 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 63.800 57.930 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 63.390 57.930 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 62.980 57.930 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 62.570 57.930 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 62.160 57.930 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 66.260 57.525 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 65.850 57.525 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 65.440 57.525 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 65.030 57.525 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 64.620 57.525 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 64.210 57.525 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 63.800 57.525 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 63.390 57.525 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 62.980 57.525 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 62.570 57.525 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 62.160 57.525 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 66.260 57.120 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 65.850 57.120 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 65.440 57.120 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 65.030 57.120 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 64.620 57.120 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 64.210 57.120 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 63.800 57.120 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 63.390 57.120 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 62.980 57.120 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 62.570 57.120 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 62.160 57.120 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 66.260 56.715 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 65.850 56.715 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 65.440 56.715 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 65.030 56.715 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 64.620 56.715 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 64.210 56.715 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 63.800 56.715 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 63.390 56.715 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 62.980 56.715 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 62.570 56.715 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 62.160 56.715 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 66.260 56.310 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 65.850 56.310 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 65.440 56.310 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 65.030 56.310 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 64.620 56.310 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 64.210 56.310 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 63.800 56.310 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 63.390 56.310 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 62.980 56.310 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 62.570 56.310 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 62.160 56.310 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 66.260 55.905 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 65.850 55.905 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 65.440 55.905 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 65.030 55.905 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 64.620 55.905 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 64.210 55.905 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 63.800 55.905 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 63.390 55.905 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 62.980 55.905 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 62.570 55.905 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 62.160 55.905 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 66.260 55.500 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 65.850 55.500 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 65.440 55.500 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 65.030 55.500 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 64.620 55.500 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 64.210 55.500 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 63.800 55.500 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 63.390 55.500 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 62.980 55.500 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 62.570 55.500 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 62.160 55.500 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 66.260 55.095 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 65.850 55.095 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 65.440 55.095 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 65.030 55.095 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 64.620 55.095 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 64.210 55.095 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 63.800 55.095 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 63.390 55.095 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 62.980 55.095 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 62.570 55.095 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 62.160 55.095 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 66.260 54.690 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 65.850 54.690 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 65.440 54.690 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 65.030 54.690 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 64.620 54.690 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 64.210 54.690 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 63.800 54.690 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 63.390 54.690 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 62.980 54.690 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 62.570 54.690 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 62.160 54.690 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 66.260 54.285 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 65.850 54.285 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 65.440 54.285 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 65.030 54.285 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 64.620 54.285 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 64.210 54.285 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 63.800 54.285 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 63.390 54.285 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 62.980 54.285 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 62.570 54.285 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 62.160 54.285 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 66.260 53.880 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 65.850 53.880 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 65.440 53.880 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 65.030 53.880 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 64.620 53.880 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 64.210 53.880 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 63.800 53.880 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 63.390 53.880 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 62.980 53.880 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 62.570 53.880 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 62.160 53.880 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 66.260 53.475 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 65.850 53.475 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 65.440 53.475 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 65.030 53.475 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 64.620 53.475 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 64.210 53.475 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 63.800 53.475 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 63.390 53.475 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 62.980 53.475 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 62.570 53.475 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 62.160 53.475 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 66.260 53.070 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 65.850 53.070 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 65.440 53.070 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 65.030 53.070 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 64.620 53.070 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 64.210 53.070 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 63.800 53.070 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 63.390 53.070 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 62.980 53.070 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 62.570 53.070 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 62.160 53.070 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 66.260 52.665 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 65.850 52.665 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 65.440 52.665 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 65.030 52.665 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 64.620 52.665 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 64.210 52.665 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 63.800 52.665 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 63.390 52.665 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 62.980 52.665 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 62.570 52.665 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 62.160 52.665 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 66.260 52.260 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 65.850 52.260 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 65.440 52.260 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 65.030 52.260 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 64.620 52.260 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 64.210 52.260 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 63.800 52.260 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 63.390 52.260 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 62.980 52.260 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 62.570 52.260 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 62.160 52.260 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 66.260 51.855 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 65.850 51.855 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 65.440 51.855 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 65.030 51.855 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 64.620 51.855 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 64.210 51.855 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 63.800 51.855 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 63.390 51.855 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 62.980 51.855 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 62.570 51.855 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 62.160 51.855 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 66.260 51.450 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 65.850 51.450 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 65.440 51.450 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 65.030 51.450 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 64.620 51.450 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 64.210 51.450 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 63.800 51.450 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 63.390 51.450 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 62.980 51.450 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 62.570 51.450 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 62.160 51.450 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 66.260 51.045 66.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 65.850 51.045 66.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 65.440 51.045 65.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 65.030 51.045 65.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 64.620 51.045 64.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 64.210 51.045 64.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 63.800 51.045 64.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 63.390 51.045 63.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 62.980 51.045 63.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 62.570 51.045 62.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 62.160 51.045 62.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 66.200 24.470 66.520 ;
      LAYER met4 ;
        RECT 24.150 66.200 24.470 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 65.790 24.470 66.110 ;
      LAYER met4 ;
        RECT 24.150 65.790 24.470 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 65.380 24.470 65.700 ;
      LAYER met4 ;
        RECT 24.150 65.380 24.470 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 64.970 24.470 65.290 ;
      LAYER met4 ;
        RECT 24.150 64.970 24.470 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 64.560 24.470 64.880 ;
      LAYER met4 ;
        RECT 24.150 64.560 24.470 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 64.150 24.470 64.470 ;
      LAYER met4 ;
        RECT 24.150 64.150 24.470 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 63.740 24.470 64.060 ;
      LAYER met4 ;
        RECT 24.150 63.740 24.470 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 63.330 24.470 63.650 ;
      LAYER met4 ;
        RECT 24.150 63.330 24.470 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 62.920 24.470 63.240 ;
      LAYER met4 ;
        RECT 24.150 62.920 24.470 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 62.510 24.470 62.830 ;
      LAYER met4 ;
        RECT 24.150 62.510 24.470 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 62.100 24.470 62.420 ;
      LAYER met4 ;
        RECT 24.150 62.100 24.470 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 66.200 24.060 66.520 ;
      LAYER met4 ;
        RECT 23.740 66.200 24.060 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 65.790 24.060 66.110 ;
      LAYER met4 ;
        RECT 23.740 65.790 24.060 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 65.380 24.060 65.700 ;
      LAYER met4 ;
        RECT 23.740 65.380 24.060 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 64.970 24.060 65.290 ;
      LAYER met4 ;
        RECT 23.740 64.970 24.060 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 64.560 24.060 64.880 ;
      LAYER met4 ;
        RECT 23.740 64.560 24.060 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 64.150 24.060 64.470 ;
      LAYER met4 ;
        RECT 23.740 64.150 24.060 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 63.740 24.060 64.060 ;
      LAYER met4 ;
        RECT 23.740 63.740 24.060 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 63.330 24.060 63.650 ;
      LAYER met4 ;
        RECT 23.740 63.330 24.060 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 62.920 24.060 63.240 ;
      LAYER met4 ;
        RECT 23.740 62.920 24.060 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 62.510 24.060 62.830 ;
      LAYER met4 ;
        RECT 23.740 62.510 24.060 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.740 62.100 24.060 62.420 ;
      LAYER met4 ;
        RECT 23.740 62.100 24.060 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 66.200 23.650 66.520 ;
      LAYER met4 ;
        RECT 23.330 66.200 23.650 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 65.790 23.650 66.110 ;
      LAYER met4 ;
        RECT 23.330 65.790 23.650 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 65.380 23.650 65.700 ;
      LAYER met4 ;
        RECT 23.330 65.380 23.650 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 64.970 23.650 65.290 ;
      LAYER met4 ;
        RECT 23.330 64.970 23.650 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 64.560 23.650 64.880 ;
      LAYER met4 ;
        RECT 23.330 64.560 23.650 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 64.150 23.650 64.470 ;
      LAYER met4 ;
        RECT 23.330 64.150 23.650 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 63.740 23.650 64.060 ;
      LAYER met4 ;
        RECT 23.330 63.740 23.650 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 63.330 23.650 63.650 ;
      LAYER met4 ;
        RECT 23.330 63.330 23.650 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 62.920 23.650 63.240 ;
      LAYER met4 ;
        RECT 23.330 62.920 23.650 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 62.510 23.650 62.830 ;
      LAYER met4 ;
        RECT 23.330 62.510 23.650 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.330 62.100 23.650 62.420 ;
      LAYER met4 ;
        RECT 23.330 62.100 23.650 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 66.200 23.240 66.520 ;
      LAYER met4 ;
        RECT 22.920 66.200 23.240 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 65.790 23.240 66.110 ;
      LAYER met4 ;
        RECT 22.920 65.790 23.240 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 65.380 23.240 65.700 ;
      LAYER met4 ;
        RECT 22.920 65.380 23.240 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 64.970 23.240 65.290 ;
      LAYER met4 ;
        RECT 22.920 64.970 23.240 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 64.560 23.240 64.880 ;
      LAYER met4 ;
        RECT 22.920 64.560 23.240 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 64.150 23.240 64.470 ;
      LAYER met4 ;
        RECT 22.920 64.150 23.240 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 63.740 23.240 64.060 ;
      LAYER met4 ;
        RECT 22.920 63.740 23.240 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 63.330 23.240 63.650 ;
      LAYER met4 ;
        RECT 22.920 63.330 23.240 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 62.920 23.240 63.240 ;
      LAYER met4 ;
        RECT 22.920 62.920 23.240 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 62.510 23.240 62.830 ;
      LAYER met4 ;
        RECT 22.920 62.510 23.240 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.920 62.100 23.240 62.420 ;
      LAYER met4 ;
        RECT 22.920 62.100 23.240 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 66.200 22.830 66.520 ;
      LAYER met4 ;
        RECT 22.510 66.200 22.830 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 65.790 22.830 66.110 ;
      LAYER met4 ;
        RECT 22.510 65.790 22.830 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 65.380 22.830 65.700 ;
      LAYER met4 ;
        RECT 22.510 65.380 22.830 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 64.970 22.830 65.290 ;
      LAYER met4 ;
        RECT 22.510 64.970 22.830 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 64.560 22.830 64.880 ;
      LAYER met4 ;
        RECT 22.510 64.560 22.830 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 64.150 22.830 64.470 ;
      LAYER met4 ;
        RECT 22.510 64.150 22.830 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 63.740 22.830 64.060 ;
      LAYER met4 ;
        RECT 22.510 63.740 22.830 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 63.330 22.830 63.650 ;
      LAYER met4 ;
        RECT 22.510 63.330 22.830 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 62.920 22.830 63.240 ;
      LAYER met4 ;
        RECT 22.510 62.920 22.830 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 62.510 22.830 62.830 ;
      LAYER met4 ;
        RECT 22.510 62.510 22.830 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.510 62.100 22.830 62.420 ;
      LAYER met4 ;
        RECT 22.510 62.100 22.830 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 66.200 22.420 66.520 ;
      LAYER met4 ;
        RECT 22.100 66.200 22.420 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 65.790 22.420 66.110 ;
      LAYER met4 ;
        RECT 22.100 65.790 22.420 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 65.380 22.420 65.700 ;
      LAYER met4 ;
        RECT 22.100 65.380 22.420 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 64.970 22.420 65.290 ;
      LAYER met4 ;
        RECT 22.100 64.970 22.420 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 64.560 22.420 64.880 ;
      LAYER met4 ;
        RECT 22.100 64.560 22.420 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 64.150 22.420 64.470 ;
      LAYER met4 ;
        RECT 22.100 64.150 22.420 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 63.740 22.420 64.060 ;
      LAYER met4 ;
        RECT 22.100 63.740 22.420 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 63.330 22.420 63.650 ;
      LAYER met4 ;
        RECT 22.100 63.330 22.420 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 62.920 22.420 63.240 ;
      LAYER met4 ;
        RECT 22.100 62.920 22.420 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 62.510 22.420 62.830 ;
      LAYER met4 ;
        RECT 22.100 62.510 22.420 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.100 62.100 22.420 62.420 ;
      LAYER met4 ;
        RECT 22.100 62.100 22.420 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 66.200 22.010 66.520 ;
      LAYER met4 ;
        RECT 21.690 66.200 22.010 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 65.790 22.010 66.110 ;
      LAYER met4 ;
        RECT 21.690 65.790 22.010 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 65.380 22.010 65.700 ;
      LAYER met4 ;
        RECT 21.690 65.380 22.010 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 64.970 22.010 65.290 ;
      LAYER met4 ;
        RECT 21.690 64.970 22.010 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 64.560 22.010 64.880 ;
      LAYER met4 ;
        RECT 21.690 64.560 22.010 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 64.150 22.010 64.470 ;
      LAYER met4 ;
        RECT 21.690 64.150 22.010 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 63.740 22.010 64.060 ;
      LAYER met4 ;
        RECT 21.690 63.740 22.010 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 63.330 22.010 63.650 ;
      LAYER met4 ;
        RECT 21.690 63.330 22.010 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 62.920 22.010 63.240 ;
      LAYER met4 ;
        RECT 21.690 62.920 22.010 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 62.510 22.010 62.830 ;
      LAYER met4 ;
        RECT 21.690 62.510 22.010 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.690 62.100 22.010 62.420 ;
      LAYER met4 ;
        RECT 21.690 62.100 22.010 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 66.200 21.605 66.520 ;
      LAYER met4 ;
        RECT 21.285 66.200 21.605 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 65.790 21.605 66.110 ;
      LAYER met4 ;
        RECT 21.285 65.790 21.605 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 65.380 21.605 65.700 ;
      LAYER met4 ;
        RECT 21.285 65.380 21.605 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 64.970 21.605 65.290 ;
      LAYER met4 ;
        RECT 21.285 64.970 21.605 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 64.560 21.605 64.880 ;
      LAYER met4 ;
        RECT 21.285 64.560 21.605 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 64.150 21.605 64.470 ;
      LAYER met4 ;
        RECT 21.285 64.150 21.605 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 63.740 21.605 64.060 ;
      LAYER met4 ;
        RECT 21.285 63.740 21.605 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 63.330 21.605 63.650 ;
      LAYER met4 ;
        RECT 21.285 63.330 21.605 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 62.920 21.605 63.240 ;
      LAYER met4 ;
        RECT 21.285 62.920 21.605 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 62.510 21.605 62.830 ;
      LAYER met4 ;
        RECT 21.285 62.510 21.605 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.285 62.100 21.605 62.420 ;
      LAYER met4 ;
        RECT 21.285 62.100 21.605 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 66.200 21.200 66.520 ;
      LAYER met4 ;
        RECT 20.880 66.200 21.200 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 65.790 21.200 66.110 ;
      LAYER met4 ;
        RECT 20.880 65.790 21.200 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 65.380 21.200 65.700 ;
      LAYER met4 ;
        RECT 20.880 65.380 21.200 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 64.970 21.200 65.290 ;
      LAYER met4 ;
        RECT 20.880 64.970 21.200 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 64.560 21.200 64.880 ;
      LAYER met4 ;
        RECT 20.880 64.560 21.200 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 64.150 21.200 64.470 ;
      LAYER met4 ;
        RECT 20.880 64.150 21.200 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 63.740 21.200 64.060 ;
      LAYER met4 ;
        RECT 20.880 63.740 21.200 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 63.330 21.200 63.650 ;
      LAYER met4 ;
        RECT 20.880 63.330 21.200 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 62.920 21.200 63.240 ;
      LAYER met4 ;
        RECT 20.880 62.920 21.200 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 62.510 21.200 62.830 ;
      LAYER met4 ;
        RECT 20.880 62.510 21.200 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.880 62.100 21.200 62.420 ;
      LAYER met4 ;
        RECT 20.880 62.100 21.200 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 66.200 20.795 66.520 ;
      LAYER met4 ;
        RECT 20.475 66.200 20.795 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 65.790 20.795 66.110 ;
      LAYER met4 ;
        RECT 20.475 65.790 20.795 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 65.380 20.795 65.700 ;
      LAYER met4 ;
        RECT 20.475 65.380 20.795 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 64.970 20.795 65.290 ;
      LAYER met4 ;
        RECT 20.475 64.970 20.795 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 64.560 20.795 64.880 ;
      LAYER met4 ;
        RECT 20.475 64.560 20.795 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 64.150 20.795 64.470 ;
      LAYER met4 ;
        RECT 20.475 64.150 20.795 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 63.740 20.795 64.060 ;
      LAYER met4 ;
        RECT 20.475 63.740 20.795 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 63.330 20.795 63.650 ;
      LAYER met4 ;
        RECT 20.475 63.330 20.795 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 62.920 20.795 63.240 ;
      LAYER met4 ;
        RECT 20.475 62.920 20.795 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 62.510 20.795 62.830 ;
      LAYER met4 ;
        RECT 20.475 62.510 20.795 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.475 62.100 20.795 62.420 ;
      LAYER met4 ;
        RECT 20.475 62.100 20.795 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 66.200 20.390 66.520 ;
      LAYER met4 ;
        RECT 20.070 66.200 20.390 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 65.790 20.390 66.110 ;
      LAYER met4 ;
        RECT 20.070 65.790 20.390 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 65.380 20.390 65.700 ;
      LAYER met4 ;
        RECT 20.070 65.380 20.390 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 64.970 20.390 65.290 ;
      LAYER met4 ;
        RECT 20.070 64.970 20.390 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 64.560 20.390 64.880 ;
      LAYER met4 ;
        RECT 20.070 64.560 20.390 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 64.150 20.390 64.470 ;
      LAYER met4 ;
        RECT 20.070 64.150 20.390 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 63.740 20.390 64.060 ;
      LAYER met4 ;
        RECT 20.070 63.740 20.390 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 63.330 20.390 63.650 ;
      LAYER met4 ;
        RECT 20.070 63.330 20.390 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 62.920 20.390 63.240 ;
      LAYER met4 ;
        RECT 20.070 62.920 20.390 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 62.510 20.390 62.830 ;
      LAYER met4 ;
        RECT 20.070 62.510 20.390 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.070 62.100 20.390 62.420 ;
      LAYER met4 ;
        RECT 20.070 62.100 20.390 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 66.200 19.985 66.520 ;
      LAYER met4 ;
        RECT 19.665 66.200 19.985 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 65.790 19.985 66.110 ;
      LAYER met4 ;
        RECT 19.665 65.790 19.985 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 65.380 19.985 65.700 ;
      LAYER met4 ;
        RECT 19.665 65.380 19.985 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 64.970 19.985 65.290 ;
      LAYER met4 ;
        RECT 19.665 64.970 19.985 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 64.560 19.985 64.880 ;
      LAYER met4 ;
        RECT 19.665 64.560 19.985 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 64.150 19.985 64.470 ;
      LAYER met4 ;
        RECT 19.665 64.150 19.985 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 63.740 19.985 64.060 ;
      LAYER met4 ;
        RECT 19.665 63.740 19.985 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 63.330 19.985 63.650 ;
      LAYER met4 ;
        RECT 19.665 63.330 19.985 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 62.920 19.985 63.240 ;
      LAYER met4 ;
        RECT 19.665 62.920 19.985 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 62.510 19.985 62.830 ;
      LAYER met4 ;
        RECT 19.665 62.510 19.985 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.665 62.100 19.985 62.420 ;
      LAYER met4 ;
        RECT 19.665 62.100 19.985 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 66.200 19.580 66.520 ;
      LAYER met4 ;
        RECT 19.260 66.200 19.580 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 65.790 19.580 66.110 ;
      LAYER met4 ;
        RECT 19.260 65.790 19.580 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 65.380 19.580 65.700 ;
      LAYER met4 ;
        RECT 19.260 65.380 19.580 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 64.970 19.580 65.290 ;
      LAYER met4 ;
        RECT 19.260 64.970 19.580 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 64.560 19.580 64.880 ;
      LAYER met4 ;
        RECT 19.260 64.560 19.580 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 64.150 19.580 64.470 ;
      LAYER met4 ;
        RECT 19.260 64.150 19.580 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 63.740 19.580 64.060 ;
      LAYER met4 ;
        RECT 19.260 63.740 19.580 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 63.330 19.580 63.650 ;
      LAYER met4 ;
        RECT 19.260 63.330 19.580 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 62.920 19.580 63.240 ;
      LAYER met4 ;
        RECT 19.260 62.920 19.580 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 62.510 19.580 62.830 ;
      LAYER met4 ;
        RECT 19.260 62.510 19.580 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.260 62.100 19.580 62.420 ;
      LAYER met4 ;
        RECT 19.260 62.100 19.580 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 66.200 19.175 66.520 ;
      LAYER met4 ;
        RECT 18.855 66.200 19.175 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 65.790 19.175 66.110 ;
      LAYER met4 ;
        RECT 18.855 65.790 19.175 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 65.380 19.175 65.700 ;
      LAYER met4 ;
        RECT 18.855 65.380 19.175 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 64.970 19.175 65.290 ;
      LAYER met4 ;
        RECT 18.855 64.970 19.175 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 64.560 19.175 64.880 ;
      LAYER met4 ;
        RECT 18.855 64.560 19.175 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 64.150 19.175 64.470 ;
      LAYER met4 ;
        RECT 18.855 64.150 19.175 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 63.740 19.175 64.060 ;
      LAYER met4 ;
        RECT 18.855 63.740 19.175 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 63.330 19.175 63.650 ;
      LAYER met4 ;
        RECT 18.855 63.330 19.175 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 62.920 19.175 63.240 ;
      LAYER met4 ;
        RECT 18.855 62.920 19.175 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 62.510 19.175 62.830 ;
      LAYER met4 ;
        RECT 18.855 62.510 19.175 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.855 62.100 19.175 62.420 ;
      LAYER met4 ;
        RECT 18.855 62.100 19.175 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 66.200 18.770 66.520 ;
      LAYER met4 ;
        RECT 18.450 66.200 18.770 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 65.790 18.770 66.110 ;
      LAYER met4 ;
        RECT 18.450 65.790 18.770 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 65.380 18.770 65.700 ;
      LAYER met4 ;
        RECT 18.450 65.380 18.770 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 64.970 18.770 65.290 ;
      LAYER met4 ;
        RECT 18.450 64.970 18.770 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 64.560 18.770 64.880 ;
      LAYER met4 ;
        RECT 18.450 64.560 18.770 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 64.150 18.770 64.470 ;
      LAYER met4 ;
        RECT 18.450 64.150 18.770 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 63.740 18.770 64.060 ;
      LAYER met4 ;
        RECT 18.450 63.740 18.770 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 63.330 18.770 63.650 ;
      LAYER met4 ;
        RECT 18.450 63.330 18.770 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 62.920 18.770 63.240 ;
      LAYER met4 ;
        RECT 18.450 62.920 18.770 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 62.510 18.770 62.830 ;
      LAYER met4 ;
        RECT 18.450 62.510 18.770 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.450 62.100 18.770 62.420 ;
      LAYER met4 ;
        RECT 18.450 62.100 18.770 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 66.200 18.365 66.520 ;
      LAYER met4 ;
        RECT 18.045 66.200 18.365 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 65.790 18.365 66.110 ;
      LAYER met4 ;
        RECT 18.045 65.790 18.365 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 65.380 18.365 65.700 ;
      LAYER met4 ;
        RECT 18.045 65.380 18.365 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 64.970 18.365 65.290 ;
      LAYER met4 ;
        RECT 18.045 64.970 18.365 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 64.560 18.365 64.880 ;
      LAYER met4 ;
        RECT 18.045 64.560 18.365 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 64.150 18.365 64.470 ;
      LAYER met4 ;
        RECT 18.045 64.150 18.365 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 63.740 18.365 64.060 ;
      LAYER met4 ;
        RECT 18.045 63.740 18.365 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 63.330 18.365 63.650 ;
      LAYER met4 ;
        RECT 18.045 63.330 18.365 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 62.920 18.365 63.240 ;
      LAYER met4 ;
        RECT 18.045 62.920 18.365 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 62.510 18.365 62.830 ;
      LAYER met4 ;
        RECT 18.045 62.510 18.365 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 62.100 18.365 62.420 ;
      LAYER met4 ;
        RECT 18.045 62.100 18.365 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 66.200 17.960 66.520 ;
      LAYER met4 ;
        RECT 17.640 66.200 17.960 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 65.790 17.960 66.110 ;
      LAYER met4 ;
        RECT 17.640 65.790 17.960 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 65.380 17.960 65.700 ;
      LAYER met4 ;
        RECT 17.640 65.380 17.960 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 64.970 17.960 65.290 ;
      LAYER met4 ;
        RECT 17.640 64.970 17.960 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 64.560 17.960 64.880 ;
      LAYER met4 ;
        RECT 17.640 64.560 17.960 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 64.150 17.960 64.470 ;
      LAYER met4 ;
        RECT 17.640 64.150 17.960 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 63.740 17.960 64.060 ;
      LAYER met4 ;
        RECT 17.640 63.740 17.960 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 63.330 17.960 63.650 ;
      LAYER met4 ;
        RECT 17.640 63.330 17.960 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 62.920 17.960 63.240 ;
      LAYER met4 ;
        RECT 17.640 62.920 17.960 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 62.510 17.960 62.830 ;
      LAYER met4 ;
        RECT 17.640 62.510 17.960 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.640 62.100 17.960 62.420 ;
      LAYER met4 ;
        RECT 17.640 62.100 17.960 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 66.200 17.555 66.520 ;
      LAYER met4 ;
        RECT 17.235 66.200 17.555 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 65.790 17.555 66.110 ;
      LAYER met4 ;
        RECT 17.235 65.790 17.555 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 65.380 17.555 65.700 ;
      LAYER met4 ;
        RECT 17.235 65.380 17.555 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 64.970 17.555 65.290 ;
      LAYER met4 ;
        RECT 17.235 64.970 17.555 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 64.560 17.555 64.880 ;
      LAYER met4 ;
        RECT 17.235 64.560 17.555 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 64.150 17.555 64.470 ;
      LAYER met4 ;
        RECT 17.235 64.150 17.555 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 63.740 17.555 64.060 ;
      LAYER met4 ;
        RECT 17.235 63.740 17.555 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 63.330 17.555 63.650 ;
      LAYER met4 ;
        RECT 17.235 63.330 17.555 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 62.920 17.555 63.240 ;
      LAYER met4 ;
        RECT 17.235 62.920 17.555 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 62.510 17.555 62.830 ;
      LAYER met4 ;
        RECT 17.235 62.510 17.555 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.235 62.100 17.555 62.420 ;
      LAYER met4 ;
        RECT 17.235 62.100 17.555 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 66.200 17.150 66.520 ;
      LAYER met4 ;
        RECT 16.830 66.200 17.150 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 65.790 17.150 66.110 ;
      LAYER met4 ;
        RECT 16.830 65.790 17.150 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 65.380 17.150 65.700 ;
      LAYER met4 ;
        RECT 16.830 65.380 17.150 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 64.970 17.150 65.290 ;
      LAYER met4 ;
        RECT 16.830 64.970 17.150 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 64.560 17.150 64.880 ;
      LAYER met4 ;
        RECT 16.830 64.560 17.150 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 64.150 17.150 64.470 ;
      LAYER met4 ;
        RECT 16.830 64.150 17.150 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 63.740 17.150 64.060 ;
      LAYER met4 ;
        RECT 16.830 63.740 17.150 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 63.330 17.150 63.650 ;
      LAYER met4 ;
        RECT 16.830 63.330 17.150 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 62.920 17.150 63.240 ;
      LAYER met4 ;
        RECT 16.830 62.920 17.150 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 62.510 17.150 62.830 ;
      LAYER met4 ;
        RECT 16.830 62.510 17.150 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.830 62.100 17.150 62.420 ;
      LAYER met4 ;
        RECT 16.830 62.100 17.150 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 66.200 16.745 66.520 ;
      LAYER met4 ;
        RECT 16.425 66.200 16.745 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 65.790 16.745 66.110 ;
      LAYER met4 ;
        RECT 16.425 65.790 16.745 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 65.380 16.745 65.700 ;
      LAYER met4 ;
        RECT 16.425 65.380 16.745 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 64.970 16.745 65.290 ;
      LAYER met4 ;
        RECT 16.425 64.970 16.745 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 64.560 16.745 64.880 ;
      LAYER met4 ;
        RECT 16.425 64.560 16.745 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 64.150 16.745 64.470 ;
      LAYER met4 ;
        RECT 16.425 64.150 16.745 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 63.740 16.745 64.060 ;
      LAYER met4 ;
        RECT 16.425 63.740 16.745 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 63.330 16.745 63.650 ;
      LAYER met4 ;
        RECT 16.425 63.330 16.745 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 62.920 16.745 63.240 ;
      LAYER met4 ;
        RECT 16.425 62.920 16.745 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 62.510 16.745 62.830 ;
      LAYER met4 ;
        RECT 16.425 62.510 16.745 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.425 62.100 16.745 62.420 ;
      LAYER met4 ;
        RECT 16.425 62.100 16.745 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 66.200 16.340 66.520 ;
      LAYER met4 ;
        RECT 16.020 66.200 16.340 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 65.790 16.340 66.110 ;
      LAYER met4 ;
        RECT 16.020 65.790 16.340 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 65.380 16.340 65.700 ;
      LAYER met4 ;
        RECT 16.020 65.380 16.340 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 64.970 16.340 65.290 ;
      LAYER met4 ;
        RECT 16.020 64.970 16.340 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 64.560 16.340 64.880 ;
      LAYER met4 ;
        RECT 16.020 64.560 16.340 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 64.150 16.340 64.470 ;
      LAYER met4 ;
        RECT 16.020 64.150 16.340 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 63.740 16.340 64.060 ;
      LAYER met4 ;
        RECT 16.020 63.740 16.340 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 63.330 16.340 63.650 ;
      LAYER met4 ;
        RECT 16.020 63.330 16.340 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 62.920 16.340 63.240 ;
      LAYER met4 ;
        RECT 16.020 62.920 16.340 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 62.510 16.340 62.830 ;
      LAYER met4 ;
        RECT 16.020 62.510 16.340 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.020 62.100 16.340 62.420 ;
      LAYER met4 ;
        RECT 16.020 62.100 16.340 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 66.200 15.935 66.520 ;
      LAYER met4 ;
        RECT 15.615 66.200 15.935 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 65.790 15.935 66.110 ;
      LAYER met4 ;
        RECT 15.615 65.790 15.935 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 65.380 15.935 65.700 ;
      LAYER met4 ;
        RECT 15.615 65.380 15.935 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 64.970 15.935 65.290 ;
      LAYER met4 ;
        RECT 15.615 64.970 15.935 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 64.560 15.935 64.880 ;
      LAYER met4 ;
        RECT 15.615 64.560 15.935 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 64.150 15.935 64.470 ;
      LAYER met4 ;
        RECT 15.615 64.150 15.935 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 63.740 15.935 64.060 ;
      LAYER met4 ;
        RECT 15.615 63.740 15.935 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 63.330 15.935 63.650 ;
      LAYER met4 ;
        RECT 15.615 63.330 15.935 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 62.920 15.935 63.240 ;
      LAYER met4 ;
        RECT 15.615 62.920 15.935 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 62.510 15.935 62.830 ;
      LAYER met4 ;
        RECT 15.615 62.510 15.935 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.615 62.100 15.935 62.420 ;
      LAYER met4 ;
        RECT 15.615 62.100 15.935 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 66.200 15.530 66.520 ;
      LAYER met4 ;
        RECT 15.210 66.200 15.530 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 65.790 15.530 66.110 ;
      LAYER met4 ;
        RECT 15.210 65.790 15.530 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 65.380 15.530 65.700 ;
      LAYER met4 ;
        RECT 15.210 65.380 15.530 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 64.970 15.530 65.290 ;
      LAYER met4 ;
        RECT 15.210 64.970 15.530 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 64.560 15.530 64.880 ;
      LAYER met4 ;
        RECT 15.210 64.560 15.530 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 64.150 15.530 64.470 ;
      LAYER met4 ;
        RECT 15.210 64.150 15.530 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 63.740 15.530 64.060 ;
      LAYER met4 ;
        RECT 15.210 63.740 15.530 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 63.330 15.530 63.650 ;
      LAYER met4 ;
        RECT 15.210 63.330 15.530 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 62.920 15.530 63.240 ;
      LAYER met4 ;
        RECT 15.210 62.920 15.530 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 62.510 15.530 62.830 ;
      LAYER met4 ;
        RECT 15.210 62.510 15.530 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.210 62.100 15.530 62.420 ;
      LAYER met4 ;
        RECT 15.210 62.100 15.530 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 66.200 15.125 66.520 ;
      LAYER met4 ;
        RECT 14.805 66.200 15.125 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 65.790 15.125 66.110 ;
      LAYER met4 ;
        RECT 14.805 65.790 15.125 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 65.380 15.125 65.700 ;
      LAYER met4 ;
        RECT 14.805 65.380 15.125 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 64.970 15.125 65.290 ;
      LAYER met4 ;
        RECT 14.805 64.970 15.125 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 64.560 15.125 64.880 ;
      LAYER met4 ;
        RECT 14.805 64.560 15.125 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 64.150 15.125 64.470 ;
      LAYER met4 ;
        RECT 14.805 64.150 15.125 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 63.740 15.125 64.060 ;
      LAYER met4 ;
        RECT 14.805 63.740 15.125 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 63.330 15.125 63.650 ;
      LAYER met4 ;
        RECT 14.805 63.330 15.125 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 62.920 15.125 63.240 ;
      LAYER met4 ;
        RECT 14.805 62.920 15.125 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 62.510 15.125 62.830 ;
      LAYER met4 ;
        RECT 14.805 62.510 15.125 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.805 62.100 15.125 62.420 ;
      LAYER met4 ;
        RECT 14.805 62.100 15.125 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 66.200 14.720 66.520 ;
      LAYER met4 ;
        RECT 14.400 66.200 14.720 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 65.790 14.720 66.110 ;
      LAYER met4 ;
        RECT 14.400 65.790 14.720 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 65.380 14.720 65.700 ;
      LAYER met4 ;
        RECT 14.400 65.380 14.720 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 64.970 14.720 65.290 ;
      LAYER met4 ;
        RECT 14.400 64.970 14.720 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 64.560 14.720 64.880 ;
      LAYER met4 ;
        RECT 14.400 64.560 14.720 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 64.150 14.720 64.470 ;
      LAYER met4 ;
        RECT 14.400 64.150 14.720 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 63.740 14.720 64.060 ;
      LAYER met4 ;
        RECT 14.400 63.740 14.720 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 63.330 14.720 63.650 ;
      LAYER met4 ;
        RECT 14.400 63.330 14.720 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 62.920 14.720 63.240 ;
      LAYER met4 ;
        RECT 14.400 62.920 14.720 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 62.510 14.720 62.830 ;
      LAYER met4 ;
        RECT 14.400 62.510 14.720 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.400 62.100 14.720 62.420 ;
      LAYER met4 ;
        RECT 14.400 62.100 14.720 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 66.200 14.315 66.520 ;
      LAYER met4 ;
        RECT 13.995 66.200 14.315 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 65.790 14.315 66.110 ;
      LAYER met4 ;
        RECT 13.995 65.790 14.315 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 65.380 14.315 65.700 ;
      LAYER met4 ;
        RECT 13.995 65.380 14.315 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 64.970 14.315 65.290 ;
      LAYER met4 ;
        RECT 13.995 64.970 14.315 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 64.560 14.315 64.880 ;
      LAYER met4 ;
        RECT 13.995 64.560 14.315 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 64.150 14.315 64.470 ;
      LAYER met4 ;
        RECT 13.995 64.150 14.315 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 63.740 14.315 64.060 ;
      LAYER met4 ;
        RECT 13.995 63.740 14.315 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 63.330 14.315 63.650 ;
      LAYER met4 ;
        RECT 13.995 63.330 14.315 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 62.920 14.315 63.240 ;
      LAYER met4 ;
        RECT 13.995 62.920 14.315 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 62.510 14.315 62.830 ;
      LAYER met4 ;
        RECT 13.995 62.510 14.315 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.995 62.100 14.315 62.420 ;
      LAYER met4 ;
        RECT 13.995 62.100 14.315 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 66.200 13.910 66.520 ;
      LAYER met4 ;
        RECT 13.590 66.200 13.910 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 65.790 13.910 66.110 ;
      LAYER met4 ;
        RECT 13.590 65.790 13.910 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 65.380 13.910 65.700 ;
      LAYER met4 ;
        RECT 13.590 65.380 13.910 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 64.970 13.910 65.290 ;
      LAYER met4 ;
        RECT 13.590 64.970 13.910 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 64.560 13.910 64.880 ;
      LAYER met4 ;
        RECT 13.590 64.560 13.910 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 64.150 13.910 64.470 ;
      LAYER met4 ;
        RECT 13.590 64.150 13.910 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 63.740 13.910 64.060 ;
      LAYER met4 ;
        RECT 13.590 63.740 13.910 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 63.330 13.910 63.650 ;
      LAYER met4 ;
        RECT 13.590 63.330 13.910 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 62.920 13.910 63.240 ;
      LAYER met4 ;
        RECT 13.590 62.920 13.910 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 62.510 13.910 62.830 ;
      LAYER met4 ;
        RECT 13.590 62.510 13.910 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.590 62.100 13.910 62.420 ;
      LAYER met4 ;
        RECT 13.590 62.100 13.910 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 66.200 13.505 66.520 ;
      LAYER met4 ;
        RECT 13.185 66.200 13.505 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 65.790 13.505 66.110 ;
      LAYER met4 ;
        RECT 13.185 65.790 13.505 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 65.380 13.505 65.700 ;
      LAYER met4 ;
        RECT 13.185 65.380 13.505 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 64.970 13.505 65.290 ;
      LAYER met4 ;
        RECT 13.185 64.970 13.505 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 64.560 13.505 64.880 ;
      LAYER met4 ;
        RECT 13.185 64.560 13.505 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 64.150 13.505 64.470 ;
      LAYER met4 ;
        RECT 13.185 64.150 13.505 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 63.740 13.505 64.060 ;
      LAYER met4 ;
        RECT 13.185 63.740 13.505 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 63.330 13.505 63.650 ;
      LAYER met4 ;
        RECT 13.185 63.330 13.505 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 62.920 13.505 63.240 ;
      LAYER met4 ;
        RECT 13.185 62.920 13.505 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 62.510 13.505 62.830 ;
      LAYER met4 ;
        RECT 13.185 62.510 13.505 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 62.100 13.505 62.420 ;
      LAYER met4 ;
        RECT 13.185 62.100 13.505 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 66.200 13.100 66.520 ;
      LAYER met4 ;
        RECT 12.780 66.200 13.100 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 65.790 13.100 66.110 ;
      LAYER met4 ;
        RECT 12.780 65.790 13.100 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 65.380 13.100 65.700 ;
      LAYER met4 ;
        RECT 12.780 65.380 13.100 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 64.970 13.100 65.290 ;
      LAYER met4 ;
        RECT 12.780 64.970 13.100 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 64.560 13.100 64.880 ;
      LAYER met4 ;
        RECT 12.780 64.560 13.100 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 64.150 13.100 64.470 ;
      LAYER met4 ;
        RECT 12.780 64.150 13.100 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 63.740 13.100 64.060 ;
      LAYER met4 ;
        RECT 12.780 63.740 13.100 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 63.330 13.100 63.650 ;
      LAYER met4 ;
        RECT 12.780 63.330 13.100 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 62.920 13.100 63.240 ;
      LAYER met4 ;
        RECT 12.780 62.920 13.100 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 62.510 13.100 62.830 ;
      LAYER met4 ;
        RECT 12.780 62.510 13.100 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.780 62.100 13.100 62.420 ;
      LAYER met4 ;
        RECT 12.780 62.100 13.100 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 66.200 12.695 66.520 ;
      LAYER met4 ;
        RECT 12.375 66.200 12.695 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 65.790 12.695 66.110 ;
      LAYER met4 ;
        RECT 12.375 65.790 12.695 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 65.380 12.695 65.700 ;
      LAYER met4 ;
        RECT 12.375 65.380 12.695 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 64.970 12.695 65.290 ;
      LAYER met4 ;
        RECT 12.375 64.970 12.695 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 64.560 12.695 64.880 ;
      LAYER met4 ;
        RECT 12.375 64.560 12.695 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 64.150 12.695 64.470 ;
      LAYER met4 ;
        RECT 12.375 64.150 12.695 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 63.740 12.695 64.060 ;
      LAYER met4 ;
        RECT 12.375 63.740 12.695 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 63.330 12.695 63.650 ;
      LAYER met4 ;
        RECT 12.375 63.330 12.695 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 62.920 12.695 63.240 ;
      LAYER met4 ;
        RECT 12.375 62.920 12.695 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 62.510 12.695 62.830 ;
      LAYER met4 ;
        RECT 12.375 62.510 12.695 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.375 62.100 12.695 62.420 ;
      LAYER met4 ;
        RECT 12.375 62.100 12.695 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 66.200 12.290 66.520 ;
      LAYER met4 ;
        RECT 11.970 66.200 12.290 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 65.790 12.290 66.110 ;
      LAYER met4 ;
        RECT 11.970 65.790 12.290 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 65.380 12.290 65.700 ;
      LAYER met4 ;
        RECT 11.970 65.380 12.290 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 64.970 12.290 65.290 ;
      LAYER met4 ;
        RECT 11.970 64.970 12.290 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 64.560 12.290 64.880 ;
      LAYER met4 ;
        RECT 11.970 64.560 12.290 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 64.150 12.290 64.470 ;
      LAYER met4 ;
        RECT 11.970 64.150 12.290 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 63.740 12.290 64.060 ;
      LAYER met4 ;
        RECT 11.970 63.740 12.290 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 63.330 12.290 63.650 ;
      LAYER met4 ;
        RECT 11.970 63.330 12.290 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 62.920 12.290 63.240 ;
      LAYER met4 ;
        RECT 11.970 62.920 12.290 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 62.510 12.290 62.830 ;
      LAYER met4 ;
        RECT 11.970 62.510 12.290 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.970 62.100 12.290 62.420 ;
      LAYER met4 ;
        RECT 11.970 62.100 12.290 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 66.200 11.885 66.520 ;
      LAYER met4 ;
        RECT 11.565 66.200 11.885 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 65.790 11.885 66.110 ;
      LAYER met4 ;
        RECT 11.565 65.790 11.885 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 65.380 11.885 65.700 ;
      LAYER met4 ;
        RECT 11.565 65.380 11.885 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 64.970 11.885 65.290 ;
      LAYER met4 ;
        RECT 11.565 64.970 11.885 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 64.560 11.885 64.880 ;
      LAYER met4 ;
        RECT 11.565 64.560 11.885 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 64.150 11.885 64.470 ;
      LAYER met4 ;
        RECT 11.565 64.150 11.885 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 63.740 11.885 64.060 ;
      LAYER met4 ;
        RECT 11.565 63.740 11.885 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 63.330 11.885 63.650 ;
      LAYER met4 ;
        RECT 11.565 63.330 11.885 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 62.920 11.885 63.240 ;
      LAYER met4 ;
        RECT 11.565 62.920 11.885 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 62.510 11.885 62.830 ;
      LAYER met4 ;
        RECT 11.565 62.510 11.885 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.565 62.100 11.885 62.420 ;
      LAYER met4 ;
        RECT 11.565 62.100 11.885 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 66.200 11.480 66.520 ;
      LAYER met4 ;
        RECT 11.160 66.200 11.480 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 65.790 11.480 66.110 ;
      LAYER met4 ;
        RECT 11.160 65.790 11.480 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 65.380 11.480 65.700 ;
      LAYER met4 ;
        RECT 11.160 65.380 11.480 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 64.970 11.480 65.290 ;
      LAYER met4 ;
        RECT 11.160 64.970 11.480 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 64.560 11.480 64.880 ;
      LAYER met4 ;
        RECT 11.160 64.560 11.480 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 64.150 11.480 64.470 ;
      LAYER met4 ;
        RECT 11.160 64.150 11.480 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 63.740 11.480 64.060 ;
      LAYER met4 ;
        RECT 11.160 63.740 11.480 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 63.330 11.480 63.650 ;
      LAYER met4 ;
        RECT 11.160 63.330 11.480 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 62.920 11.480 63.240 ;
      LAYER met4 ;
        RECT 11.160 62.920 11.480 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 62.510 11.480 62.830 ;
      LAYER met4 ;
        RECT 11.160 62.510 11.480 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.160 62.100 11.480 62.420 ;
      LAYER met4 ;
        RECT 11.160 62.100 11.480 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 66.200 11.075 66.520 ;
      LAYER met4 ;
        RECT 10.755 66.200 11.075 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 65.790 11.075 66.110 ;
      LAYER met4 ;
        RECT 10.755 65.790 11.075 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 65.380 11.075 65.700 ;
      LAYER met4 ;
        RECT 10.755 65.380 11.075 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 64.970 11.075 65.290 ;
      LAYER met4 ;
        RECT 10.755 64.970 11.075 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 64.560 11.075 64.880 ;
      LAYER met4 ;
        RECT 10.755 64.560 11.075 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 64.150 11.075 64.470 ;
      LAYER met4 ;
        RECT 10.755 64.150 11.075 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 63.740 11.075 64.060 ;
      LAYER met4 ;
        RECT 10.755 63.740 11.075 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 63.330 11.075 63.650 ;
      LAYER met4 ;
        RECT 10.755 63.330 11.075 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 62.920 11.075 63.240 ;
      LAYER met4 ;
        RECT 10.755 62.920 11.075 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 62.510 11.075 62.830 ;
      LAYER met4 ;
        RECT 10.755 62.510 11.075 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.755 62.100 11.075 62.420 ;
      LAYER met4 ;
        RECT 10.755 62.100 11.075 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 66.200 10.670 66.520 ;
      LAYER met4 ;
        RECT 10.350 66.200 10.670 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 65.790 10.670 66.110 ;
      LAYER met4 ;
        RECT 10.350 65.790 10.670 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 65.380 10.670 65.700 ;
      LAYER met4 ;
        RECT 10.350 65.380 10.670 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 64.970 10.670 65.290 ;
      LAYER met4 ;
        RECT 10.350 64.970 10.670 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 64.560 10.670 64.880 ;
      LAYER met4 ;
        RECT 10.350 64.560 10.670 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 64.150 10.670 64.470 ;
      LAYER met4 ;
        RECT 10.350 64.150 10.670 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 63.740 10.670 64.060 ;
      LAYER met4 ;
        RECT 10.350 63.740 10.670 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 63.330 10.670 63.650 ;
      LAYER met4 ;
        RECT 10.350 63.330 10.670 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 62.920 10.670 63.240 ;
      LAYER met4 ;
        RECT 10.350 62.920 10.670 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 62.510 10.670 62.830 ;
      LAYER met4 ;
        RECT 10.350 62.510 10.670 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.350 62.100 10.670 62.420 ;
      LAYER met4 ;
        RECT 10.350 62.100 10.670 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 66.200 10.265 66.520 ;
      LAYER met4 ;
        RECT 9.945 66.200 10.265 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 65.790 10.265 66.110 ;
      LAYER met4 ;
        RECT 9.945 65.790 10.265 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 65.380 10.265 65.700 ;
      LAYER met4 ;
        RECT 9.945 65.380 10.265 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 64.970 10.265 65.290 ;
      LAYER met4 ;
        RECT 9.945 64.970 10.265 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 64.560 10.265 64.880 ;
      LAYER met4 ;
        RECT 9.945 64.560 10.265 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 64.150 10.265 64.470 ;
      LAYER met4 ;
        RECT 9.945 64.150 10.265 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 63.740 10.265 64.060 ;
      LAYER met4 ;
        RECT 9.945 63.740 10.265 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 63.330 10.265 63.650 ;
      LAYER met4 ;
        RECT 9.945 63.330 10.265 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 62.920 10.265 63.240 ;
      LAYER met4 ;
        RECT 9.945 62.920 10.265 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 62.510 10.265 62.830 ;
      LAYER met4 ;
        RECT 9.945 62.510 10.265 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.945 62.100 10.265 62.420 ;
      LAYER met4 ;
        RECT 9.945 62.100 10.265 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 66.200 9.860 66.520 ;
      LAYER met4 ;
        RECT 9.540 66.200 9.860 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 65.790 9.860 66.110 ;
      LAYER met4 ;
        RECT 9.540 65.790 9.860 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 65.380 9.860 65.700 ;
      LAYER met4 ;
        RECT 9.540 65.380 9.860 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 64.970 9.860 65.290 ;
      LAYER met4 ;
        RECT 9.540 64.970 9.860 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 64.560 9.860 64.880 ;
      LAYER met4 ;
        RECT 9.540 64.560 9.860 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 64.150 9.860 64.470 ;
      LAYER met4 ;
        RECT 9.540 64.150 9.860 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 63.740 9.860 64.060 ;
      LAYER met4 ;
        RECT 9.540 63.740 9.860 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 63.330 9.860 63.650 ;
      LAYER met4 ;
        RECT 9.540 63.330 9.860 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 62.920 9.860 63.240 ;
      LAYER met4 ;
        RECT 9.540 62.920 9.860 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 62.510 9.860 62.830 ;
      LAYER met4 ;
        RECT 9.540 62.510 9.860 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.540 62.100 9.860 62.420 ;
      LAYER met4 ;
        RECT 9.540 62.100 9.860 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 66.200 9.455 66.520 ;
      LAYER met4 ;
        RECT 9.135 66.200 9.455 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 65.790 9.455 66.110 ;
      LAYER met4 ;
        RECT 9.135 65.790 9.455 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 65.380 9.455 65.700 ;
      LAYER met4 ;
        RECT 9.135 65.380 9.455 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 64.970 9.455 65.290 ;
      LAYER met4 ;
        RECT 9.135 64.970 9.455 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 64.560 9.455 64.880 ;
      LAYER met4 ;
        RECT 9.135 64.560 9.455 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 64.150 9.455 64.470 ;
      LAYER met4 ;
        RECT 9.135 64.150 9.455 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 63.740 9.455 64.060 ;
      LAYER met4 ;
        RECT 9.135 63.740 9.455 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 63.330 9.455 63.650 ;
      LAYER met4 ;
        RECT 9.135 63.330 9.455 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 62.920 9.455 63.240 ;
      LAYER met4 ;
        RECT 9.135 62.920 9.455 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 62.510 9.455 62.830 ;
      LAYER met4 ;
        RECT 9.135 62.510 9.455 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.135 62.100 9.455 62.420 ;
      LAYER met4 ;
        RECT 9.135 62.100 9.455 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 66.200 9.050 66.520 ;
      LAYER met4 ;
        RECT 8.730 66.200 9.050 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 65.790 9.050 66.110 ;
      LAYER met4 ;
        RECT 8.730 65.790 9.050 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 65.380 9.050 65.700 ;
      LAYER met4 ;
        RECT 8.730 65.380 9.050 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 64.970 9.050 65.290 ;
      LAYER met4 ;
        RECT 8.730 64.970 9.050 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 64.560 9.050 64.880 ;
      LAYER met4 ;
        RECT 8.730 64.560 9.050 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 64.150 9.050 64.470 ;
      LAYER met4 ;
        RECT 8.730 64.150 9.050 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 63.740 9.050 64.060 ;
      LAYER met4 ;
        RECT 8.730 63.740 9.050 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 63.330 9.050 63.650 ;
      LAYER met4 ;
        RECT 8.730 63.330 9.050 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 62.920 9.050 63.240 ;
      LAYER met4 ;
        RECT 8.730 62.920 9.050 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 62.510 9.050 62.830 ;
      LAYER met4 ;
        RECT 8.730 62.510 9.050 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.730 62.100 9.050 62.420 ;
      LAYER met4 ;
        RECT 8.730 62.100 9.050 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 66.200 8.645 66.520 ;
      LAYER met4 ;
        RECT 8.325 66.200 8.645 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 65.790 8.645 66.110 ;
      LAYER met4 ;
        RECT 8.325 65.790 8.645 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 65.380 8.645 65.700 ;
      LAYER met4 ;
        RECT 8.325 65.380 8.645 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 64.970 8.645 65.290 ;
      LAYER met4 ;
        RECT 8.325 64.970 8.645 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 64.560 8.645 64.880 ;
      LAYER met4 ;
        RECT 8.325 64.560 8.645 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 64.150 8.645 64.470 ;
      LAYER met4 ;
        RECT 8.325 64.150 8.645 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 63.740 8.645 64.060 ;
      LAYER met4 ;
        RECT 8.325 63.740 8.645 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 63.330 8.645 63.650 ;
      LAYER met4 ;
        RECT 8.325 63.330 8.645 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 62.920 8.645 63.240 ;
      LAYER met4 ;
        RECT 8.325 62.920 8.645 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 62.510 8.645 62.830 ;
      LAYER met4 ;
        RECT 8.325 62.510 8.645 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.325 62.100 8.645 62.420 ;
      LAYER met4 ;
        RECT 8.325 62.100 8.645 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 66.200 8.240 66.520 ;
      LAYER met4 ;
        RECT 7.920 66.200 8.240 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 65.790 8.240 66.110 ;
      LAYER met4 ;
        RECT 7.920 65.790 8.240 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 65.380 8.240 65.700 ;
      LAYER met4 ;
        RECT 7.920 65.380 8.240 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 64.970 8.240 65.290 ;
      LAYER met4 ;
        RECT 7.920 64.970 8.240 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 64.560 8.240 64.880 ;
      LAYER met4 ;
        RECT 7.920 64.560 8.240 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 64.150 8.240 64.470 ;
      LAYER met4 ;
        RECT 7.920 64.150 8.240 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 63.740 8.240 64.060 ;
      LAYER met4 ;
        RECT 7.920 63.740 8.240 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 63.330 8.240 63.650 ;
      LAYER met4 ;
        RECT 7.920 63.330 8.240 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 62.920 8.240 63.240 ;
      LAYER met4 ;
        RECT 7.920 62.920 8.240 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 62.510 8.240 62.830 ;
      LAYER met4 ;
        RECT 7.920 62.510 8.240 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.920 62.100 8.240 62.420 ;
      LAYER met4 ;
        RECT 7.920 62.100 8.240 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 66.200 7.835 66.520 ;
      LAYER met4 ;
        RECT 7.515 66.200 7.835 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 65.790 7.835 66.110 ;
      LAYER met4 ;
        RECT 7.515 65.790 7.835 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 65.380 7.835 65.700 ;
      LAYER met4 ;
        RECT 7.515 65.380 7.835 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 64.970 7.835 65.290 ;
      LAYER met4 ;
        RECT 7.515 64.970 7.835 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 64.560 7.835 64.880 ;
      LAYER met4 ;
        RECT 7.515 64.560 7.835 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 64.150 7.835 64.470 ;
      LAYER met4 ;
        RECT 7.515 64.150 7.835 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 63.740 7.835 64.060 ;
      LAYER met4 ;
        RECT 7.515 63.740 7.835 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 63.330 7.835 63.650 ;
      LAYER met4 ;
        RECT 7.515 63.330 7.835 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 62.920 7.835 63.240 ;
      LAYER met4 ;
        RECT 7.515 62.920 7.835 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 62.510 7.835 62.830 ;
      LAYER met4 ;
        RECT 7.515 62.510 7.835 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.515 62.100 7.835 62.420 ;
      LAYER met4 ;
        RECT 7.515 62.100 7.835 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 66.200 7.430 66.520 ;
      LAYER met4 ;
        RECT 7.110 66.200 7.430 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 65.790 7.430 66.110 ;
      LAYER met4 ;
        RECT 7.110 65.790 7.430 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 65.380 7.430 65.700 ;
      LAYER met4 ;
        RECT 7.110 65.380 7.430 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 64.970 7.430 65.290 ;
      LAYER met4 ;
        RECT 7.110 64.970 7.430 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 64.560 7.430 64.880 ;
      LAYER met4 ;
        RECT 7.110 64.560 7.430 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 64.150 7.430 64.470 ;
      LAYER met4 ;
        RECT 7.110 64.150 7.430 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 63.740 7.430 64.060 ;
      LAYER met4 ;
        RECT 7.110 63.740 7.430 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 63.330 7.430 63.650 ;
      LAYER met4 ;
        RECT 7.110 63.330 7.430 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 62.920 7.430 63.240 ;
      LAYER met4 ;
        RECT 7.110 62.920 7.430 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 62.510 7.430 62.830 ;
      LAYER met4 ;
        RECT 7.110 62.510 7.430 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.110 62.100 7.430 62.420 ;
      LAYER met4 ;
        RECT 7.110 62.100 7.430 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 66.200 7.025 66.520 ;
      LAYER met4 ;
        RECT 6.705 66.200 7.025 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 65.790 7.025 66.110 ;
      LAYER met4 ;
        RECT 6.705 65.790 7.025 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 65.380 7.025 65.700 ;
      LAYER met4 ;
        RECT 6.705 65.380 7.025 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 64.970 7.025 65.290 ;
      LAYER met4 ;
        RECT 6.705 64.970 7.025 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 64.560 7.025 64.880 ;
      LAYER met4 ;
        RECT 6.705 64.560 7.025 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 64.150 7.025 64.470 ;
      LAYER met4 ;
        RECT 6.705 64.150 7.025 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 63.740 7.025 64.060 ;
      LAYER met4 ;
        RECT 6.705 63.740 7.025 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 63.330 7.025 63.650 ;
      LAYER met4 ;
        RECT 6.705 63.330 7.025 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 62.920 7.025 63.240 ;
      LAYER met4 ;
        RECT 6.705 62.920 7.025 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 62.510 7.025 62.830 ;
      LAYER met4 ;
        RECT 6.705 62.510 7.025 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.705 62.100 7.025 62.420 ;
      LAYER met4 ;
        RECT 6.705 62.100 7.025 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 66.200 6.620 66.520 ;
      LAYER met4 ;
        RECT 6.300 66.200 6.620 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 65.790 6.620 66.110 ;
      LAYER met4 ;
        RECT 6.300 65.790 6.620 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 65.380 6.620 65.700 ;
      LAYER met4 ;
        RECT 6.300 65.380 6.620 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 64.970 6.620 65.290 ;
      LAYER met4 ;
        RECT 6.300 64.970 6.620 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 64.560 6.620 64.880 ;
      LAYER met4 ;
        RECT 6.300 64.560 6.620 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 64.150 6.620 64.470 ;
      LAYER met4 ;
        RECT 6.300 64.150 6.620 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 63.740 6.620 64.060 ;
      LAYER met4 ;
        RECT 6.300 63.740 6.620 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 63.330 6.620 63.650 ;
      LAYER met4 ;
        RECT 6.300 63.330 6.620 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 62.920 6.620 63.240 ;
      LAYER met4 ;
        RECT 6.300 62.920 6.620 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 62.510 6.620 62.830 ;
      LAYER met4 ;
        RECT 6.300 62.510 6.620 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.300 62.100 6.620 62.420 ;
      LAYER met4 ;
        RECT 6.300 62.100 6.620 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 66.200 6.215 66.520 ;
      LAYER met4 ;
        RECT 5.895 66.200 6.215 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 65.790 6.215 66.110 ;
      LAYER met4 ;
        RECT 5.895 65.790 6.215 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 65.380 6.215 65.700 ;
      LAYER met4 ;
        RECT 5.895 65.380 6.215 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 64.970 6.215 65.290 ;
      LAYER met4 ;
        RECT 5.895 64.970 6.215 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 64.560 6.215 64.880 ;
      LAYER met4 ;
        RECT 5.895 64.560 6.215 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 64.150 6.215 64.470 ;
      LAYER met4 ;
        RECT 5.895 64.150 6.215 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 63.740 6.215 64.060 ;
      LAYER met4 ;
        RECT 5.895 63.740 6.215 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 63.330 6.215 63.650 ;
      LAYER met4 ;
        RECT 5.895 63.330 6.215 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 62.920 6.215 63.240 ;
      LAYER met4 ;
        RECT 5.895 62.920 6.215 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 62.510 6.215 62.830 ;
      LAYER met4 ;
        RECT 5.895 62.510 6.215 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.895 62.100 6.215 62.420 ;
      LAYER met4 ;
        RECT 5.895 62.100 6.215 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 66.200 5.810 66.520 ;
      LAYER met4 ;
        RECT 5.490 66.200 5.810 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 65.790 5.810 66.110 ;
      LAYER met4 ;
        RECT 5.490 65.790 5.810 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 65.380 5.810 65.700 ;
      LAYER met4 ;
        RECT 5.490 65.380 5.810 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 64.970 5.810 65.290 ;
      LAYER met4 ;
        RECT 5.490 64.970 5.810 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 64.560 5.810 64.880 ;
      LAYER met4 ;
        RECT 5.490 64.560 5.810 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 64.150 5.810 64.470 ;
      LAYER met4 ;
        RECT 5.490 64.150 5.810 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 63.740 5.810 64.060 ;
      LAYER met4 ;
        RECT 5.490 63.740 5.810 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 63.330 5.810 63.650 ;
      LAYER met4 ;
        RECT 5.490 63.330 5.810 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 62.920 5.810 63.240 ;
      LAYER met4 ;
        RECT 5.490 62.920 5.810 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 62.510 5.810 62.830 ;
      LAYER met4 ;
        RECT 5.490 62.510 5.810 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.490 62.100 5.810 62.420 ;
      LAYER met4 ;
        RECT 5.490 62.100 5.810 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 66.200 5.405 66.520 ;
      LAYER met4 ;
        RECT 5.085 66.200 5.405 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 65.790 5.405 66.110 ;
      LAYER met4 ;
        RECT 5.085 65.790 5.405 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 65.380 5.405 65.700 ;
      LAYER met4 ;
        RECT 5.085 65.380 5.405 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 64.970 5.405 65.290 ;
      LAYER met4 ;
        RECT 5.085 64.970 5.405 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 64.560 5.405 64.880 ;
      LAYER met4 ;
        RECT 5.085 64.560 5.405 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 64.150 5.405 64.470 ;
      LAYER met4 ;
        RECT 5.085 64.150 5.405 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 63.740 5.405 64.060 ;
      LAYER met4 ;
        RECT 5.085 63.740 5.405 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 63.330 5.405 63.650 ;
      LAYER met4 ;
        RECT 5.085 63.330 5.405 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 62.920 5.405 63.240 ;
      LAYER met4 ;
        RECT 5.085 62.920 5.405 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 62.510 5.405 62.830 ;
      LAYER met4 ;
        RECT 5.085 62.510 5.405 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.085 62.100 5.405 62.420 ;
      LAYER met4 ;
        RECT 5.085 62.100 5.405 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 66.200 5.000 66.520 ;
      LAYER met4 ;
        RECT 4.680 66.200 5.000 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 65.790 5.000 66.110 ;
      LAYER met4 ;
        RECT 4.680 65.790 5.000 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 65.380 5.000 65.700 ;
      LAYER met4 ;
        RECT 4.680 65.380 5.000 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 64.970 5.000 65.290 ;
      LAYER met4 ;
        RECT 4.680 64.970 5.000 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 64.560 5.000 64.880 ;
      LAYER met4 ;
        RECT 4.680 64.560 5.000 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 64.150 5.000 64.470 ;
      LAYER met4 ;
        RECT 4.680 64.150 5.000 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 63.740 5.000 64.060 ;
      LAYER met4 ;
        RECT 4.680 63.740 5.000 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 63.330 5.000 63.650 ;
      LAYER met4 ;
        RECT 4.680 63.330 5.000 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 62.920 5.000 63.240 ;
      LAYER met4 ;
        RECT 4.680 62.920 5.000 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 62.510 5.000 62.830 ;
      LAYER met4 ;
        RECT 4.680 62.510 5.000 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.680 62.100 5.000 62.420 ;
      LAYER met4 ;
        RECT 4.680 62.100 5.000 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 66.200 4.595 66.520 ;
      LAYER met4 ;
        RECT 4.275 66.200 4.595 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 65.790 4.595 66.110 ;
      LAYER met4 ;
        RECT 4.275 65.790 4.595 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 65.380 4.595 65.700 ;
      LAYER met4 ;
        RECT 4.275 65.380 4.595 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 64.970 4.595 65.290 ;
      LAYER met4 ;
        RECT 4.275 64.970 4.595 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 64.560 4.595 64.880 ;
      LAYER met4 ;
        RECT 4.275 64.560 4.595 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 64.150 4.595 64.470 ;
      LAYER met4 ;
        RECT 4.275 64.150 4.595 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 63.740 4.595 64.060 ;
      LAYER met4 ;
        RECT 4.275 63.740 4.595 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 63.330 4.595 63.650 ;
      LAYER met4 ;
        RECT 4.275 63.330 4.595 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 62.920 4.595 63.240 ;
      LAYER met4 ;
        RECT 4.275 62.920 4.595 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 62.510 4.595 62.830 ;
      LAYER met4 ;
        RECT 4.275 62.510 4.595 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.275 62.100 4.595 62.420 ;
      LAYER met4 ;
        RECT 4.275 62.100 4.595 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 66.200 4.190 66.520 ;
      LAYER met4 ;
        RECT 3.870 66.200 4.190 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 65.790 4.190 66.110 ;
      LAYER met4 ;
        RECT 3.870 65.790 4.190 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 65.380 4.190 65.700 ;
      LAYER met4 ;
        RECT 3.870 65.380 4.190 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 64.970 4.190 65.290 ;
      LAYER met4 ;
        RECT 3.870 64.970 4.190 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 64.560 4.190 64.880 ;
      LAYER met4 ;
        RECT 3.870 64.560 4.190 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 64.150 4.190 64.470 ;
      LAYER met4 ;
        RECT 3.870 64.150 4.190 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 63.740 4.190 64.060 ;
      LAYER met4 ;
        RECT 3.870 63.740 4.190 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 63.330 4.190 63.650 ;
      LAYER met4 ;
        RECT 3.870 63.330 4.190 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 62.920 4.190 63.240 ;
      LAYER met4 ;
        RECT 3.870 62.920 4.190 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 62.510 4.190 62.830 ;
      LAYER met4 ;
        RECT 3.870 62.510 4.190 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.870 62.100 4.190 62.420 ;
      LAYER met4 ;
        RECT 3.870 62.100 4.190 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 66.200 3.785 66.520 ;
      LAYER met4 ;
        RECT 3.465 66.200 3.785 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 65.790 3.785 66.110 ;
      LAYER met4 ;
        RECT 3.465 65.790 3.785 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 65.380 3.785 65.700 ;
      LAYER met4 ;
        RECT 3.465 65.380 3.785 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 64.970 3.785 65.290 ;
      LAYER met4 ;
        RECT 3.465 64.970 3.785 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 64.560 3.785 64.880 ;
      LAYER met4 ;
        RECT 3.465 64.560 3.785 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 64.150 3.785 64.470 ;
      LAYER met4 ;
        RECT 3.465 64.150 3.785 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 63.740 3.785 64.060 ;
      LAYER met4 ;
        RECT 3.465 63.740 3.785 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 63.330 3.785 63.650 ;
      LAYER met4 ;
        RECT 3.465 63.330 3.785 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 62.920 3.785 63.240 ;
      LAYER met4 ;
        RECT 3.465 62.920 3.785 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 62.510 3.785 62.830 ;
      LAYER met4 ;
        RECT 3.465 62.510 3.785 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.465 62.100 3.785 62.420 ;
      LAYER met4 ;
        RECT 3.465 62.100 3.785 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 66.200 3.380 66.520 ;
      LAYER met4 ;
        RECT 3.060 66.200 3.380 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 65.790 3.380 66.110 ;
      LAYER met4 ;
        RECT 3.060 65.790 3.380 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 65.380 3.380 65.700 ;
      LAYER met4 ;
        RECT 3.060 65.380 3.380 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 64.970 3.380 65.290 ;
      LAYER met4 ;
        RECT 3.060 64.970 3.380 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 64.560 3.380 64.880 ;
      LAYER met4 ;
        RECT 3.060 64.560 3.380 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 64.150 3.380 64.470 ;
      LAYER met4 ;
        RECT 3.060 64.150 3.380 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 63.740 3.380 64.060 ;
      LAYER met4 ;
        RECT 3.060 63.740 3.380 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 63.330 3.380 63.650 ;
      LAYER met4 ;
        RECT 3.060 63.330 3.380 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 62.920 3.380 63.240 ;
      LAYER met4 ;
        RECT 3.060 62.920 3.380 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 62.510 3.380 62.830 ;
      LAYER met4 ;
        RECT 3.060 62.510 3.380 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.060 62.100 3.380 62.420 ;
      LAYER met4 ;
        RECT 3.060 62.100 3.380 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 66.200 2.975 66.520 ;
      LAYER met4 ;
        RECT 2.655 66.200 2.975 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 65.790 2.975 66.110 ;
      LAYER met4 ;
        RECT 2.655 65.790 2.975 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 65.380 2.975 65.700 ;
      LAYER met4 ;
        RECT 2.655 65.380 2.975 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 64.970 2.975 65.290 ;
      LAYER met4 ;
        RECT 2.655 64.970 2.975 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 64.560 2.975 64.880 ;
      LAYER met4 ;
        RECT 2.655 64.560 2.975 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 64.150 2.975 64.470 ;
      LAYER met4 ;
        RECT 2.655 64.150 2.975 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 63.740 2.975 64.060 ;
      LAYER met4 ;
        RECT 2.655 63.740 2.975 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 63.330 2.975 63.650 ;
      LAYER met4 ;
        RECT 2.655 63.330 2.975 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 62.920 2.975 63.240 ;
      LAYER met4 ;
        RECT 2.655 62.920 2.975 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 62.510 2.975 62.830 ;
      LAYER met4 ;
        RECT 2.655 62.510 2.975 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.655 62.100 2.975 62.420 ;
      LAYER met4 ;
        RECT 2.655 62.100 2.975 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 66.200 2.570 66.520 ;
      LAYER met4 ;
        RECT 2.250 66.200 2.570 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 65.790 2.570 66.110 ;
      LAYER met4 ;
        RECT 2.250 65.790 2.570 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 65.380 2.570 65.700 ;
      LAYER met4 ;
        RECT 2.250 65.380 2.570 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 64.970 2.570 65.290 ;
      LAYER met4 ;
        RECT 2.250 64.970 2.570 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 64.560 2.570 64.880 ;
      LAYER met4 ;
        RECT 2.250 64.560 2.570 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 64.150 2.570 64.470 ;
      LAYER met4 ;
        RECT 2.250 64.150 2.570 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 63.740 2.570 64.060 ;
      LAYER met4 ;
        RECT 2.250 63.740 2.570 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 63.330 2.570 63.650 ;
      LAYER met4 ;
        RECT 2.250 63.330 2.570 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 62.920 2.570 63.240 ;
      LAYER met4 ;
        RECT 2.250 62.920 2.570 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 62.510 2.570 62.830 ;
      LAYER met4 ;
        RECT 2.250 62.510 2.570 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.250 62.100 2.570 62.420 ;
      LAYER met4 ;
        RECT 2.250 62.100 2.570 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 66.200 2.165 66.520 ;
      LAYER met4 ;
        RECT 1.845 66.200 2.165 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 65.790 2.165 66.110 ;
      LAYER met4 ;
        RECT 1.845 65.790 2.165 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 65.380 2.165 65.700 ;
      LAYER met4 ;
        RECT 1.845 65.380 2.165 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 64.970 2.165 65.290 ;
      LAYER met4 ;
        RECT 1.845 64.970 2.165 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 64.560 2.165 64.880 ;
      LAYER met4 ;
        RECT 1.845 64.560 2.165 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 64.150 2.165 64.470 ;
      LAYER met4 ;
        RECT 1.845 64.150 2.165 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 63.740 2.165 64.060 ;
      LAYER met4 ;
        RECT 1.845 63.740 2.165 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 63.330 2.165 63.650 ;
      LAYER met4 ;
        RECT 1.845 63.330 2.165 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 62.920 2.165 63.240 ;
      LAYER met4 ;
        RECT 1.845 62.920 2.165 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 62.510 2.165 62.830 ;
      LAYER met4 ;
        RECT 1.845 62.510 2.165 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.845 62.100 2.165 62.420 ;
      LAYER met4 ;
        RECT 1.845 62.100 2.165 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 66.200 1.760 66.520 ;
      LAYER met4 ;
        RECT 1.440 66.200 1.760 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 65.790 1.760 66.110 ;
      LAYER met4 ;
        RECT 1.440 65.790 1.760 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 65.380 1.760 65.700 ;
      LAYER met4 ;
        RECT 1.440 65.380 1.760 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 64.970 1.760 65.290 ;
      LAYER met4 ;
        RECT 1.440 64.970 1.760 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 64.560 1.760 64.880 ;
      LAYER met4 ;
        RECT 1.440 64.560 1.760 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 64.150 1.760 64.470 ;
      LAYER met4 ;
        RECT 1.440 64.150 1.760 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 63.740 1.760 64.060 ;
      LAYER met4 ;
        RECT 1.440 63.740 1.760 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 63.330 1.760 63.650 ;
      LAYER met4 ;
        RECT 1.440 63.330 1.760 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 62.920 1.760 63.240 ;
      LAYER met4 ;
        RECT 1.440 62.920 1.760 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 62.510 1.760 62.830 ;
      LAYER met4 ;
        RECT 1.440 62.510 1.760 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.440 62.100 1.760 62.420 ;
      LAYER met4 ;
        RECT 1.440 62.100 1.760 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 66.200 1.355 66.520 ;
      LAYER met4 ;
        RECT 1.270 66.200 1.355 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 65.790 1.355 66.110 ;
      LAYER met4 ;
        RECT 1.270 65.790 1.355 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 65.380 1.355 65.700 ;
      LAYER met4 ;
        RECT 1.270 65.380 1.355 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 64.970 1.355 65.290 ;
      LAYER met4 ;
        RECT 1.270 64.970 1.355 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 64.560 1.355 64.880 ;
      LAYER met4 ;
        RECT 1.270 64.560 1.355 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 64.150 1.355 64.470 ;
      LAYER met4 ;
        RECT 1.270 64.150 1.355 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 63.740 1.355 64.060 ;
      LAYER met4 ;
        RECT 1.270 63.740 1.355 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 63.330 1.355 63.650 ;
      LAYER met4 ;
        RECT 1.270 63.330 1.355 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 62.920 1.355 63.240 ;
      LAYER met4 ;
        RECT 1.270 62.920 1.355 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 62.510 1.355 62.830 ;
      LAYER met4 ;
        RECT 1.270 62.510 1.355 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.035 62.100 1.355 62.420 ;
      LAYER met4 ;
        RECT 1.270 62.100 1.355 62.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 66.200 0.950 66.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 65.790 0.950 66.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 65.380 0.950 65.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 64.970 0.950 65.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 64.560 0.950 64.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 64.150 0.950 64.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 63.740 0.950 64.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 63.330 0.950 63.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 62.920 0.950 63.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 62.510 0.950 62.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.630 62.100 0.950 62.420 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
  END VSSD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.600 17.790 24.500 22.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 17.790 74.655 22.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.055 92.865 74.660 92.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 91.735 61.055 92.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.940 90.845 59.830 91.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.650 89.555 58.940 90.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.260 88.165 57.650 89.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.135 87.040 56.260 88.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 85.615 55.135 87.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.405 84.310 53.710 85.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.760 82.665 52.405 84.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.760 68.035 74.660 82.665 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.255 90.950 15.365 91.710 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.270 88.345 16.250 90.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.375 82.990 18.855 88.140 ;
    END
    PORT
      LAYER met4 ;
        RECT 16.415 88.365 17.525 89.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.995 85.810 20.065 87.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.170 82.945 21.450 85.590 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.650 82.855 22.770 84.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 52.485 82.855 53.605 84.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.805 82.945 56.085 85.590 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.190 85.810 56.260 87.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.400 82.990 60.880 88.140 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.730 88.365 58.840 89.530 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.005 88.345 60.985 90.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 59.890 90.950 61.000 91.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 22.160 74.565 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 21.730 74.565 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 21.300 74.565 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 20.870 74.565 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 20.440 74.565 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 20.010 74.565 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 19.580 74.565 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 19.150 74.565 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 18.720 74.565 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 18.290 74.565 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 17.860 74.565 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.320 92.695 74.520 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 92.225 74.580 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 91.815 74.580 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 91.405 74.580 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 90.995 74.580 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 90.585 74.580 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 90.175 74.580 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 89.765 74.580 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 89.355 74.580 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 88.945 74.580 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 88.535 74.580 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 88.125 74.580 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 87.715 74.580 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 87.305 74.580 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 86.895 74.580 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 86.485 74.580 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 86.075 74.580 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 85.665 74.580 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 85.255 74.580 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 84.845 74.580 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 84.435 74.580 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 84.025 74.580 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 83.615 74.580 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 83.205 74.580 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.260 82.795 74.580 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 82.360 74.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 81.955 74.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 81.550 74.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 81.145 74.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 80.740 74.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 80.335 74.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 79.930 74.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 79.525 74.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 79.120 74.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 78.715 74.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 78.310 74.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 77.905 74.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 77.500 74.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 77.095 74.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 76.690 74.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 76.285 74.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 75.880 74.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 75.475 74.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 75.070 74.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 74.665 74.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 74.260 74.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 73.855 74.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 73.450 74.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 73.045 74.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 72.635 74.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 72.225 74.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 71.815 74.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 71.405 74.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 70.995 74.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 70.585 74.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 70.175 74.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 69.765 74.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 69.355 74.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 68.945 74.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 68.535 74.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.210 68.125 74.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 22.160 74.155 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 21.730 74.155 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 21.300 74.155 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 20.870 74.155 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 20.440 74.155 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 20.010 74.155 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 19.580 74.155 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 19.150 74.155 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 18.720 74.155 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 18.290 74.155 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 17.860 74.155 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.910 92.695 74.110 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 92.225 74.170 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 91.815 74.170 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 91.405 74.170 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 90.995 74.170 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 90.585 74.170 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 90.175 74.170 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 89.765 74.170 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 89.355 74.170 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 88.945 74.170 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 88.535 74.170 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 88.125 74.170 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 87.715 74.170 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 87.305 74.170 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 86.895 74.170 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 86.485 74.170 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 86.075 74.170 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 85.665 74.170 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 85.255 74.170 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 84.845 74.170 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 84.435 74.170 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 84.025 74.170 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 83.615 74.170 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 83.205 74.170 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.850 82.795 74.170 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 82.360 74.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 81.955 74.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 81.550 74.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 81.145 74.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 80.740 74.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 80.335 74.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 79.930 74.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 79.525 74.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 79.120 74.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 78.715 74.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 78.310 74.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 77.905 74.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 77.500 74.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 77.095 74.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 76.690 74.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 76.285 74.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 75.880 74.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 75.475 74.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 75.070 74.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 74.665 74.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 74.260 74.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 73.855 74.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 73.450 74.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 73.045 74.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 72.635 74.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 72.225 74.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 71.815 74.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 71.405 74.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 70.995 74.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 70.585 74.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 70.175 74.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 69.765 74.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 69.355 74.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 68.945 74.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 68.535 74.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.810 68.125 74.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 22.160 73.745 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 21.730 73.745 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 21.300 73.745 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 20.870 73.745 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 20.440 73.745 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 20.010 73.745 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 19.580 73.745 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 19.150 73.745 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 18.720 73.745 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 18.290 73.745 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.545 17.860 73.745 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.500 92.695 73.700 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 92.225 73.760 92.545 ;
      LAYER met4 ;
        RECT 73.440 92.225 73.730 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 91.815 73.760 92.135 ;
      LAYER met4 ;
        RECT 73.440 91.815 73.730 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 91.405 73.760 91.725 ;
      LAYER met4 ;
        RECT 73.440 91.405 73.730 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 90.995 73.760 91.315 ;
      LAYER met4 ;
        RECT 73.440 90.995 73.730 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 90.585 73.760 90.905 ;
      LAYER met4 ;
        RECT 73.440 90.585 73.730 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 90.175 73.760 90.495 ;
      LAYER met4 ;
        RECT 73.440 90.175 73.730 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 89.765 73.760 90.085 ;
      LAYER met4 ;
        RECT 73.440 89.765 73.730 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 89.355 73.760 89.675 ;
      LAYER met4 ;
        RECT 73.440 89.355 73.730 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 88.945 73.760 89.265 ;
      LAYER met4 ;
        RECT 73.440 88.945 73.730 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 88.535 73.760 88.855 ;
      LAYER met4 ;
        RECT 73.440 88.535 73.730 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 88.125 73.760 88.445 ;
      LAYER met4 ;
        RECT 73.440 88.125 73.730 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 87.715 73.760 88.035 ;
      LAYER met4 ;
        RECT 73.440 87.715 73.730 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 87.305 73.760 87.625 ;
      LAYER met4 ;
        RECT 73.440 87.305 73.730 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 86.895 73.760 87.215 ;
      LAYER met4 ;
        RECT 73.440 86.895 73.730 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 86.485 73.760 86.805 ;
      LAYER met4 ;
        RECT 73.440 86.485 73.730 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 86.075 73.760 86.395 ;
      LAYER met4 ;
        RECT 73.440 86.075 73.730 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 85.665 73.760 85.985 ;
      LAYER met4 ;
        RECT 73.440 85.665 73.730 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 85.255 73.760 85.575 ;
      LAYER met4 ;
        RECT 73.440 85.255 73.730 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 84.845 73.760 85.165 ;
      LAYER met4 ;
        RECT 73.440 84.845 73.730 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 84.435 73.760 84.755 ;
      LAYER met4 ;
        RECT 73.440 84.435 73.730 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 84.025 73.760 84.345 ;
      LAYER met4 ;
        RECT 73.440 84.025 73.730 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 83.615 73.760 83.935 ;
      LAYER met4 ;
        RECT 73.440 83.615 73.730 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 83.205 73.760 83.525 ;
      LAYER met4 ;
        RECT 73.440 83.205 73.730 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.440 82.795 73.760 83.115 ;
      LAYER met4 ;
        RECT 73.440 82.795 73.730 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 82.360 73.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 81.955 73.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 81.550 73.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 81.145 73.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 80.740 73.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 80.335 73.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 79.930 73.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 79.525 73.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 79.120 73.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 78.715 73.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 78.310 73.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 77.905 73.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 77.500 73.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 77.095 73.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 76.690 73.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 76.285 73.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 75.880 73.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 75.475 73.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 75.070 73.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 74.665 73.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 74.260 73.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 73.855 73.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 73.450 73.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 73.045 73.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 72.635 73.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 72.225 73.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 71.815 73.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 71.405 73.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 70.995 73.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 70.585 73.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 70.175 73.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 69.765 73.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 69.355 73.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 68.945 73.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 68.535 73.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.410 68.125 73.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 22.160 73.335 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 21.730 73.335 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 21.300 73.335 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 20.870 73.335 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 20.440 73.335 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 20.010 73.335 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 19.580 73.335 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 19.150 73.335 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 18.720 73.335 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 18.290 73.335 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.135 17.860 73.335 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.090 92.695 73.290 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 92.225 73.350 92.545 ;
      LAYER met4 ;
        RECT 73.030 92.225 73.350 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 91.815 73.350 92.135 ;
      LAYER met4 ;
        RECT 73.030 91.815 73.350 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 91.405 73.350 91.725 ;
      LAYER met4 ;
        RECT 73.030 91.405 73.350 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 90.995 73.350 91.315 ;
      LAYER met4 ;
        RECT 73.030 90.995 73.350 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 90.585 73.350 90.905 ;
      LAYER met4 ;
        RECT 73.030 90.585 73.350 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 90.175 73.350 90.495 ;
      LAYER met4 ;
        RECT 73.030 90.175 73.350 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 89.765 73.350 90.085 ;
      LAYER met4 ;
        RECT 73.030 89.765 73.350 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 89.355 73.350 89.675 ;
      LAYER met4 ;
        RECT 73.030 89.355 73.350 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 88.945 73.350 89.265 ;
      LAYER met4 ;
        RECT 73.030 88.945 73.350 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 88.535 73.350 88.855 ;
      LAYER met4 ;
        RECT 73.030 88.535 73.350 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 88.125 73.350 88.445 ;
      LAYER met4 ;
        RECT 73.030 88.125 73.350 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 87.715 73.350 88.035 ;
      LAYER met4 ;
        RECT 73.030 87.715 73.350 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 87.305 73.350 87.625 ;
      LAYER met4 ;
        RECT 73.030 87.305 73.350 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 86.895 73.350 87.215 ;
      LAYER met4 ;
        RECT 73.030 86.895 73.350 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 86.485 73.350 86.805 ;
      LAYER met4 ;
        RECT 73.030 86.485 73.350 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 86.075 73.350 86.395 ;
      LAYER met4 ;
        RECT 73.030 86.075 73.350 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 85.665 73.350 85.985 ;
      LAYER met4 ;
        RECT 73.030 85.665 73.350 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 85.255 73.350 85.575 ;
      LAYER met4 ;
        RECT 73.030 85.255 73.350 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 84.845 73.350 85.165 ;
      LAYER met4 ;
        RECT 73.030 84.845 73.350 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 84.435 73.350 84.755 ;
      LAYER met4 ;
        RECT 73.030 84.435 73.350 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 84.025 73.350 84.345 ;
      LAYER met4 ;
        RECT 73.030 84.025 73.350 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 83.615 73.350 83.935 ;
      LAYER met4 ;
        RECT 73.030 83.615 73.350 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 83.205 73.350 83.525 ;
      LAYER met4 ;
        RECT 73.030 83.205 73.350 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.030 82.795 73.350 83.115 ;
      LAYER met4 ;
        RECT 73.030 82.795 73.350 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 82.360 73.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 81.955 73.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 81.550 73.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 81.145 73.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 80.740 73.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 80.335 73.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 79.930 73.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 79.525 73.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 79.120 73.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 78.715 73.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 78.310 73.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 77.905 73.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 77.500 73.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 77.095 73.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 76.690 73.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 76.285 73.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 75.880 73.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 75.475 73.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 75.070 73.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 74.665 73.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 74.260 73.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 73.855 73.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 73.450 73.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 73.045 73.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 72.635 73.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 72.225 73.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 71.815 73.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 71.405 73.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 70.995 73.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 70.585 73.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 70.175 73.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 69.765 73.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 69.355 73.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 68.945 73.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 68.535 73.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.010 68.125 73.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 22.160 72.925 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 21.730 72.925 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 21.300 72.925 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 20.870 72.925 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 20.440 72.925 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 20.010 72.925 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 19.580 72.925 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 19.150 72.925 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 18.720 72.925 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 18.290 72.925 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 17.860 72.925 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.680 92.695 72.880 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 92.225 72.940 92.545 ;
      LAYER met4 ;
        RECT 72.620 92.225 72.940 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 91.815 72.940 92.135 ;
      LAYER met4 ;
        RECT 72.620 91.815 72.940 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 91.405 72.940 91.725 ;
      LAYER met4 ;
        RECT 72.620 91.405 72.940 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 90.995 72.940 91.315 ;
      LAYER met4 ;
        RECT 72.620 90.995 72.940 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 90.585 72.940 90.905 ;
      LAYER met4 ;
        RECT 72.620 90.585 72.940 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 90.175 72.940 90.495 ;
      LAYER met4 ;
        RECT 72.620 90.175 72.940 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 89.765 72.940 90.085 ;
      LAYER met4 ;
        RECT 72.620 89.765 72.940 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 89.355 72.940 89.675 ;
      LAYER met4 ;
        RECT 72.620 89.355 72.940 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 88.945 72.940 89.265 ;
      LAYER met4 ;
        RECT 72.620 88.945 72.940 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 88.535 72.940 88.855 ;
      LAYER met4 ;
        RECT 72.620 88.535 72.940 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 88.125 72.940 88.445 ;
      LAYER met4 ;
        RECT 72.620 88.125 72.940 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 87.715 72.940 88.035 ;
      LAYER met4 ;
        RECT 72.620 87.715 72.940 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 87.305 72.940 87.625 ;
      LAYER met4 ;
        RECT 72.620 87.305 72.940 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 86.895 72.940 87.215 ;
      LAYER met4 ;
        RECT 72.620 86.895 72.940 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 86.485 72.940 86.805 ;
      LAYER met4 ;
        RECT 72.620 86.485 72.940 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 86.075 72.940 86.395 ;
      LAYER met4 ;
        RECT 72.620 86.075 72.940 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 85.665 72.940 85.985 ;
      LAYER met4 ;
        RECT 72.620 85.665 72.940 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 85.255 72.940 85.575 ;
      LAYER met4 ;
        RECT 72.620 85.255 72.940 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 84.845 72.940 85.165 ;
      LAYER met4 ;
        RECT 72.620 84.845 72.940 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 84.435 72.940 84.755 ;
      LAYER met4 ;
        RECT 72.620 84.435 72.940 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 84.025 72.940 84.345 ;
      LAYER met4 ;
        RECT 72.620 84.025 72.940 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 83.615 72.940 83.935 ;
      LAYER met4 ;
        RECT 72.620 83.615 72.940 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 83.205 72.940 83.525 ;
      LAYER met4 ;
        RECT 72.620 83.205 72.940 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.620 82.795 72.940 83.115 ;
      LAYER met4 ;
        RECT 72.620 82.795 72.940 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 82.360 72.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 81.955 72.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 81.550 72.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 81.145 72.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 80.740 72.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 80.335 72.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 79.930 72.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 79.525 72.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 79.120 72.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 78.715 72.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 78.310 72.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 77.905 72.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 77.500 72.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 77.095 72.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 76.690 72.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 76.285 72.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 75.880 72.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 75.475 72.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 75.070 72.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 74.665 72.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 74.260 72.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 73.855 72.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 73.450 72.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 73.045 72.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 72.635 72.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 72.225 72.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 71.815 72.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 71.405 72.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 70.995 72.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 70.585 72.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 70.175 72.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 69.765 72.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 69.355 72.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 68.945 72.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 68.535 72.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.610 68.125 72.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 22.160 72.515 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 21.730 72.515 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 21.300 72.515 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 20.870 72.515 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 20.440 72.515 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 20.010 72.515 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 19.580 72.515 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 19.150 72.515 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 18.720 72.515 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 18.290 72.515 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.315 17.860 72.515 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.270 92.695 72.470 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 92.225 72.530 92.545 ;
      LAYER met4 ;
        RECT 72.210 92.225 72.530 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 91.815 72.530 92.135 ;
      LAYER met4 ;
        RECT 72.210 91.815 72.530 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 91.405 72.530 91.725 ;
      LAYER met4 ;
        RECT 72.210 91.405 72.530 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 90.995 72.530 91.315 ;
      LAYER met4 ;
        RECT 72.210 90.995 72.530 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 90.585 72.530 90.905 ;
      LAYER met4 ;
        RECT 72.210 90.585 72.530 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 90.175 72.530 90.495 ;
      LAYER met4 ;
        RECT 72.210 90.175 72.530 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 89.765 72.530 90.085 ;
      LAYER met4 ;
        RECT 72.210 89.765 72.530 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 89.355 72.530 89.675 ;
      LAYER met4 ;
        RECT 72.210 89.355 72.530 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 88.945 72.530 89.265 ;
      LAYER met4 ;
        RECT 72.210 88.945 72.530 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 88.535 72.530 88.855 ;
      LAYER met4 ;
        RECT 72.210 88.535 72.530 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 88.125 72.530 88.445 ;
      LAYER met4 ;
        RECT 72.210 88.125 72.530 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 87.715 72.530 88.035 ;
      LAYER met4 ;
        RECT 72.210 87.715 72.530 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 87.305 72.530 87.625 ;
      LAYER met4 ;
        RECT 72.210 87.305 72.530 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 86.895 72.530 87.215 ;
      LAYER met4 ;
        RECT 72.210 86.895 72.530 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 86.485 72.530 86.805 ;
      LAYER met4 ;
        RECT 72.210 86.485 72.530 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 86.075 72.530 86.395 ;
      LAYER met4 ;
        RECT 72.210 86.075 72.530 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 85.665 72.530 85.985 ;
      LAYER met4 ;
        RECT 72.210 85.665 72.530 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 85.255 72.530 85.575 ;
      LAYER met4 ;
        RECT 72.210 85.255 72.530 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 84.845 72.530 85.165 ;
      LAYER met4 ;
        RECT 72.210 84.845 72.530 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 84.435 72.530 84.755 ;
      LAYER met4 ;
        RECT 72.210 84.435 72.530 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 84.025 72.530 84.345 ;
      LAYER met4 ;
        RECT 72.210 84.025 72.530 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 83.615 72.530 83.935 ;
      LAYER met4 ;
        RECT 72.210 83.615 72.530 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 83.205 72.530 83.525 ;
      LAYER met4 ;
        RECT 72.210 83.205 72.530 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 82.795 72.530 83.115 ;
      LAYER met4 ;
        RECT 72.210 82.795 72.530 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 82.360 72.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 81.955 72.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 81.550 72.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 81.145 72.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 80.740 72.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 80.335 72.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 79.930 72.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 79.525 72.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 79.120 72.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 78.715 72.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 78.310 72.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 77.905 72.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 77.500 72.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 77.095 72.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 76.690 72.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 76.285 72.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 75.880 72.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 75.475 72.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 75.070 72.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 74.665 72.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 74.260 72.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 73.855 72.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 73.450 72.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 73.045 72.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 72.635 72.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 72.225 72.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 71.815 72.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 71.405 72.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 70.995 72.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 70.585 72.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 70.175 72.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 69.765 72.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 69.355 72.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 68.945 72.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 68.535 72.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.210 68.125 72.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 22.160 72.105 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 21.730 72.105 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 21.300 72.105 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 20.870 72.105 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 20.440 72.105 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 20.010 72.105 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 19.580 72.105 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 19.150 72.105 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 18.720 72.105 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 18.290 72.105 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.905 17.860 72.105 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.860 92.695 72.060 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 92.225 72.120 92.545 ;
      LAYER met4 ;
        RECT 71.800 92.225 72.120 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 91.815 72.120 92.135 ;
      LAYER met4 ;
        RECT 71.800 91.815 72.120 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 91.405 72.120 91.725 ;
      LAYER met4 ;
        RECT 71.800 91.405 72.120 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 90.995 72.120 91.315 ;
      LAYER met4 ;
        RECT 71.800 90.995 72.120 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 90.585 72.120 90.905 ;
      LAYER met4 ;
        RECT 71.800 90.585 72.120 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 90.175 72.120 90.495 ;
      LAYER met4 ;
        RECT 71.800 90.175 72.120 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 89.765 72.120 90.085 ;
      LAYER met4 ;
        RECT 71.800 89.765 72.120 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 89.355 72.120 89.675 ;
      LAYER met4 ;
        RECT 71.800 89.355 72.120 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 88.945 72.120 89.265 ;
      LAYER met4 ;
        RECT 71.800 88.945 72.120 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 88.535 72.120 88.855 ;
      LAYER met4 ;
        RECT 71.800 88.535 72.120 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 88.125 72.120 88.445 ;
      LAYER met4 ;
        RECT 71.800 88.125 72.120 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 87.715 72.120 88.035 ;
      LAYER met4 ;
        RECT 71.800 87.715 72.120 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 87.305 72.120 87.625 ;
      LAYER met4 ;
        RECT 71.800 87.305 72.120 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 86.895 72.120 87.215 ;
      LAYER met4 ;
        RECT 71.800 86.895 72.120 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 86.485 72.120 86.805 ;
      LAYER met4 ;
        RECT 71.800 86.485 72.120 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 86.075 72.120 86.395 ;
      LAYER met4 ;
        RECT 71.800 86.075 72.120 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 85.665 72.120 85.985 ;
      LAYER met4 ;
        RECT 71.800 85.665 72.120 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 85.255 72.120 85.575 ;
      LAYER met4 ;
        RECT 71.800 85.255 72.120 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 84.845 72.120 85.165 ;
      LAYER met4 ;
        RECT 71.800 84.845 72.120 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 84.435 72.120 84.755 ;
      LAYER met4 ;
        RECT 71.800 84.435 72.120 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 84.025 72.120 84.345 ;
      LAYER met4 ;
        RECT 71.800 84.025 72.120 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 83.615 72.120 83.935 ;
      LAYER met4 ;
        RECT 71.800 83.615 72.120 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 83.205 72.120 83.525 ;
      LAYER met4 ;
        RECT 71.800 83.205 72.120 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.800 82.795 72.120 83.115 ;
      LAYER met4 ;
        RECT 71.800 82.795 72.120 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 82.360 72.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 81.955 72.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 81.550 72.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 81.145 72.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 80.740 72.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 80.335 72.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 79.930 72.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 79.525 72.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 79.120 72.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 78.715 72.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 78.310 72.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 77.905 72.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 77.500 72.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 77.095 72.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 76.690 72.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 76.285 72.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 75.880 72.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 75.475 72.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 75.070 72.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 74.665 72.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 74.260 72.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 73.855 72.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 73.450 72.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 73.045 72.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 72.635 72.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 72.225 72.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 71.815 72.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 71.405 72.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 70.995 72.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 70.585 72.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 70.175 72.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 69.765 72.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 69.355 72.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 68.945 72.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 68.535 72.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.810 68.125 72.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 22.160 71.700 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 21.730 71.700 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 21.300 71.700 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 20.870 71.700 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 20.440 71.700 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 20.010 71.700 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 19.580 71.700 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 19.150 71.700 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 18.720 71.700 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 18.290 71.700 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.500 17.860 71.700 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.450 92.695 71.650 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 92.225 71.710 92.545 ;
      LAYER met4 ;
        RECT 71.390 92.225 71.710 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 91.815 71.710 92.135 ;
      LAYER met4 ;
        RECT 71.390 91.815 71.710 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 91.405 71.710 91.725 ;
      LAYER met4 ;
        RECT 71.390 91.405 71.710 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 90.995 71.710 91.315 ;
      LAYER met4 ;
        RECT 71.390 90.995 71.710 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 90.585 71.710 90.905 ;
      LAYER met4 ;
        RECT 71.390 90.585 71.710 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 90.175 71.710 90.495 ;
      LAYER met4 ;
        RECT 71.390 90.175 71.710 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 89.765 71.710 90.085 ;
      LAYER met4 ;
        RECT 71.390 89.765 71.710 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 89.355 71.710 89.675 ;
      LAYER met4 ;
        RECT 71.390 89.355 71.710 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 88.945 71.710 89.265 ;
      LAYER met4 ;
        RECT 71.390 88.945 71.710 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 88.535 71.710 88.855 ;
      LAYER met4 ;
        RECT 71.390 88.535 71.710 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 88.125 71.710 88.445 ;
      LAYER met4 ;
        RECT 71.390 88.125 71.710 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 87.715 71.710 88.035 ;
      LAYER met4 ;
        RECT 71.390 87.715 71.710 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 87.305 71.710 87.625 ;
      LAYER met4 ;
        RECT 71.390 87.305 71.710 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 86.895 71.710 87.215 ;
      LAYER met4 ;
        RECT 71.390 86.895 71.710 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 86.485 71.710 86.805 ;
      LAYER met4 ;
        RECT 71.390 86.485 71.710 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 86.075 71.710 86.395 ;
      LAYER met4 ;
        RECT 71.390 86.075 71.710 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 85.665 71.710 85.985 ;
      LAYER met4 ;
        RECT 71.390 85.665 71.710 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 85.255 71.710 85.575 ;
      LAYER met4 ;
        RECT 71.390 85.255 71.710 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 84.845 71.710 85.165 ;
      LAYER met4 ;
        RECT 71.390 84.845 71.710 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 84.435 71.710 84.755 ;
      LAYER met4 ;
        RECT 71.390 84.435 71.710 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 84.025 71.710 84.345 ;
      LAYER met4 ;
        RECT 71.390 84.025 71.710 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 83.615 71.710 83.935 ;
      LAYER met4 ;
        RECT 71.390 83.615 71.710 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 83.205 71.710 83.525 ;
      LAYER met4 ;
        RECT 71.390 83.205 71.710 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.390 82.795 71.710 83.115 ;
      LAYER met4 ;
        RECT 71.390 82.795 71.710 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 82.360 71.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 81.955 71.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 81.550 71.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 81.145 71.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 80.740 71.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 80.335 71.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 79.930 71.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 79.525 71.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 79.120 71.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 78.715 71.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 78.310 71.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 77.905 71.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 77.500 71.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 77.095 71.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 76.690 71.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 76.285 71.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 75.880 71.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 75.475 71.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 75.070 71.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 74.665 71.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 74.260 71.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 73.855 71.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 73.450 71.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 73.045 71.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 72.635 71.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 72.225 71.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 71.815 71.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 71.405 71.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 70.995 71.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 70.585 71.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 70.175 71.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 69.765 71.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 69.355 71.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 68.945 71.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 68.535 71.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.410 68.125 71.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 22.160 71.295 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 21.730 71.295 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 21.300 71.295 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 20.870 71.295 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 20.440 71.295 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 20.010 71.295 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 19.580 71.295 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 19.150 71.295 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 18.720 71.295 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 18.290 71.295 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.095 17.860 71.295 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.040 92.695 71.240 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 92.225 71.300 92.545 ;
      LAYER met4 ;
        RECT 70.980 92.225 71.300 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 91.815 71.300 92.135 ;
      LAYER met4 ;
        RECT 70.980 91.815 71.300 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 91.405 71.300 91.725 ;
      LAYER met4 ;
        RECT 70.980 91.405 71.300 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 90.995 71.300 91.315 ;
      LAYER met4 ;
        RECT 70.980 90.995 71.300 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 90.585 71.300 90.905 ;
      LAYER met4 ;
        RECT 70.980 90.585 71.300 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 90.175 71.300 90.495 ;
      LAYER met4 ;
        RECT 70.980 90.175 71.300 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 89.765 71.300 90.085 ;
      LAYER met4 ;
        RECT 70.980 89.765 71.300 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 89.355 71.300 89.675 ;
      LAYER met4 ;
        RECT 70.980 89.355 71.300 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 88.945 71.300 89.265 ;
      LAYER met4 ;
        RECT 70.980 88.945 71.300 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 88.535 71.300 88.855 ;
      LAYER met4 ;
        RECT 70.980 88.535 71.300 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 88.125 71.300 88.445 ;
      LAYER met4 ;
        RECT 70.980 88.125 71.300 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 87.715 71.300 88.035 ;
      LAYER met4 ;
        RECT 70.980 87.715 71.300 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 87.305 71.300 87.625 ;
      LAYER met4 ;
        RECT 70.980 87.305 71.300 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 86.895 71.300 87.215 ;
      LAYER met4 ;
        RECT 70.980 86.895 71.300 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 86.485 71.300 86.805 ;
      LAYER met4 ;
        RECT 70.980 86.485 71.300 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 86.075 71.300 86.395 ;
      LAYER met4 ;
        RECT 70.980 86.075 71.300 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 85.665 71.300 85.985 ;
      LAYER met4 ;
        RECT 70.980 85.665 71.300 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 85.255 71.300 85.575 ;
      LAYER met4 ;
        RECT 70.980 85.255 71.300 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 84.845 71.300 85.165 ;
      LAYER met4 ;
        RECT 70.980 84.845 71.300 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 84.435 71.300 84.755 ;
      LAYER met4 ;
        RECT 70.980 84.435 71.300 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 84.025 71.300 84.345 ;
      LAYER met4 ;
        RECT 70.980 84.025 71.300 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 83.615 71.300 83.935 ;
      LAYER met4 ;
        RECT 70.980 83.615 71.300 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 83.205 71.300 83.525 ;
      LAYER met4 ;
        RECT 70.980 83.205 71.300 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.980 82.795 71.300 83.115 ;
      LAYER met4 ;
        RECT 70.980 82.795 71.300 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 82.360 71.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 81.955 71.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 81.550 71.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 81.145 71.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 80.740 71.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 80.335 71.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 79.930 71.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 79.525 71.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 79.120 71.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 78.715 71.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 78.310 71.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 77.905 71.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 77.500 71.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 77.095 71.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 76.690 71.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 76.285 71.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 75.880 71.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 75.475 71.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 75.070 71.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 74.665 71.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 74.260 71.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 73.855 71.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 73.450 71.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 73.045 71.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 72.635 71.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 72.225 71.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 71.815 71.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 71.405 71.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 70.995 71.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 70.585 71.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 70.175 71.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 69.765 71.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 69.355 71.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 68.945 71.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 68.535 71.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.010 68.125 71.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 22.160 70.890 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 21.730 70.890 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 21.300 70.890 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 20.870 70.890 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 20.440 70.890 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 20.010 70.890 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 19.580 70.890 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 19.150 70.890 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 18.720 70.890 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 18.290 70.890 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.690 17.860 70.890 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.630 92.695 70.830 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 92.225 70.890 92.545 ;
      LAYER met4 ;
        RECT 70.570 92.225 70.890 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 91.815 70.890 92.135 ;
      LAYER met4 ;
        RECT 70.570 91.815 70.890 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 91.405 70.890 91.725 ;
      LAYER met4 ;
        RECT 70.570 91.405 70.890 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 90.995 70.890 91.315 ;
      LAYER met4 ;
        RECT 70.570 90.995 70.890 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 90.585 70.890 90.905 ;
      LAYER met4 ;
        RECT 70.570 90.585 70.890 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 90.175 70.890 90.495 ;
      LAYER met4 ;
        RECT 70.570 90.175 70.890 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 89.765 70.890 90.085 ;
      LAYER met4 ;
        RECT 70.570 89.765 70.890 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 89.355 70.890 89.675 ;
      LAYER met4 ;
        RECT 70.570 89.355 70.890 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 88.945 70.890 89.265 ;
      LAYER met4 ;
        RECT 70.570 88.945 70.890 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 88.535 70.890 88.855 ;
      LAYER met4 ;
        RECT 70.570 88.535 70.890 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 88.125 70.890 88.445 ;
      LAYER met4 ;
        RECT 70.570 88.125 70.890 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 87.715 70.890 88.035 ;
      LAYER met4 ;
        RECT 70.570 87.715 70.890 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 87.305 70.890 87.625 ;
      LAYER met4 ;
        RECT 70.570 87.305 70.890 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 86.895 70.890 87.215 ;
      LAYER met4 ;
        RECT 70.570 86.895 70.890 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 86.485 70.890 86.805 ;
      LAYER met4 ;
        RECT 70.570 86.485 70.890 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 86.075 70.890 86.395 ;
      LAYER met4 ;
        RECT 70.570 86.075 70.890 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 85.665 70.890 85.985 ;
      LAYER met4 ;
        RECT 70.570 85.665 70.890 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 85.255 70.890 85.575 ;
      LAYER met4 ;
        RECT 70.570 85.255 70.890 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 84.845 70.890 85.165 ;
      LAYER met4 ;
        RECT 70.570 84.845 70.890 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 84.435 70.890 84.755 ;
      LAYER met4 ;
        RECT 70.570 84.435 70.890 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 84.025 70.890 84.345 ;
      LAYER met4 ;
        RECT 70.570 84.025 70.890 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 83.615 70.890 83.935 ;
      LAYER met4 ;
        RECT 70.570 83.615 70.890 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 83.205 70.890 83.525 ;
      LAYER met4 ;
        RECT 70.570 83.205 70.890 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.570 82.795 70.890 83.115 ;
      LAYER met4 ;
        RECT 70.570 82.795 70.890 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 82.360 70.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 81.955 70.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 81.550 70.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 81.145 70.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 80.740 70.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 80.335 70.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 79.930 70.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 79.525 70.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 79.120 70.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 78.715 70.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 78.310 70.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 77.905 70.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 77.500 70.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 77.095 70.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 76.690 70.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 76.285 70.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 75.880 70.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 75.475 70.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 75.070 70.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 74.665 70.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 74.260 70.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 73.855 70.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 73.450 70.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 73.045 70.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 72.635 70.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 72.225 70.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 71.815 70.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 71.405 70.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 70.995 70.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 70.585 70.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 70.175 70.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 69.765 70.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 69.355 70.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 68.945 70.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 68.535 70.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.610 68.125 70.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 22.160 70.485 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 21.730 70.485 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 21.300 70.485 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 20.870 70.485 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 20.440 70.485 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 20.010 70.485 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 19.580 70.485 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 19.150 70.485 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 18.720 70.485 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 18.290 70.485 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.285 17.860 70.485 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.220 92.695 70.420 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 92.225 70.480 92.545 ;
      LAYER met4 ;
        RECT 70.160 92.225 70.480 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 91.815 70.480 92.135 ;
      LAYER met4 ;
        RECT 70.160 91.815 70.480 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 91.405 70.480 91.725 ;
      LAYER met4 ;
        RECT 70.160 91.405 70.480 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 90.995 70.480 91.315 ;
      LAYER met4 ;
        RECT 70.160 90.995 70.480 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 90.585 70.480 90.905 ;
      LAYER met4 ;
        RECT 70.160 90.585 70.480 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 90.175 70.480 90.495 ;
      LAYER met4 ;
        RECT 70.160 90.175 70.480 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 89.765 70.480 90.085 ;
      LAYER met4 ;
        RECT 70.160 89.765 70.480 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 89.355 70.480 89.675 ;
      LAYER met4 ;
        RECT 70.160 89.355 70.480 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 88.945 70.480 89.265 ;
      LAYER met4 ;
        RECT 70.160 88.945 70.480 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 88.535 70.480 88.855 ;
      LAYER met4 ;
        RECT 70.160 88.535 70.480 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 88.125 70.480 88.445 ;
      LAYER met4 ;
        RECT 70.160 88.125 70.480 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 87.715 70.480 88.035 ;
      LAYER met4 ;
        RECT 70.160 87.715 70.480 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 87.305 70.480 87.625 ;
      LAYER met4 ;
        RECT 70.160 87.305 70.480 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 86.895 70.480 87.215 ;
      LAYER met4 ;
        RECT 70.160 86.895 70.480 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 86.485 70.480 86.805 ;
      LAYER met4 ;
        RECT 70.160 86.485 70.480 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 86.075 70.480 86.395 ;
      LAYER met4 ;
        RECT 70.160 86.075 70.480 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 85.665 70.480 85.985 ;
      LAYER met4 ;
        RECT 70.160 85.665 70.480 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 85.255 70.480 85.575 ;
      LAYER met4 ;
        RECT 70.160 85.255 70.480 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 84.845 70.480 85.165 ;
      LAYER met4 ;
        RECT 70.160 84.845 70.480 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 84.435 70.480 84.755 ;
      LAYER met4 ;
        RECT 70.160 84.435 70.480 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 84.025 70.480 84.345 ;
      LAYER met4 ;
        RECT 70.160 84.025 70.480 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 83.615 70.480 83.935 ;
      LAYER met4 ;
        RECT 70.160 83.615 70.480 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 83.205 70.480 83.525 ;
      LAYER met4 ;
        RECT 70.160 83.205 70.480 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.160 82.795 70.480 83.115 ;
      LAYER met4 ;
        RECT 70.160 82.795 70.480 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 82.360 70.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 81.955 70.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 81.550 70.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 81.145 70.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 80.740 70.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 80.335 70.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 79.930 70.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 79.525 70.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 79.120 70.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 78.715 70.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 78.310 70.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 77.905 70.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 77.500 70.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 77.095 70.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 76.690 70.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 76.285 70.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 75.880 70.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 75.475 70.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 75.070 70.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 74.665 70.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 74.260 70.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 73.855 70.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 73.450 70.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 73.045 70.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 72.635 70.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 72.225 70.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 71.815 70.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 71.405 70.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 70.995 70.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 70.585 70.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 70.175 70.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 69.765 70.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 69.355 70.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 68.945 70.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 68.535 70.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.210 68.125 70.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 22.160 70.080 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 21.730 70.080 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 21.300 70.080 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 20.870 70.080 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 20.440 70.080 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 20.010 70.080 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 19.580 70.080 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 19.150 70.080 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 18.720 70.080 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 18.290 70.080 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.880 17.860 70.080 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 92.695 70.010 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 92.225 70.070 92.545 ;
      LAYER met4 ;
        RECT 69.750 92.225 70.070 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 91.815 70.070 92.135 ;
      LAYER met4 ;
        RECT 69.750 91.815 70.070 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 91.405 70.070 91.725 ;
      LAYER met4 ;
        RECT 69.750 91.405 70.070 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 90.995 70.070 91.315 ;
      LAYER met4 ;
        RECT 69.750 90.995 70.070 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 90.585 70.070 90.905 ;
      LAYER met4 ;
        RECT 69.750 90.585 70.070 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 90.175 70.070 90.495 ;
      LAYER met4 ;
        RECT 69.750 90.175 70.070 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 89.765 70.070 90.085 ;
      LAYER met4 ;
        RECT 69.750 89.765 70.070 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 89.355 70.070 89.675 ;
      LAYER met4 ;
        RECT 69.750 89.355 70.070 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 88.945 70.070 89.265 ;
      LAYER met4 ;
        RECT 69.750 88.945 70.070 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 88.535 70.070 88.855 ;
      LAYER met4 ;
        RECT 69.750 88.535 70.070 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 88.125 70.070 88.445 ;
      LAYER met4 ;
        RECT 69.750 88.125 70.070 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 87.715 70.070 88.035 ;
      LAYER met4 ;
        RECT 69.750 87.715 70.070 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 87.305 70.070 87.625 ;
      LAYER met4 ;
        RECT 69.750 87.305 70.070 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 86.895 70.070 87.215 ;
      LAYER met4 ;
        RECT 69.750 86.895 70.070 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 86.485 70.070 86.805 ;
      LAYER met4 ;
        RECT 69.750 86.485 70.070 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 86.075 70.070 86.395 ;
      LAYER met4 ;
        RECT 69.750 86.075 70.070 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 85.665 70.070 85.985 ;
      LAYER met4 ;
        RECT 69.750 85.665 70.070 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 85.255 70.070 85.575 ;
      LAYER met4 ;
        RECT 69.750 85.255 70.070 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 84.845 70.070 85.165 ;
      LAYER met4 ;
        RECT 69.750 84.845 70.070 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 84.435 70.070 84.755 ;
      LAYER met4 ;
        RECT 69.750 84.435 70.070 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 84.025 70.070 84.345 ;
      LAYER met4 ;
        RECT 69.750 84.025 70.070 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 83.615 70.070 83.935 ;
      LAYER met4 ;
        RECT 69.750 83.615 70.070 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 83.205 70.070 83.525 ;
      LAYER met4 ;
        RECT 69.750 83.205 70.070 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.750 82.795 70.070 83.115 ;
      LAYER met4 ;
        RECT 69.750 82.795 70.070 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 82.360 70.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 81.955 70.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 81.550 70.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 81.145 70.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 80.740 70.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 80.335 70.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 79.930 70.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 79.525 70.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 79.120 70.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 78.715 70.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 78.310 70.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 77.905 70.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 77.500 70.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 77.095 70.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 76.690 70.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 76.285 70.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 75.880 70.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 75.475 70.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 75.070 70.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 74.665 70.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 74.260 70.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 73.855 70.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 73.450 70.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 73.045 70.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 72.635 70.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 72.225 70.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 71.815 70.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 71.405 70.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 70.995 70.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 70.585 70.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 70.175 70.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 69.765 70.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 69.355 70.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 68.945 70.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 68.535 70.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.810 68.125 70.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 22.160 69.675 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 21.730 69.675 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 21.300 69.675 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 20.870 69.675 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 20.440 69.675 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 20.010 69.675 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 19.580 69.675 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 19.150 69.675 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 18.720 69.675 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 18.290 69.675 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.475 17.860 69.675 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 82.360 69.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 81.955 69.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 81.550 69.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 81.145 69.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 80.740 69.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 80.335 69.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 79.930 69.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 79.525 69.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 79.120 69.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 78.715 69.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 78.310 69.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 77.905 69.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 77.500 69.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 77.095 69.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 76.690 69.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 76.285 69.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 75.880 69.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 75.475 69.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 75.070 69.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 74.665 69.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 74.260 69.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 73.855 69.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 73.450 69.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 73.045 69.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 72.635 69.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 72.225 69.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 71.815 69.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 71.405 69.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 70.995 69.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 70.585 69.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 70.175 69.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 69.765 69.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 69.355 69.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 68.945 69.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 68.535 69.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.410 68.125 69.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.400 92.695 69.600 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 92.225 69.660 92.545 ;
      LAYER met4 ;
        RECT 69.340 92.225 69.660 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 91.815 69.660 92.135 ;
      LAYER met4 ;
        RECT 69.340 91.815 69.660 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 91.405 69.660 91.725 ;
      LAYER met4 ;
        RECT 69.340 91.405 69.660 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 90.995 69.660 91.315 ;
      LAYER met4 ;
        RECT 69.340 90.995 69.660 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 90.585 69.660 90.905 ;
      LAYER met4 ;
        RECT 69.340 90.585 69.660 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 90.175 69.660 90.495 ;
      LAYER met4 ;
        RECT 69.340 90.175 69.660 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 89.765 69.660 90.085 ;
      LAYER met4 ;
        RECT 69.340 89.765 69.660 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 89.355 69.660 89.675 ;
      LAYER met4 ;
        RECT 69.340 89.355 69.660 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 88.945 69.660 89.265 ;
      LAYER met4 ;
        RECT 69.340 88.945 69.660 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 88.535 69.660 88.855 ;
      LAYER met4 ;
        RECT 69.340 88.535 69.660 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 88.125 69.660 88.445 ;
      LAYER met4 ;
        RECT 69.340 88.125 69.660 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 87.715 69.660 88.035 ;
      LAYER met4 ;
        RECT 69.340 87.715 69.660 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 87.305 69.660 87.625 ;
      LAYER met4 ;
        RECT 69.340 87.305 69.660 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 86.895 69.660 87.215 ;
      LAYER met4 ;
        RECT 69.340 86.895 69.660 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 86.485 69.660 86.805 ;
      LAYER met4 ;
        RECT 69.340 86.485 69.660 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 86.075 69.660 86.395 ;
      LAYER met4 ;
        RECT 69.340 86.075 69.660 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 85.665 69.660 85.985 ;
      LAYER met4 ;
        RECT 69.340 85.665 69.660 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 85.255 69.660 85.575 ;
      LAYER met4 ;
        RECT 69.340 85.255 69.660 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 84.845 69.660 85.165 ;
      LAYER met4 ;
        RECT 69.340 84.845 69.660 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 84.435 69.660 84.755 ;
      LAYER met4 ;
        RECT 69.340 84.435 69.660 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 84.025 69.660 84.345 ;
      LAYER met4 ;
        RECT 69.340 84.025 69.660 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 83.615 69.660 83.935 ;
      LAYER met4 ;
        RECT 69.340 83.615 69.660 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 83.205 69.660 83.525 ;
      LAYER met4 ;
        RECT 69.340 83.205 69.660 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.340 82.795 69.660 83.115 ;
      LAYER met4 ;
        RECT 69.340 82.795 69.660 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 22.160 69.270 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 21.730 69.270 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 21.300 69.270 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 20.870 69.270 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 20.440 69.270 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 20.010 69.270 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 19.580 69.270 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 19.150 69.270 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 18.720 69.270 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 18.290 69.270 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.070 17.860 69.270 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 82.360 69.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 81.955 69.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 81.550 69.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 81.145 69.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 80.740 69.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 80.335 69.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 79.930 69.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 79.525 69.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 79.120 69.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 78.715 69.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 78.310 69.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 77.905 69.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 77.500 69.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 77.095 69.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 76.690 69.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 76.285 69.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 75.880 69.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 75.475 69.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 75.070 69.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 74.665 69.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 74.260 69.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 73.855 69.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 73.450 69.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 73.045 69.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 72.635 69.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 72.225 69.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 71.815 69.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 71.405 69.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 70.995 69.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 70.585 69.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 70.175 69.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 69.765 69.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 69.355 69.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 68.945 69.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 68.535 69.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.010 68.125 69.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.990 92.695 69.190 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 92.225 69.250 92.545 ;
      LAYER met4 ;
        RECT 68.930 92.225 69.250 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 91.815 69.250 92.135 ;
      LAYER met4 ;
        RECT 68.930 91.815 69.250 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 91.405 69.250 91.725 ;
      LAYER met4 ;
        RECT 68.930 91.405 69.250 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 90.995 69.250 91.315 ;
      LAYER met4 ;
        RECT 68.930 90.995 69.250 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 90.585 69.250 90.905 ;
      LAYER met4 ;
        RECT 68.930 90.585 69.250 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 90.175 69.250 90.495 ;
      LAYER met4 ;
        RECT 68.930 90.175 69.250 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 89.765 69.250 90.085 ;
      LAYER met4 ;
        RECT 68.930 89.765 69.250 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 89.355 69.250 89.675 ;
      LAYER met4 ;
        RECT 68.930 89.355 69.250 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 88.945 69.250 89.265 ;
      LAYER met4 ;
        RECT 68.930 88.945 69.250 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 88.535 69.250 88.855 ;
      LAYER met4 ;
        RECT 68.930 88.535 69.250 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 88.125 69.250 88.445 ;
      LAYER met4 ;
        RECT 68.930 88.125 69.250 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 87.715 69.250 88.035 ;
      LAYER met4 ;
        RECT 68.930 87.715 69.250 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 87.305 69.250 87.625 ;
      LAYER met4 ;
        RECT 68.930 87.305 69.250 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 86.895 69.250 87.215 ;
      LAYER met4 ;
        RECT 68.930 86.895 69.250 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 86.485 69.250 86.805 ;
      LAYER met4 ;
        RECT 68.930 86.485 69.250 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 86.075 69.250 86.395 ;
      LAYER met4 ;
        RECT 68.930 86.075 69.250 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 85.665 69.250 85.985 ;
      LAYER met4 ;
        RECT 68.930 85.665 69.250 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 85.255 69.250 85.575 ;
      LAYER met4 ;
        RECT 68.930 85.255 69.250 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 84.845 69.250 85.165 ;
      LAYER met4 ;
        RECT 68.930 84.845 69.250 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 84.435 69.250 84.755 ;
      LAYER met4 ;
        RECT 68.930 84.435 69.250 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 84.025 69.250 84.345 ;
      LAYER met4 ;
        RECT 68.930 84.025 69.250 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 83.615 69.250 83.935 ;
      LAYER met4 ;
        RECT 68.930 83.615 69.250 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 83.205 69.250 83.525 ;
      LAYER met4 ;
        RECT 68.930 83.205 69.250 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.930 82.795 69.250 83.115 ;
      LAYER met4 ;
        RECT 68.930 82.795 69.250 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 22.160 68.865 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 21.730 68.865 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 21.300 68.865 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 20.870 68.865 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 20.440 68.865 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 20.010 68.865 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 19.580 68.865 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 19.150 68.865 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 18.720 68.865 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 18.290 68.865 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.665 17.860 68.865 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 82.360 68.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 81.955 68.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 81.550 68.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 81.145 68.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 80.740 68.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 80.335 68.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 79.930 68.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 79.525 68.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 79.120 68.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 78.715 68.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 78.310 68.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 77.905 68.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 77.500 68.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 77.095 68.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 76.690 68.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 76.285 68.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 75.880 68.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 75.475 68.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 75.070 68.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 74.665 68.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 74.260 68.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 73.855 68.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 73.450 68.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 73.045 68.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 72.635 68.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 72.225 68.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 71.815 68.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 71.405 68.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 70.995 68.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 70.585 68.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 70.175 68.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 69.765 68.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 69.355 68.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 68.945 68.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 68.535 68.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.610 68.125 68.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.580 92.695 68.780 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 92.225 68.840 92.545 ;
      LAYER met4 ;
        RECT 68.520 92.225 68.840 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 91.815 68.840 92.135 ;
      LAYER met4 ;
        RECT 68.520 91.815 68.840 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 91.405 68.840 91.725 ;
      LAYER met4 ;
        RECT 68.520 91.405 68.840 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 90.995 68.840 91.315 ;
      LAYER met4 ;
        RECT 68.520 90.995 68.840 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 90.585 68.840 90.905 ;
      LAYER met4 ;
        RECT 68.520 90.585 68.840 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 90.175 68.840 90.495 ;
      LAYER met4 ;
        RECT 68.520 90.175 68.840 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 89.765 68.840 90.085 ;
      LAYER met4 ;
        RECT 68.520 89.765 68.840 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 89.355 68.840 89.675 ;
      LAYER met4 ;
        RECT 68.520 89.355 68.840 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 88.945 68.840 89.265 ;
      LAYER met4 ;
        RECT 68.520 88.945 68.840 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 88.535 68.840 88.855 ;
      LAYER met4 ;
        RECT 68.520 88.535 68.840 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 88.125 68.840 88.445 ;
      LAYER met4 ;
        RECT 68.520 88.125 68.840 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 87.715 68.840 88.035 ;
      LAYER met4 ;
        RECT 68.520 87.715 68.840 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 87.305 68.840 87.625 ;
      LAYER met4 ;
        RECT 68.520 87.305 68.840 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 86.895 68.840 87.215 ;
      LAYER met4 ;
        RECT 68.520 86.895 68.840 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 86.485 68.840 86.805 ;
      LAYER met4 ;
        RECT 68.520 86.485 68.840 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 86.075 68.840 86.395 ;
      LAYER met4 ;
        RECT 68.520 86.075 68.840 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 85.665 68.840 85.985 ;
      LAYER met4 ;
        RECT 68.520 85.665 68.840 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 85.255 68.840 85.575 ;
      LAYER met4 ;
        RECT 68.520 85.255 68.840 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 84.845 68.840 85.165 ;
      LAYER met4 ;
        RECT 68.520 84.845 68.840 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 84.435 68.840 84.755 ;
      LAYER met4 ;
        RECT 68.520 84.435 68.840 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 84.025 68.840 84.345 ;
      LAYER met4 ;
        RECT 68.520 84.025 68.840 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 83.615 68.840 83.935 ;
      LAYER met4 ;
        RECT 68.520 83.615 68.840 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 83.205 68.840 83.525 ;
      LAYER met4 ;
        RECT 68.520 83.205 68.840 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.520 82.795 68.840 83.115 ;
      LAYER met4 ;
        RECT 68.520 82.795 68.840 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 22.160 68.460 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 21.730 68.460 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 21.300 68.460 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 20.870 68.460 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 20.440 68.460 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 20.010 68.460 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 19.580 68.460 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 19.150 68.460 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 18.720 68.460 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 18.290 68.460 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.260 17.860 68.460 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 82.360 68.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 81.955 68.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 81.550 68.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 81.145 68.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 80.740 68.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 80.335 68.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 79.930 68.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 79.525 68.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 79.120 68.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 78.715 68.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 78.310 68.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 77.905 68.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 77.500 68.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 77.095 68.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 76.690 68.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 76.285 68.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 75.880 68.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 75.475 68.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 75.070 68.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 74.665 68.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 74.260 68.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 73.855 68.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 73.450 68.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 73.045 68.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 72.635 68.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 72.225 68.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 71.815 68.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 71.405 68.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 70.995 68.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 70.585 68.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 70.175 68.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 69.765 68.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 69.355 68.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 68.945 68.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 68.535 68.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.210 68.125 68.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.170 92.695 68.370 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 92.225 68.430 92.545 ;
      LAYER met4 ;
        RECT 68.110 92.225 68.430 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 91.815 68.430 92.135 ;
      LAYER met4 ;
        RECT 68.110 91.815 68.430 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 91.405 68.430 91.725 ;
      LAYER met4 ;
        RECT 68.110 91.405 68.430 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 90.995 68.430 91.315 ;
      LAYER met4 ;
        RECT 68.110 90.995 68.430 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 90.585 68.430 90.905 ;
      LAYER met4 ;
        RECT 68.110 90.585 68.430 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 90.175 68.430 90.495 ;
      LAYER met4 ;
        RECT 68.110 90.175 68.430 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 89.765 68.430 90.085 ;
      LAYER met4 ;
        RECT 68.110 89.765 68.430 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 89.355 68.430 89.675 ;
      LAYER met4 ;
        RECT 68.110 89.355 68.430 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 88.945 68.430 89.265 ;
      LAYER met4 ;
        RECT 68.110 88.945 68.430 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 88.535 68.430 88.855 ;
      LAYER met4 ;
        RECT 68.110 88.535 68.430 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 88.125 68.430 88.445 ;
      LAYER met4 ;
        RECT 68.110 88.125 68.430 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 87.715 68.430 88.035 ;
      LAYER met4 ;
        RECT 68.110 87.715 68.430 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 87.305 68.430 87.625 ;
      LAYER met4 ;
        RECT 68.110 87.305 68.430 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 86.895 68.430 87.215 ;
      LAYER met4 ;
        RECT 68.110 86.895 68.430 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 86.485 68.430 86.805 ;
      LAYER met4 ;
        RECT 68.110 86.485 68.430 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 86.075 68.430 86.395 ;
      LAYER met4 ;
        RECT 68.110 86.075 68.430 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 85.665 68.430 85.985 ;
      LAYER met4 ;
        RECT 68.110 85.665 68.430 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 85.255 68.430 85.575 ;
      LAYER met4 ;
        RECT 68.110 85.255 68.430 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 84.845 68.430 85.165 ;
      LAYER met4 ;
        RECT 68.110 84.845 68.430 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 84.435 68.430 84.755 ;
      LAYER met4 ;
        RECT 68.110 84.435 68.430 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 84.025 68.430 84.345 ;
      LAYER met4 ;
        RECT 68.110 84.025 68.430 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 83.615 68.430 83.935 ;
      LAYER met4 ;
        RECT 68.110 83.615 68.430 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 83.205 68.430 83.525 ;
      LAYER met4 ;
        RECT 68.110 83.205 68.430 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.110 82.795 68.430 83.115 ;
      LAYER met4 ;
        RECT 68.110 82.795 68.430 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 22.160 68.055 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 21.730 68.055 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 21.300 68.055 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 20.870 68.055 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 20.440 68.055 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 20.010 68.055 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 19.580 68.055 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 19.150 68.055 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 18.720 68.055 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 18.290 68.055 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.855 17.860 68.055 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 82.360 68.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 81.955 68.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 81.550 68.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 81.145 68.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 80.740 68.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 80.335 68.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 79.930 68.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 79.525 68.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 79.120 68.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 78.715 68.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 78.310 68.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 77.905 68.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 77.500 68.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 77.095 68.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 76.690 68.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 76.285 68.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 75.880 68.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 75.475 68.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 75.070 68.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 74.665 68.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 74.260 68.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 73.855 68.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 73.450 68.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 73.045 68.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 72.635 68.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 72.225 68.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 71.815 68.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 71.405 68.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 70.995 68.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 70.585 68.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 70.175 68.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 69.765 68.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 69.355 68.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 68.945 68.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 68.535 68.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 68.125 68.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.760 92.695 67.960 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 92.225 68.020 92.545 ;
      LAYER met4 ;
        RECT 67.700 92.225 68.020 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 91.815 68.020 92.135 ;
      LAYER met4 ;
        RECT 67.700 91.815 68.020 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 91.405 68.020 91.725 ;
      LAYER met4 ;
        RECT 67.700 91.405 68.020 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 90.995 68.020 91.315 ;
      LAYER met4 ;
        RECT 67.700 90.995 68.020 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 90.585 68.020 90.905 ;
      LAYER met4 ;
        RECT 67.700 90.585 68.020 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 90.175 68.020 90.495 ;
      LAYER met4 ;
        RECT 67.700 90.175 68.020 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 89.765 68.020 90.085 ;
      LAYER met4 ;
        RECT 67.700 89.765 68.020 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 89.355 68.020 89.675 ;
      LAYER met4 ;
        RECT 67.700 89.355 68.020 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 88.945 68.020 89.265 ;
      LAYER met4 ;
        RECT 67.700 88.945 68.020 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 88.535 68.020 88.855 ;
      LAYER met4 ;
        RECT 67.700 88.535 68.020 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 88.125 68.020 88.445 ;
      LAYER met4 ;
        RECT 67.700 88.125 68.020 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 87.715 68.020 88.035 ;
      LAYER met4 ;
        RECT 67.700 87.715 68.020 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 87.305 68.020 87.625 ;
      LAYER met4 ;
        RECT 67.700 87.305 68.020 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 86.895 68.020 87.215 ;
      LAYER met4 ;
        RECT 67.700 86.895 68.020 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 86.485 68.020 86.805 ;
      LAYER met4 ;
        RECT 67.700 86.485 68.020 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 86.075 68.020 86.395 ;
      LAYER met4 ;
        RECT 67.700 86.075 68.020 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 85.665 68.020 85.985 ;
      LAYER met4 ;
        RECT 67.700 85.665 68.020 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 85.255 68.020 85.575 ;
      LAYER met4 ;
        RECT 67.700 85.255 68.020 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 84.845 68.020 85.165 ;
      LAYER met4 ;
        RECT 67.700 84.845 68.020 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 84.435 68.020 84.755 ;
      LAYER met4 ;
        RECT 67.700 84.435 68.020 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 84.025 68.020 84.345 ;
      LAYER met4 ;
        RECT 67.700 84.025 68.020 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 83.615 68.020 83.935 ;
      LAYER met4 ;
        RECT 67.700 83.615 68.020 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 83.205 68.020 83.525 ;
      LAYER met4 ;
        RECT 67.700 83.205 68.020 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.700 82.795 68.020 83.115 ;
      LAYER met4 ;
        RECT 67.700 82.795 68.020 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 22.160 67.650 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 21.730 67.650 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 21.300 67.650 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 20.870 67.650 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 20.440 67.650 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 20.010 67.650 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 19.580 67.650 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 19.150 67.650 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 18.720 67.650 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 18.290 67.650 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.450 17.860 67.650 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 82.360 67.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 81.955 67.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 81.550 67.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 81.145 67.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 80.740 67.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 80.335 67.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 79.930 67.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 79.525 67.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 79.120 67.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 78.715 67.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 78.310 67.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 77.905 67.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 77.500 67.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 77.095 67.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 76.690 67.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 76.285 67.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 75.880 67.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 75.475 67.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 75.070 67.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 74.665 67.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 74.260 67.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 73.855 67.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 73.450 67.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 73.045 67.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 72.635 67.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 72.225 67.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 71.815 67.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 71.405 67.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 70.995 67.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 70.585 67.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 70.175 67.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 69.765 67.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 69.355 67.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 68.945 67.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 68.535 67.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.410 68.125 67.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.350 92.695 67.550 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 92.225 67.610 92.545 ;
      LAYER met4 ;
        RECT 67.290 92.225 67.610 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 91.815 67.610 92.135 ;
      LAYER met4 ;
        RECT 67.290 91.815 67.610 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 91.405 67.610 91.725 ;
      LAYER met4 ;
        RECT 67.290 91.405 67.610 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 90.995 67.610 91.315 ;
      LAYER met4 ;
        RECT 67.290 90.995 67.610 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 90.585 67.610 90.905 ;
      LAYER met4 ;
        RECT 67.290 90.585 67.610 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 90.175 67.610 90.495 ;
      LAYER met4 ;
        RECT 67.290 90.175 67.610 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 89.765 67.610 90.085 ;
      LAYER met4 ;
        RECT 67.290 89.765 67.610 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 89.355 67.610 89.675 ;
      LAYER met4 ;
        RECT 67.290 89.355 67.610 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 88.945 67.610 89.265 ;
      LAYER met4 ;
        RECT 67.290 88.945 67.610 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 88.535 67.610 88.855 ;
      LAYER met4 ;
        RECT 67.290 88.535 67.610 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 88.125 67.610 88.445 ;
      LAYER met4 ;
        RECT 67.290 88.125 67.610 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 87.715 67.610 88.035 ;
      LAYER met4 ;
        RECT 67.290 87.715 67.610 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 87.305 67.610 87.625 ;
      LAYER met4 ;
        RECT 67.290 87.305 67.610 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 86.895 67.610 87.215 ;
      LAYER met4 ;
        RECT 67.290 86.895 67.610 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 86.485 67.610 86.805 ;
      LAYER met4 ;
        RECT 67.290 86.485 67.610 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 86.075 67.610 86.395 ;
      LAYER met4 ;
        RECT 67.290 86.075 67.610 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 85.665 67.610 85.985 ;
      LAYER met4 ;
        RECT 67.290 85.665 67.610 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 85.255 67.610 85.575 ;
      LAYER met4 ;
        RECT 67.290 85.255 67.610 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 84.845 67.610 85.165 ;
      LAYER met4 ;
        RECT 67.290 84.845 67.610 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 84.435 67.610 84.755 ;
      LAYER met4 ;
        RECT 67.290 84.435 67.610 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 84.025 67.610 84.345 ;
      LAYER met4 ;
        RECT 67.290 84.025 67.610 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 83.615 67.610 83.935 ;
      LAYER met4 ;
        RECT 67.290 83.615 67.610 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 83.205 67.610 83.525 ;
      LAYER met4 ;
        RECT 67.290 83.205 67.610 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.290 82.795 67.610 83.115 ;
      LAYER met4 ;
        RECT 67.290 82.795 67.610 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 22.160 67.245 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 21.730 67.245 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 21.300 67.245 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 20.870 67.245 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 20.440 67.245 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 20.010 67.245 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 19.580 67.245 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 19.150 67.245 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 18.720 67.245 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 18.290 67.245 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.045 17.860 67.245 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 82.360 67.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 81.955 67.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 81.550 67.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 81.145 67.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 80.740 67.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 80.335 67.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 79.930 67.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 79.525 67.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 79.120 67.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 78.715 67.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 78.310 67.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 77.905 67.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 77.500 67.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 77.095 67.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 76.690 67.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 76.285 67.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 75.880 67.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 75.475 67.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 75.070 67.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 74.665 67.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 74.260 67.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 73.855 67.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 73.450 67.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 73.045 67.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 72.635 67.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 72.225 67.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 71.815 67.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 71.405 67.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 70.995 67.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 70.585 67.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 70.175 67.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 69.765 67.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 69.355 67.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 68.945 67.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 68.535 67.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.010 68.125 67.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.940 92.695 67.140 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 92.225 67.200 92.545 ;
      LAYER met4 ;
        RECT 66.880 92.225 67.200 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 91.815 67.200 92.135 ;
      LAYER met4 ;
        RECT 66.880 91.815 67.200 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 91.405 67.200 91.725 ;
      LAYER met4 ;
        RECT 66.880 91.405 67.200 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 90.995 67.200 91.315 ;
      LAYER met4 ;
        RECT 66.880 90.995 67.200 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 90.585 67.200 90.905 ;
      LAYER met4 ;
        RECT 66.880 90.585 67.200 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 90.175 67.200 90.495 ;
      LAYER met4 ;
        RECT 66.880 90.175 67.200 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 89.765 67.200 90.085 ;
      LAYER met4 ;
        RECT 66.880 89.765 67.200 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 89.355 67.200 89.675 ;
      LAYER met4 ;
        RECT 66.880 89.355 67.200 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 88.945 67.200 89.265 ;
      LAYER met4 ;
        RECT 66.880 88.945 67.200 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 88.535 67.200 88.855 ;
      LAYER met4 ;
        RECT 66.880 88.535 67.200 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 88.125 67.200 88.445 ;
      LAYER met4 ;
        RECT 66.880 88.125 67.200 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 87.715 67.200 88.035 ;
      LAYER met4 ;
        RECT 66.880 87.715 67.200 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 87.305 67.200 87.625 ;
      LAYER met4 ;
        RECT 66.880 87.305 67.200 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 86.895 67.200 87.215 ;
      LAYER met4 ;
        RECT 66.880 86.895 67.200 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 86.485 67.200 86.805 ;
      LAYER met4 ;
        RECT 66.880 86.485 67.200 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 86.075 67.200 86.395 ;
      LAYER met4 ;
        RECT 66.880 86.075 67.200 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 85.665 67.200 85.985 ;
      LAYER met4 ;
        RECT 66.880 85.665 67.200 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 85.255 67.200 85.575 ;
      LAYER met4 ;
        RECT 66.880 85.255 67.200 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 84.845 67.200 85.165 ;
      LAYER met4 ;
        RECT 66.880 84.845 67.200 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 84.435 67.200 84.755 ;
      LAYER met4 ;
        RECT 66.880 84.435 67.200 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 84.025 67.200 84.345 ;
      LAYER met4 ;
        RECT 66.880 84.025 67.200 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 83.615 67.200 83.935 ;
      LAYER met4 ;
        RECT 66.880 83.615 67.200 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 83.205 67.200 83.525 ;
      LAYER met4 ;
        RECT 66.880 83.205 67.200 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.880 82.795 67.200 83.115 ;
      LAYER met4 ;
        RECT 66.880 82.795 67.200 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 22.160 66.840 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 21.730 66.840 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 21.300 66.840 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 20.870 66.840 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 20.440 66.840 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 20.010 66.840 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 19.580 66.840 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 19.150 66.840 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 18.720 66.840 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 18.290 66.840 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.640 17.860 66.840 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 82.360 66.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 81.955 66.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 81.550 66.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 81.145 66.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 80.740 66.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 80.335 66.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 79.930 66.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 79.525 66.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 79.120 66.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 78.715 66.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 78.310 66.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 77.905 66.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 77.500 66.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 77.095 66.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 76.690 66.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 76.285 66.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 75.880 66.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 75.475 66.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 75.070 66.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 74.665 66.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 74.260 66.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 73.855 66.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 73.450 66.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 73.045 66.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 72.635 66.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 72.225 66.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 71.815 66.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 71.405 66.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 70.995 66.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 70.585 66.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 70.175 66.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 69.765 66.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 69.355 66.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 68.945 66.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 68.535 66.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.610 68.125 66.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.530 92.695 66.730 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 92.225 66.790 92.545 ;
      LAYER met4 ;
        RECT 66.470 92.225 66.790 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 91.815 66.790 92.135 ;
      LAYER met4 ;
        RECT 66.470 91.815 66.790 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 91.405 66.790 91.725 ;
      LAYER met4 ;
        RECT 66.470 91.405 66.790 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 90.995 66.790 91.315 ;
      LAYER met4 ;
        RECT 66.470 90.995 66.790 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 90.585 66.790 90.905 ;
      LAYER met4 ;
        RECT 66.470 90.585 66.790 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 90.175 66.790 90.495 ;
      LAYER met4 ;
        RECT 66.470 90.175 66.790 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 89.765 66.790 90.085 ;
      LAYER met4 ;
        RECT 66.470 89.765 66.790 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 89.355 66.790 89.675 ;
      LAYER met4 ;
        RECT 66.470 89.355 66.790 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 88.945 66.790 89.265 ;
      LAYER met4 ;
        RECT 66.470 88.945 66.790 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 88.535 66.790 88.855 ;
      LAYER met4 ;
        RECT 66.470 88.535 66.790 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 88.125 66.790 88.445 ;
      LAYER met4 ;
        RECT 66.470 88.125 66.790 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 87.715 66.790 88.035 ;
      LAYER met4 ;
        RECT 66.470 87.715 66.790 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 87.305 66.790 87.625 ;
      LAYER met4 ;
        RECT 66.470 87.305 66.790 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 86.895 66.790 87.215 ;
      LAYER met4 ;
        RECT 66.470 86.895 66.790 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 86.485 66.790 86.805 ;
      LAYER met4 ;
        RECT 66.470 86.485 66.790 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 86.075 66.790 86.395 ;
      LAYER met4 ;
        RECT 66.470 86.075 66.790 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 85.665 66.790 85.985 ;
      LAYER met4 ;
        RECT 66.470 85.665 66.790 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 85.255 66.790 85.575 ;
      LAYER met4 ;
        RECT 66.470 85.255 66.790 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 84.845 66.790 85.165 ;
      LAYER met4 ;
        RECT 66.470 84.845 66.790 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 84.435 66.790 84.755 ;
      LAYER met4 ;
        RECT 66.470 84.435 66.790 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 84.025 66.790 84.345 ;
      LAYER met4 ;
        RECT 66.470 84.025 66.790 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 83.615 66.790 83.935 ;
      LAYER met4 ;
        RECT 66.470 83.615 66.790 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 83.205 66.790 83.525 ;
      LAYER met4 ;
        RECT 66.470 83.205 66.790 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.470 82.795 66.790 83.115 ;
      LAYER met4 ;
        RECT 66.470 82.795 66.790 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 22.160 66.435 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 21.730 66.435 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 21.300 66.435 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 20.870 66.435 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 20.440 66.435 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 20.010 66.435 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 19.580 66.435 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 19.150 66.435 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 18.720 66.435 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 18.290 66.435 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.235 17.860 66.435 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 82.360 66.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 81.955 66.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 81.550 66.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 81.145 66.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 80.740 66.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 80.335 66.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 79.930 66.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 79.525 66.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 79.120 66.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 78.715 66.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 78.310 66.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 77.905 66.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 77.500 66.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 77.095 66.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 76.690 66.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 76.285 66.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 75.880 66.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 75.475 66.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 75.070 66.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 74.665 66.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 74.260 66.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 73.855 66.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 73.450 66.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 73.045 66.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 72.635 66.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 72.225 66.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 71.815 66.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 71.405 66.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 70.995 66.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 70.585 66.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 70.175 66.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 69.765 66.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 69.355 66.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 68.945 66.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 68.535 66.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.210 68.125 66.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.120 92.695 66.320 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 92.225 66.380 92.545 ;
      LAYER met4 ;
        RECT 66.060 92.225 66.380 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 91.815 66.380 92.135 ;
      LAYER met4 ;
        RECT 66.060 91.815 66.380 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 91.405 66.380 91.725 ;
      LAYER met4 ;
        RECT 66.060 91.405 66.380 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 90.995 66.380 91.315 ;
      LAYER met4 ;
        RECT 66.060 90.995 66.380 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 90.585 66.380 90.905 ;
      LAYER met4 ;
        RECT 66.060 90.585 66.380 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 90.175 66.380 90.495 ;
      LAYER met4 ;
        RECT 66.060 90.175 66.380 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 89.765 66.380 90.085 ;
      LAYER met4 ;
        RECT 66.060 89.765 66.380 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 89.355 66.380 89.675 ;
      LAYER met4 ;
        RECT 66.060 89.355 66.380 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 88.945 66.380 89.265 ;
      LAYER met4 ;
        RECT 66.060 88.945 66.380 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 88.535 66.380 88.855 ;
      LAYER met4 ;
        RECT 66.060 88.535 66.380 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 88.125 66.380 88.445 ;
      LAYER met4 ;
        RECT 66.060 88.125 66.380 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 87.715 66.380 88.035 ;
      LAYER met4 ;
        RECT 66.060 87.715 66.380 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 87.305 66.380 87.625 ;
      LAYER met4 ;
        RECT 66.060 87.305 66.380 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 86.895 66.380 87.215 ;
      LAYER met4 ;
        RECT 66.060 86.895 66.380 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 86.485 66.380 86.805 ;
      LAYER met4 ;
        RECT 66.060 86.485 66.380 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 86.075 66.380 86.395 ;
      LAYER met4 ;
        RECT 66.060 86.075 66.380 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 85.665 66.380 85.985 ;
      LAYER met4 ;
        RECT 66.060 85.665 66.380 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 85.255 66.380 85.575 ;
      LAYER met4 ;
        RECT 66.060 85.255 66.380 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 84.845 66.380 85.165 ;
      LAYER met4 ;
        RECT 66.060 84.845 66.380 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 84.435 66.380 84.755 ;
      LAYER met4 ;
        RECT 66.060 84.435 66.380 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 84.025 66.380 84.345 ;
      LAYER met4 ;
        RECT 66.060 84.025 66.380 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 83.615 66.380 83.935 ;
      LAYER met4 ;
        RECT 66.060 83.615 66.380 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 83.205 66.380 83.525 ;
      LAYER met4 ;
        RECT 66.060 83.205 66.380 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.060 82.795 66.380 83.115 ;
      LAYER met4 ;
        RECT 66.060 82.795 66.380 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 22.160 66.030 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 21.730 66.030 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 21.300 66.030 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 20.870 66.030 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 20.440 66.030 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 20.010 66.030 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 19.580 66.030 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 19.150 66.030 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 18.720 66.030 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 18.290 66.030 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 17.860 66.030 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 82.360 66.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 81.955 66.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 81.550 66.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 81.145 66.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 80.740 66.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 80.335 66.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 79.930 66.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 79.525 66.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 79.120 66.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 78.715 66.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 78.310 66.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 77.905 66.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 77.500 66.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 77.095 66.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 76.690 66.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 76.285 66.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 75.880 66.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 75.475 66.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 75.070 66.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 74.665 66.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 74.260 66.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 73.855 66.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 73.450 66.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 73.045 66.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 72.635 66.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 72.225 66.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 71.815 66.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 71.405 66.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 70.995 66.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 70.585 66.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 70.175 66.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 69.765 66.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 69.355 66.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 68.945 66.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 68.535 66.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.810 68.125 66.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.710 92.695 65.910 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 92.225 65.970 92.545 ;
      LAYER met4 ;
        RECT 65.650 92.225 65.970 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 91.815 65.970 92.135 ;
      LAYER met4 ;
        RECT 65.650 91.815 65.970 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 91.405 65.970 91.725 ;
      LAYER met4 ;
        RECT 65.650 91.405 65.970 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 90.995 65.970 91.315 ;
      LAYER met4 ;
        RECT 65.650 90.995 65.970 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 90.585 65.970 90.905 ;
      LAYER met4 ;
        RECT 65.650 90.585 65.970 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 90.175 65.970 90.495 ;
      LAYER met4 ;
        RECT 65.650 90.175 65.970 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 89.765 65.970 90.085 ;
      LAYER met4 ;
        RECT 65.650 89.765 65.970 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 89.355 65.970 89.675 ;
      LAYER met4 ;
        RECT 65.650 89.355 65.970 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 88.945 65.970 89.265 ;
      LAYER met4 ;
        RECT 65.650 88.945 65.970 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 88.535 65.970 88.855 ;
      LAYER met4 ;
        RECT 65.650 88.535 65.970 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 88.125 65.970 88.445 ;
      LAYER met4 ;
        RECT 65.650 88.125 65.970 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 87.715 65.970 88.035 ;
      LAYER met4 ;
        RECT 65.650 87.715 65.970 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 87.305 65.970 87.625 ;
      LAYER met4 ;
        RECT 65.650 87.305 65.970 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 86.895 65.970 87.215 ;
      LAYER met4 ;
        RECT 65.650 86.895 65.970 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 86.485 65.970 86.805 ;
      LAYER met4 ;
        RECT 65.650 86.485 65.970 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 86.075 65.970 86.395 ;
      LAYER met4 ;
        RECT 65.650 86.075 65.970 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 85.665 65.970 85.985 ;
      LAYER met4 ;
        RECT 65.650 85.665 65.970 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 85.255 65.970 85.575 ;
      LAYER met4 ;
        RECT 65.650 85.255 65.970 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 84.845 65.970 85.165 ;
      LAYER met4 ;
        RECT 65.650 84.845 65.970 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 84.435 65.970 84.755 ;
      LAYER met4 ;
        RECT 65.650 84.435 65.970 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 84.025 65.970 84.345 ;
      LAYER met4 ;
        RECT 65.650 84.025 65.970 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 83.615 65.970 83.935 ;
      LAYER met4 ;
        RECT 65.650 83.615 65.970 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 83.205 65.970 83.525 ;
      LAYER met4 ;
        RECT 65.650 83.205 65.970 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.650 82.795 65.970 83.115 ;
      LAYER met4 ;
        RECT 65.650 82.795 65.970 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 22.160 65.625 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 21.730 65.625 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 21.300 65.625 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 20.870 65.625 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 20.440 65.625 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 20.010 65.625 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 19.580 65.625 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 19.150 65.625 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 18.720 65.625 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 18.290 65.625 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.425 17.860 65.625 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 82.360 65.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 81.955 65.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 81.550 65.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 81.145 65.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 80.740 65.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 80.335 65.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 79.930 65.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 79.525 65.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 79.120 65.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 78.715 65.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 78.310 65.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 77.905 65.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 77.500 65.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 77.095 65.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 76.690 65.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 76.285 65.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 75.880 65.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 75.475 65.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 75.070 65.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 74.665 65.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 74.260 65.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 73.855 65.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 73.450 65.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 73.045 65.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 72.635 65.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 72.225 65.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 71.815 65.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 71.405 65.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 70.995 65.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 70.585 65.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 70.175 65.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 69.765 65.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 69.355 65.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 68.945 65.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 68.535 65.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.410 68.125 65.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.300 92.695 65.500 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 92.225 65.560 92.545 ;
      LAYER met4 ;
        RECT 65.240 92.225 65.560 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 91.815 65.560 92.135 ;
      LAYER met4 ;
        RECT 65.240 91.815 65.560 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 91.405 65.560 91.725 ;
      LAYER met4 ;
        RECT 65.240 91.405 65.560 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 90.995 65.560 91.315 ;
      LAYER met4 ;
        RECT 65.240 90.995 65.560 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 90.585 65.560 90.905 ;
      LAYER met4 ;
        RECT 65.240 90.585 65.560 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 90.175 65.560 90.495 ;
      LAYER met4 ;
        RECT 65.240 90.175 65.560 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 89.765 65.560 90.085 ;
      LAYER met4 ;
        RECT 65.240 89.765 65.560 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 89.355 65.560 89.675 ;
      LAYER met4 ;
        RECT 65.240 89.355 65.560 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 88.945 65.560 89.265 ;
      LAYER met4 ;
        RECT 65.240 88.945 65.560 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 88.535 65.560 88.855 ;
      LAYER met4 ;
        RECT 65.240 88.535 65.560 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 88.125 65.560 88.445 ;
      LAYER met4 ;
        RECT 65.240 88.125 65.560 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 87.715 65.560 88.035 ;
      LAYER met4 ;
        RECT 65.240 87.715 65.560 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 87.305 65.560 87.625 ;
      LAYER met4 ;
        RECT 65.240 87.305 65.560 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 86.895 65.560 87.215 ;
      LAYER met4 ;
        RECT 65.240 86.895 65.560 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 86.485 65.560 86.805 ;
      LAYER met4 ;
        RECT 65.240 86.485 65.560 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 86.075 65.560 86.395 ;
      LAYER met4 ;
        RECT 65.240 86.075 65.560 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 85.665 65.560 85.985 ;
      LAYER met4 ;
        RECT 65.240 85.665 65.560 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 85.255 65.560 85.575 ;
      LAYER met4 ;
        RECT 65.240 85.255 65.560 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 84.845 65.560 85.165 ;
      LAYER met4 ;
        RECT 65.240 84.845 65.560 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 84.435 65.560 84.755 ;
      LAYER met4 ;
        RECT 65.240 84.435 65.560 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 84.025 65.560 84.345 ;
      LAYER met4 ;
        RECT 65.240 84.025 65.560 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 83.615 65.560 83.935 ;
      LAYER met4 ;
        RECT 65.240 83.615 65.560 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 83.205 65.560 83.525 ;
      LAYER met4 ;
        RECT 65.240 83.205 65.560 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.240 82.795 65.560 83.115 ;
      LAYER met4 ;
        RECT 65.240 82.795 65.560 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 22.160 65.220 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 21.730 65.220 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 21.300 65.220 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 20.870 65.220 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 20.440 65.220 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 20.010 65.220 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 19.580 65.220 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 19.150 65.220 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 18.720 65.220 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 18.290 65.220 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.020 17.860 65.220 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 82.360 65.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 81.955 65.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 81.550 65.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 81.145 65.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 80.740 65.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 80.335 65.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 79.930 65.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 79.525 65.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 79.120 65.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 78.715 65.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 78.310 65.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 77.905 65.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 77.500 65.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 77.095 65.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 76.690 65.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 76.285 65.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 75.880 65.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 75.475 65.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 75.070 65.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 74.665 65.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 74.260 65.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 73.855 65.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 73.450 65.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 73.045 65.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 72.635 65.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 72.225 65.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 71.815 65.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 71.405 65.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 70.995 65.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 70.585 65.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 70.175 65.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 69.765 65.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 69.355 65.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 68.945 65.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 68.535 65.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 68.125 65.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.890 92.695 65.090 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 92.225 65.150 92.545 ;
      LAYER met4 ;
        RECT 64.830 92.225 65.150 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 91.815 65.150 92.135 ;
      LAYER met4 ;
        RECT 64.830 91.815 65.150 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 91.405 65.150 91.725 ;
      LAYER met4 ;
        RECT 64.830 91.405 65.150 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 90.995 65.150 91.315 ;
      LAYER met4 ;
        RECT 64.830 90.995 65.150 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 90.585 65.150 90.905 ;
      LAYER met4 ;
        RECT 64.830 90.585 65.150 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 90.175 65.150 90.495 ;
      LAYER met4 ;
        RECT 64.830 90.175 65.150 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 89.765 65.150 90.085 ;
      LAYER met4 ;
        RECT 64.830 89.765 65.150 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 89.355 65.150 89.675 ;
      LAYER met4 ;
        RECT 64.830 89.355 65.150 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 88.945 65.150 89.265 ;
      LAYER met4 ;
        RECT 64.830 88.945 65.150 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 88.535 65.150 88.855 ;
      LAYER met4 ;
        RECT 64.830 88.535 65.150 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 88.125 65.150 88.445 ;
      LAYER met4 ;
        RECT 64.830 88.125 65.150 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 87.715 65.150 88.035 ;
      LAYER met4 ;
        RECT 64.830 87.715 65.150 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 87.305 65.150 87.625 ;
      LAYER met4 ;
        RECT 64.830 87.305 65.150 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 86.895 65.150 87.215 ;
      LAYER met4 ;
        RECT 64.830 86.895 65.150 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 86.485 65.150 86.805 ;
      LAYER met4 ;
        RECT 64.830 86.485 65.150 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 86.075 65.150 86.395 ;
      LAYER met4 ;
        RECT 64.830 86.075 65.150 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 85.665 65.150 85.985 ;
      LAYER met4 ;
        RECT 64.830 85.665 65.150 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 85.255 65.150 85.575 ;
      LAYER met4 ;
        RECT 64.830 85.255 65.150 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 84.845 65.150 85.165 ;
      LAYER met4 ;
        RECT 64.830 84.845 65.150 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 84.435 65.150 84.755 ;
      LAYER met4 ;
        RECT 64.830 84.435 65.150 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 84.025 65.150 84.345 ;
      LAYER met4 ;
        RECT 64.830 84.025 65.150 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 83.615 65.150 83.935 ;
      LAYER met4 ;
        RECT 64.830 83.615 65.150 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 83.205 65.150 83.525 ;
      LAYER met4 ;
        RECT 64.830 83.205 65.150 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.830 82.795 65.150 83.115 ;
      LAYER met4 ;
        RECT 64.830 82.795 65.150 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 22.160 64.815 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 21.730 64.815 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 21.300 64.815 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 20.870 64.815 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 20.440 64.815 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 20.010 64.815 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 19.580 64.815 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 19.150 64.815 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 18.720 64.815 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 18.290 64.815 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.615 17.860 64.815 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 82.360 64.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 81.955 64.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 81.550 64.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 81.145 64.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 80.740 64.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 80.335 64.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 79.930 64.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 79.525 64.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 79.120 64.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 78.715 64.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 78.310 64.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 77.905 64.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 77.500 64.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 77.095 64.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 76.690 64.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 76.285 64.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 75.880 64.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 75.475 64.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 75.070 64.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 74.665 64.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 74.260 64.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 73.855 64.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 73.450 64.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 73.045 64.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 72.635 64.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 72.225 64.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 71.815 64.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 71.405 64.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 70.995 64.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 70.585 64.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 70.175 64.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 69.765 64.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 69.355 64.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 68.945 64.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 68.535 64.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.610 68.125 64.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.480 92.695 64.680 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 92.225 64.740 92.545 ;
      LAYER met4 ;
        RECT 64.420 92.225 64.740 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 91.815 64.740 92.135 ;
      LAYER met4 ;
        RECT 64.420 91.815 64.740 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 91.405 64.740 91.725 ;
      LAYER met4 ;
        RECT 64.420 91.405 64.740 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 90.995 64.740 91.315 ;
      LAYER met4 ;
        RECT 64.420 90.995 64.740 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 90.585 64.740 90.905 ;
      LAYER met4 ;
        RECT 64.420 90.585 64.740 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 90.175 64.740 90.495 ;
      LAYER met4 ;
        RECT 64.420 90.175 64.740 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 89.765 64.740 90.085 ;
      LAYER met4 ;
        RECT 64.420 89.765 64.740 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 89.355 64.740 89.675 ;
      LAYER met4 ;
        RECT 64.420 89.355 64.740 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 88.945 64.740 89.265 ;
      LAYER met4 ;
        RECT 64.420 88.945 64.740 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 88.535 64.740 88.855 ;
      LAYER met4 ;
        RECT 64.420 88.535 64.740 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 88.125 64.740 88.445 ;
      LAYER met4 ;
        RECT 64.420 88.125 64.740 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 87.715 64.740 88.035 ;
      LAYER met4 ;
        RECT 64.420 87.715 64.740 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 87.305 64.740 87.625 ;
      LAYER met4 ;
        RECT 64.420 87.305 64.740 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 86.895 64.740 87.215 ;
      LAYER met4 ;
        RECT 64.420 86.895 64.740 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 86.485 64.740 86.805 ;
      LAYER met4 ;
        RECT 64.420 86.485 64.740 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 86.075 64.740 86.395 ;
      LAYER met4 ;
        RECT 64.420 86.075 64.740 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 85.665 64.740 85.985 ;
      LAYER met4 ;
        RECT 64.420 85.665 64.740 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 85.255 64.740 85.575 ;
      LAYER met4 ;
        RECT 64.420 85.255 64.740 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 84.845 64.740 85.165 ;
      LAYER met4 ;
        RECT 64.420 84.845 64.740 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 84.435 64.740 84.755 ;
      LAYER met4 ;
        RECT 64.420 84.435 64.740 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 84.025 64.740 84.345 ;
      LAYER met4 ;
        RECT 64.420 84.025 64.740 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 83.615 64.740 83.935 ;
      LAYER met4 ;
        RECT 64.420 83.615 64.740 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 83.205 64.740 83.525 ;
      LAYER met4 ;
        RECT 64.420 83.205 64.740 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.420 82.795 64.740 83.115 ;
      LAYER met4 ;
        RECT 64.420 82.795 64.740 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 82.360 64.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 81.955 64.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 81.550 64.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 81.145 64.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 80.740 64.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 80.335 64.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 79.930 64.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 79.525 64.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 79.120 64.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 78.715 64.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 78.310 64.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 77.905 64.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 77.500 64.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 77.095 64.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 76.690 64.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 76.285 64.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 75.880 64.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 75.475 64.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 75.070 64.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 74.665 64.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 74.260 64.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 73.855 64.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 73.450 64.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 73.045 64.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 72.635 64.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 72.225 64.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 71.815 64.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 71.405 64.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 70.995 64.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 70.585 64.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 70.175 64.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 69.765 64.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 69.355 64.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 68.945 64.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 68.535 64.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 68.125 64.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 22.160 64.410 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 21.730 64.410 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 21.300 64.410 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 20.870 64.410 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 20.440 64.410 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 20.010 64.410 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 19.580 64.410 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 19.150 64.410 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 18.720 64.410 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 18.290 64.410 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.210 17.860 64.410 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.070 92.695 64.270 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 92.225 64.330 92.545 ;
      LAYER met4 ;
        RECT 64.010 92.225 64.330 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 91.815 64.330 92.135 ;
      LAYER met4 ;
        RECT 64.010 91.815 64.330 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 91.405 64.330 91.725 ;
      LAYER met4 ;
        RECT 64.010 91.405 64.330 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 90.995 64.330 91.315 ;
      LAYER met4 ;
        RECT 64.010 90.995 64.330 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 90.585 64.330 90.905 ;
      LAYER met4 ;
        RECT 64.010 90.585 64.330 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 90.175 64.330 90.495 ;
      LAYER met4 ;
        RECT 64.010 90.175 64.330 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 89.765 64.330 90.085 ;
      LAYER met4 ;
        RECT 64.010 89.765 64.330 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 89.355 64.330 89.675 ;
      LAYER met4 ;
        RECT 64.010 89.355 64.330 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 88.945 64.330 89.265 ;
      LAYER met4 ;
        RECT 64.010 88.945 64.330 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 88.535 64.330 88.855 ;
      LAYER met4 ;
        RECT 64.010 88.535 64.330 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 88.125 64.330 88.445 ;
      LAYER met4 ;
        RECT 64.010 88.125 64.330 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 87.715 64.330 88.035 ;
      LAYER met4 ;
        RECT 64.010 87.715 64.330 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 87.305 64.330 87.625 ;
      LAYER met4 ;
        RECT 64.010 87.305 64.330 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 86.895 64.330 87.215 ;
      LAYER met4 ;
        RECT 64.010 86.895 64.330 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 86.485 64.330 86.805 ;
      LAYER met4 ;
        RECT 64.010 86.485 64.330 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 86.075 64.330 86.395 ;
      LAYER met4 ;
        RECT 64.010 86.075 64.330 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 85.665 64.330 85.985 ;
      LAYER met4 ;
        RECT 64.010 85.665 64.330 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 85.255 64.330 85.575 ;
      LAYER met4 ;
        RECT 64.010 85.255 64.330 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 84.845 64.330 85.165 ;
      LAYER met4 ;
        RECT 64.010 84.845 64.330 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 84.435 64.330 84.755 ;
      LAYER met4 ;
        RECT 64.010 84.435 64.330 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 84.025 64.330 84.345 ;
      LAYER met4 ;
        RECT 64.010 84.025 64.330 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 83.615 64.330 83.935 ;
      LAYER met4 ;
        RECT 64.010 83.615 64.330 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 83.205 64.330 83.525 ;
      LAYER met4 ;
        RECT 64.010 83.205 64.330 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.010 82.795 64.330 83.115 ;
      LAYER met4 ;
        RECT 64.010 82.795 64.330 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 82.360 64.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 81.955 64.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 81.550 64.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 81.145 64.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 80.740 64.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 80.335 64.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 79.930 64.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 79.525 64.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 79.120 64.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 78.715 64.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 78.310 64.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 77.905 64.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 77.500 64.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 77.095 64.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 76.690 64.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 76.285 64.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 75.880 64.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 75.475 64.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 75.070 64.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 74.665 64.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 74.260 64.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 73.855 64.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 73.450 64.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 73.045 64.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 72.635 64.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 72.225 64.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 71.815 64.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 71.405 64.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 70.995 64.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 70.585 64.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 70.175 64.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 69.765 64.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 69.355 64.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 68.945 64.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 68.535 64.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.810 68.125 64.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 22.160 64.005 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 21.730 64.005 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 21.300 64.005 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 20.870 64.005 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 20.440 64.005 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 20.010 64.005 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 19.580 64.005 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 19.150 64.005 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 18.720 64.005 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 18.290 64.005 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.805 17.860 64.005 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.660 92.695 63.860 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 92.225 63.920 92.545 ;
      LAYER met4 ;
        RECT 63.600 92.225 63.920 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 91.815 63.920 92.135 ;
      LAYER met4 ;
        RECT 63.600 91.815 63.920 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 91.405 63.920 91.725 ;
      LAYER met4 ;
        RECT 63.600 91.405 63.920 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 90.995 63.920 91.315 ;
      LAYER met4 ;
        RECT 63.600 90.995 63.920 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 90.585 63.920 90.905 ;
      LAYER met4 ;
        RECT 63.600 90.585 63.920 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 90.175 63.920 90.495 ;
      LAYER met4 ;
        RECT 63.600 90.175 63.920 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 89.765 63.920 90.085 ;
      LAYER met4 ;
        RECT 63.600 89.765 63.920 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 89.355 63.920 89.675 ;
      LAYER met4 ;
        RECT 63.600 89.355 63.920 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 88.945 63.920 89.265 ;
      LAYER met4 ;
        RECT 63.600 88.945 63.920 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 88.535 63.920 88.855 ;
      LAYER met4 ;
        RECT 63.600 88.535 63.920 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 88.125 63.920 88.445 ;
      LAYER met4 ;
        RECT 63.600 88.125 63.920 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 87.715 63.920 88.035 ;
      LAYER met4 ;
        RECT 63.600 87.715 63.920 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 87.305 63.920 87.625 ;
      LAYER met4 ;
        RECT 63.600 87.305 63.920 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 86.895 63.920 87.215 ;
      LAYER met4 ;
        RECT 63.600 86.895 63.920 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 86.485 63.920 86.805 ;
      LAYER met4 ;
        RECT 63.600 86.485 63.920 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 86.075 63.920 86.395 ;
      LAYER met4 ;
        RECT 63.600 86.075 63.920 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 85.665 63.920 85.985 ;
      LAYER met4 ;
        RECT 63.600 85.665 63.920 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 85.255 63.920 85.575 ;
      LAYER met4 ;
        RECT 63.600 85.255 63.920 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 84.845 63.920 85.165 ;
      LAYER met4 ;
        RECT 63.600 84.845 63.920 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 84.435 63.920 84.755 ;
      LAYER met4 ;
        RECT 63.600 84.435 63.920 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 84.025 63.920 84.345 ;
      LAYER met4 ;
        RECT 63.600 84.025 63.920 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 83.615 63.920 83.935 ;
      LAYER met4 ;
        RECT 63.600 83.615 63.920 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 83.205 63.920 83.525 ;
      LAYER met4 ;
        RECT 63.600 83.205 63.920 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.600 82.795 63.920 83.115 ;
      LAYER met4 ;
        RECT 63.600 82.795 63.920 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 82.360 63.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 81.955 63.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 81.550 63.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 81.145 63.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 80.740 63.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 80.335 63.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 79.930 63.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 79.525 63.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 79.120 63.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 78.715 63.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 78.310 63.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 77.905 63.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 77.500 63.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 77.095 63.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 76.690 63.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 76.285 63.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 75.880 63.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 75.475 63.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 75.070 63.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 74.665 63.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 74.260 63.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 73.855 63.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 73.450 63.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 73.045 63.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 72.635 63.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 72.225 63.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 71.815 63.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 71.405 63.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 70.995 63.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 70.585 63.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 70.175 63.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 69.765 63.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 69.355 63.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 68.945 63.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 68.535 63.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 68.125 63.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 22.160 63.600 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 21.730 63.600 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 21.300 63.600 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 20.870 63.600 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 20.440 63.600 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 20.010 63.600 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 19.580 63.600 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 19.150 63.600 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 18.720 63.600 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 18.290 63.600 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.400 17.860 63.600 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.250 92.695 63.450 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 92.225 63.510 92.545 ;
      LAYER met4 ;
        RECT 63.190 92.225 63.510 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 91.815 63.510 92.135 ;
      LAYER met4 ;
        RECT 63.190 91.815 63.510 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 91.405 63.510 91.725 ;
      LAYER met4 ;
        RECT 63.190 91.405 63.510 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 90.995 63.510 91.315 ;
      LAYER met4 ;
        RECT 63.190 90.995 63.510 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 90.585 63.510 90.905 ;
      LAYER met4 ;
        RECT 63.190 90.585 63.510 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 90.175 63.510 90.495 ;
      LAYER met4 ;
        RECT 63.190 90.175 63.510 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 89.765 63.510 90.085 ;
      LAYER met4 ;
        RECT 63.190 89.765 63.510 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 89.355 63.510 89.675 ;
      LAYER met4 ;
        RECT 63.190 89.355 63.510 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 88.945 63.510 89.265 ;
      LAYER met4 ;
        RECT 63.190 88.945 63.510 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 88.535 63.510 88.855 ;
      LAYER met4 ;
        RECT 63.190 88.535 63.510 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 88.125 63.510 88.445 ;
      LAYER met4 ;
        RECT 63.190 88.125 63.510 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 87.715 63.510 88.035 ;
      LAYER met4 ;
        RECT 63.190 87.715 63.510 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 87.305 63.510 87.625 ;
      LAYER met4 ;
        RECT 63.190 87.305 63.510 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 86.895 63.510 87.215 ;
      LAYER met4 ;
        RECT 63.190 86.895 63.510 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 86.485 63.510 86.805 ;
      LAYER met4 ;
        RECT 63.190 86.485 63.510 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 86.075 63.510 86.395 ;
      LAYER met4 ;
        RECT 63.190 86.075 63.510 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 85.665 63.510 85.985 ;
      LAYER met4 ;
        RECT 63.190 85.665 63.510 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 85.255 63.510 85.575 ;
      LAYER met4 ;
        RECT 63.190 85.255 63.510 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 84.845 63.510 85.165 ;
      LAYER met4 ;
        RECT 63.190 84.845 63.510 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 84.435 63.510 84.755 ;
      LAYER met4 ;
        RECT 63.190 84.435 63.510 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 84.025 63.510 84.345 ;
      LAYER met4 ;
        RECT 63.190 84.025 63.510 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 83.615 63.510 83.935 ;
      LAYER met4 ;
        RECT 63.190 83.615 63.510 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 83.205 63.510 83.525 ;
      LAYER met4 ;
        RECT 63.190 83.205 63.510 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.190 82.795 63.510 83.115 ;
      LAYER met4 ;
        RECT 63.190 82.795 63.510 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 82.360 63.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 81.955 63.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 81.550 63.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 81.145 63.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 80.740 63.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 80.335 63.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 79.930 63.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 79.525 63.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 79.120 63.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 78.715 63.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 78.310 63.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 77.905 63.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 77.500 63.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 77.095 63.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 76.690 63.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 76.285 63.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 75.880 63.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 75.475 63.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 75.070 63.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 74.665 63.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 74.260 63.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 73.855 63.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 73.450 63.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 73.045 63.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 72.635 63.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 72.225 63.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 71.815 63.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 71.405 63.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 70.995 63.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 70.585 63.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 70.175 63.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 69.765 63.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 69.355 63.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 68.945 63.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 68.535 63.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.010 68.125 63.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 22.160 63.195 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 21.730 63.195 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 21.300 63.195 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 20.870 63.195 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 20.440 63.195 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 20.010 63.195 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 19.580 63.195 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 19.150 63.195 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 18.720 63.195 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 18.290 63.195 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.995 17.860 63.195 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.840 92.695 63.040 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 92.225 63.100 92.545 ;
      LAYER met4 ;
        RECT 62.780 92.225 63.100 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 91.815 63.100 92.135 ;
      LAYER met4 ;
        RECT 62.780 91.815 63.100 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 91.405 63.100 91.725 ;
      LAYER met4 ;
        RECT 62.780 91.405 63.100 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 90.995 63.100 91.315 ;
      LAYER met4 ;
        RECT 62.780 90.995 63.100 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 90.585 63.100 90.905 ;
      LAYER met4 ;
        RECT 62.780 90.585 63.100 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 90.175 63.100 90.495 ;
      LAYER met4 ;
        RECT 62.780 90.175 63.100 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 89.765 63.100 90.085 ;
      LAYER met4 ;
        RECT 62.780 89.765 63.100 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 89.355 63.100 89.675 ;
      LAYER met4 ;
        RECT 62.780 89.355 63.100 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 88.945 63.100 89.265 ;
      LAYER met4 ;
        RECT 62.780 88.945 63.100 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 88.535 63.100 88.855 ;
      LAYER met4 ;
        RECT 62.780 88.535 63.100 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 88.125 63.100 88.445 ;
      LAYER met4 ;
        RECT 62.780 88.125 63.100 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 87.715 63.100 88.035 ;
      LAYER met4 ;
        RECT 62.780 87.715 63.100 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 87.305 63.100 87.625 ;
      LAYER met4 ;
        RECT 62.780 87.305 63.100 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 86.895 63.100 87.215 ;
      LAYER met4 ;
        RECT 62.780 86.895 63.100 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 86.485 63.100 86.805 ;
      LAYER met4 ;
        RECT 62.780 86.485 63.100 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 86.075 63.100 86.395 ;
      LAYER met4 ;
        RECT 62.780 86.075 63.100 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 85.665 63.100 85.985 ;
      LAYER met4 ;
        RECT 62.780 85.665 63.100 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 85.255 63.100 85.575 ;
      LAYER met4 ;
        RECT 62.780 85.255 63.100 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 84.845 63.100 85.165 ;
      LAYER met4 ;
        RECT 62.780 84.845 63.100 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 84.435 63.100 84.755 ;
      LAYER met4 ;
        RECT 62.780 84.435 63.100 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 84.025 63.100 84.345 ;
      LAYER met4 ;
        RECT 62.780 84.025 63.100 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 83.615 63.100 83.935 ;
      LAYER met4 ;
        RECT 62.780 83.615 63.100 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 83.205 63.100 83.525 ;
      LAYER met4 ;
        RECT 62.780 83.205 63.100 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.780 82.795 63.100 83.115 ;
      LAYER met4 ;
        RECT 62.780 82.795 63.100 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 82.360 62.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 81.955 62.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 81.550 62.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 81.145 62.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 80.740 62.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 80.335 62.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 79.930 62.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 79.525 62.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 79.120 62.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 78.715 62.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 78.310 62.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 77.905 62.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 77.500 62.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 77.095 62.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 76.690 62.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 76.285 62.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 75.880 62.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 75.475 62.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 75.070 62.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 74.665 62.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 74.260 62.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 73.855 62.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 73.450 62.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 73.045 62.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 72.635 62.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 72.225 62.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 71.815 62.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 71.405 62.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 70.995 62.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 70.585 62.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 70.175 62.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 69.765 62.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 69.355 62.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 68.945 62.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 68.535 62.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.610 68.125 62.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 22.160 62.790 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 21.730 62.790 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 21.300 62.790 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 20.870 62.790 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 20.440 62.790 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 20.010 62.790 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 19.580 62.790 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 19.150 62.790 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 18.720 62.790 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 18.290 62.790 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.590 17.860 62.790 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.430 92.695 62.630 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 92.225 62.690 92.545 ;
      LAYER met4 ;
        RECT 62.370 92.225 62.690 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 91.815 62.690 92.135 ;
      LAYER met4 ;
        RECT 62.370 91.815 62.690 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 91.405 62.690 91.725 ;
      LAYER met4 ;
        RECT 62.370 91.405 62.690 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 90.995 62.690 91.315 ;
      LAYER met4 ;
        RECT 62.370 90.995 62.690 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 90.585 62.690 90.905 ;
      LAYER met4 ;
        RECT 62.370 90.585 62.690 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 90.175 62.690 90.495 ;
      LAYER met4 ;
        RECT 62.370 90.175 62.690 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 89.765 62.690 90.085 ;
      LAYER met4 ;
        RECT 62.370 89.765 62.690 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 89.355 62.690 89.675 ;
      LAYER met4 ;
        RECT 62.370 89.355 62.690 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 88.945 62.690 89.265 ;
      LAYER met4 ;
        RECT 62.370 88.945 62.690 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 88.535 62.690 88.855 ;
      LAYER met4 ;
        RECT 62.370 88.535 62.690 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 88.125 62.690 88.445 ;
      LAYER met4 ;
        RECT 62.370 88.125 62.690 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 87.715 62.690 88.035 ;
      LAYER met4 ;
        RECT 62.370 87.715 62.690 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 87.305 62.690 87.625 ;
      LAYER met4 ;
        RECT 62.370 87.305 62.690 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 86.895 62.690 87.215 ;
      LAYER met4 ;
        RECT 62.370 86.895 62.690 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 86.485 62.690 86.805 ;
      LAYER met4 ;
        RECT 62.370 86.485 62.690 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 86.075 62.690 86.395 ;
      LAYER met4 ;
        RECT 62.370 86.075 62.690 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 85.665 62.690 85.985 ;
      LAYER met4 ;
        RECT 62.370 85.665 62.690 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 85.255 62.690 85.575 ;
      LAYER met4 ;
        RECT 62.370 85.255 62.690 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 84.845 62.690 85.165 ;
      LAYER met4 ;
        RECT 62.370 84.845 62.690 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 84.435 62.690 84.755 ;
      LAYER met4 ;
        RECT 62.370 84.435 62.690 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 84.025 62.690 84.345 ;
      LAYER met4 ;
        RECT 62.370 84.025 62.690 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 83.615 62.690 83.935 ;
      LAYER met4 ;
        RECT 62.370 83.615 62.690 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 83.205 62.690 83.525 ;
      LAYER met4 ;
        RECT 62.370 83.205 62.690 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.370 82.795 62.690 83.115 ;
      LAYER met4 ;
        RECT 62.370 82.795 62.690 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 82.360 62.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 81.955 62.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 81.550 62.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 81.145 62.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 80.740 62.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 80.335 62.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 79.930 62.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 79.525 62.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 79.120 62.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 78.715 62.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 78.310 62.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 77.905 62.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 77.500 62.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 77.095 62.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 76.690 62.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 76.285 62.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 75.880 62.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 75.475 62.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 75.070 62.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 74.665 62.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 74.260 62.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 73.855 62.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 73.450 62.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 73.045 62.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 72.635 62.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 72.225 62.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 71.815 62.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 71.405 62.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 70.995 62.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 70.585 62.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 70.175 62.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 69.765 62.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 69.355 62.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 68.945 62.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 68.535 62.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.210 68.125 62.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 22.160 62.385 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 21.730 62.385 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 21.300 62.385 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 20.870 62.385 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 20.440 62.385 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 20.010 62.385 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 19.580 62.385 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 19.150 62.385 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 18.720 62.385 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 18.290 62.385 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.185 17.860 62.385 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.025 92.695 62.225 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 92.225 62.285 92.545 ;
      LAYER met4 ;
        RECT 61.965 92.225 62.285 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 91.815 62.285 92.135 ;
      LAYER met4 ;
        RECT 61.965 91.815 62.285 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 91.405 62.285 91.725 ;
      LAYER met4 ;
        RECT 61.965 91.405 62.285 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 90.995 62.285 91.315 ;
      LAYER met4 ;
        RECT 61.965 90.995 62.285 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 90.585 62.285 90.905 ;
      LAYER met4 ;
        RECT 61.965 90.585 62.285 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 90.175 62.285 90.495 ;
      LAYER met4 ;
        RECT 61.965 90.175 62.285 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 89.765 62.285 90.085 ;
      LAYER met4 ;
        RECT 61.965 89.765 62.285 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 89.355 62.285 89.675 ;
      LAYER met4 ;
        RECT 61.965 89.355 62.285 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 88.945 62.285 89.265 ;
      LAYER met4 ;
        RECT 61.965 88.945 62.285 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 88.535 62.285 88.855 ;
      LAYER met4 ;
        RECT 61.965 88.535 62.285 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 88.125 62.285 88.445 ;
      LAYER met4 ;
        RECT 61.965 88.125 62.285 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 87.715 62.285 88.035 ;
      LAYER met4 ;
        RECT 61.965 87.715 62.285 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 87.305 62.285 87.625 ;
      LAYER met4 ;
        RECT 61.965 87.305 62.285 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 86.895 62.285 87.215 ;
      LAYER met4 ;
        RECT 61.965 86.895 62.285 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 86.485 62.285 86.805 ;
      LAYER met4 ;
        RECT 61.965 86.485 62.285 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 86.075 62.285 86.395 ;
      LAYER met4 ;
        RECT 61.965 86.075 62.285 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 85.665 62.285 85.985 ;
      LAYER met4 ;
        RECT 61.965 85.665 62.285 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 85.255 62.285 85.575 ;
      LAYER met4 ;
        RECT 61.965 85.255 62.285 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 84.845 62.285 85.165 ;
      LAYER met4 ;
        RECT 61.965 84.845 62.285 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 84.435 62.285 84.755 ;
      LAYER met4 ;
        RECT 61.965 84.435 62.285 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 84.025 62.285 84.345 ;
      LAYER met4 ;
        RECT 61.965 84.025 62.285 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 83.615 62.285 83.935 ;
      LAYER met4 ;
        RECT 61.965 83.615 62.285 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 83.205 62.285 83.525 ;
      LAYER met4 ;
        RECT 61.965 83.205 62.285 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.965 82.795 62.285 83.115 ;
      LAYER met4 ;
        RECT 61.965 82.795 62.285 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 82.360 62.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 81.955 62.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 81.550 62.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 81.145 62.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 80.740 62.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 80.335 62.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 79.930 62.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 79.525 62.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 79.120 62.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 78.715 62.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 78.310 62.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 77.905 62.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 77.500 62.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 77.095 62.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 76.690 62.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 76.285 62.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 75.880 62.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 75.475 62.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 75.070 62.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 74.665 62.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 74.260 62.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 73.855 62.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 73.450 62.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 73.045 62.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 72.635 62.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 72.225 62.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 71.815 62.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 71.405 62.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 70.995 62.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 70.585 62.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 70.175 62.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 69.765 62.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 69.355 62.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 68.945 62.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 68.535 62.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 68.125 62.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 22.160 61.980 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 21.730 61.980 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 21.300 61.980 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 20.870 61.980 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 20.440 61.980 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 20.010 61.980 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 19.580 61.980 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 19.150 61.980 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 18.720 61.980 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 18.290 61.980 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.780 17.860 61.980 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.620 92.695 61.820 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 92.225 61.880 92.545 ;
      LAYER met4 ;
        RECT 61.560 92.225 61.880 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 91.815 61.880 92.135 ;
      LAYER met4 ;
        RECT 61.560 91.815 61.880 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 91.405 61.880 91.725 ;
      LAYER met4 ;
        RECT 61.560 91.405 61.880 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 90.995 61.880 91.315 ;
      LAYER met4 ;
        RECT 61.560 90.995 61.880 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 90.585 61.880 90.905 ;
      LAYER met4 ;
        RECT 61.560 90.585 61.880 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 90.175 61.880 90.495 ;
      LAYER met4 ;
        RECT 61.560 90.175 61.880 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 89.765 61.880 90.085 ;
      LAYER met4 ;
        RECT 61.560 89.765 61.880 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 89.355 61.880 89.675 ;
      LAYER met4 ;
        RECT 61.560 89.355 61.880 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 88.945 61.880 89.265 ;
      LAYER met4 ;
        RECT 61.560 88.945 61.880 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 88.535 61.880 88.855 ;
      LAYER met4 ;
        RECT 61.560 88.535 61.880 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 88.125 61.880 88.445 ;
      LAYER met4 ;
        RECT 61.560 88.125 61.880 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 87.715 61.880 88.035 ;
      LAYER met4 ;
        RECT 61.560 87.715 61.880 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 87.305 61.880 87.625 ;
      LAYER met4 ;
        RECT 61.560 87.305 61.880 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 86.895 61.880 87.215 ;
      LAYER met4 ;
        RECT 61.560 86.895 61.880 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 86.485 61.880 86.805 ;
      LAYER met4 ;
        RECT 61.560 86.485 61.880 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 86.075 61.880 86.395 ;
      LAYER met4 ;
        RECT 61.560 86.075 61.880 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 85.665 61.880 85.985 ;
      LAYER met4 ;
        RECT 61.560 85.665 61.880 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 85.255 61.880 85.575 ;
      LAYER met4 ;
        RECT 61.560 85.255 61.880 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 84.845 61.880 85.165 ;
      LAYER met4 ;
        RECT 61.560 84.845 61.880 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 84.435 61.880 84.755 ;
      LAYER met4 ;
        RECT 61.560 84.435 61.880 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 84.025 61.880 84.345 ;
      LAYER met4 ;
        RECT 61.560 84.025 61.880 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 83.615 61.880 83.935 ;
      LAYER met4 ;
        RECT 61.560 83.615 61.880 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 83.205 61.880 83.525 ;
      LAYER met4 ;
        RECT 61.560 83.205 61.880 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.560 82.795 61.880 83.115 ;
      LAYER met4 ;
        RECT 61.560 82.795 61.880 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 82.360 61.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 81.955 61.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 81.550 61.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 81.145 61.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 80.740 61.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 80.335 61.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 79.930 61.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 79.525 61.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 79.120 61.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 78.715 61.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 78.310 61.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 77.905 61.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 77.500 61.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 77.095 61.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 76.690 61.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 76.285 61.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 75.880 61.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 75.475 61.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 75.070 61.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 74.665 61.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 74.260 61.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 73.855 61.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 73.450 61.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 73.045 61.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 72.635 61.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 72.225 61.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 71.815 61.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 71.405 61.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 70.995 61.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 70.585 61.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 70.175 61.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 69.765 61.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 69.355 61.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 68.945 61.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 68.535 61.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.410 68.125 61.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 22.160 61.575 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 21.730 61.575 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 21.300 61.575 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 20.870 61.575 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 20.440 61.575 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 20.010 61.575 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 19.580 61.575 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 19.150 61.575 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 18.720 61.575 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 18.290 61.575 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.375 17.860 61.575 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.215 92.695 61.415 92.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 92.225 61.475 92.545 ;
      LAYER met4 ;
        RECT 61.155 92.225 61.475 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 91.815 61.475 92.135 ;
      LAYER met4 ;
        RECT 61.155 91.815 61.475 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 91.405 61.475 91.725 ;
      LAYER met4 ;
        RECT 61.155 91.405 61.475 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 90.995 61.475 91.315 ;
      LAYER met4 ;
        RECT 61.155 90.995 61.475 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 90.585 61.475 90.905 ;
      LAYER met4 ;
        RECT 61.155 90.585 61.475 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 90.175 61.475 90.495 ;
      LAYER met4 ;
        RECT 61.155 90.175 61.475 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 89.765 61.475 90.085 ;
      LAYER met4 ;
        RECT 61.155 89.765 61.475 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 89.355 61.475 89.675 ;
      LAYER met4 ;
        RECT 61.155 89.355 61.475 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 88.945 61.475 89.265 ;
      LAYER met4 ;
        RECT 61.155 88.945 61.475 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 88.535 61.475 88.855 ;
      LAYER met4 ;
        RECT 61.155 88.535 61.475 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 88.125 61.475 88.445 ;
      LAYER met4 ;
        RECT 61.155 88.125 61.475 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 87.715 61.475 88.035 ;
      LAYER met4 ;
        RECT 61.155 87.715 61.475 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 87.305 61.475 87.625 ;
      LAYER met4 ;
        RECT 61.155 87.305 61.475 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 86.895 61.475 87.215 ;
      LAYER met4 ;
        RECT 61.155 86.895 61.475 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 86.485 61.475 86.805 ;
      LAYER met4 ;
        RECT 61.155 86.485 61.475 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 86.075 61.475 86.395 ;
      LAYER met4 ;
        RECT 61.155 86.075 61.475 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 85.665 61.475 85.985 ;
      LAYER met4 ;
        RECT 61.155 85.665 61.475 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 85.255 61.475 85.575 ;
      LAYER met4 ;
        RECT 61.155 85.255 61.475 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 84.845 61.475 85.165 ;
      LAYER met4 ;
        RECT 61.155 84.845 61.475 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 84.435 61.475 84.755 ;
      LAYER met4 ;
        RECT 61.155 84.435 61.475 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 84.025 61.475 84.345 ;
      LAYER met4 ;
        RECT 61.155 84.025 61.475 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 83.615 61.475 83.935 ;
      LAYER met4 ;
        RECT 61.155 83.615 61.475 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 83.205 61.475 83.525 ;
      LAYER met4 ;
        RECT 61.155 83.205 61.475 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.155 82.795 61.475 83.115 ;
      LAYER met4 ;
        RECT 61.155 82.795 61.475 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 82.360 61.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 81.955 61.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 81.550 61.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 81.145 61.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 80.740 61.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 80.335 61.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 79.930 61.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 79.525 61.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 79.120 61.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 78.715 61.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 78.310 61.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 77.905 61.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 77.500 61.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 77.095 61.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 76.690 61.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 76.285 61.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 75.880 61.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 75.475 61.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 75.070 61.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 74.665 61.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 74.260 61.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 73.855 61.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 73.450 61.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 73.045 61.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 72.635 61.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 72.225 61.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 71.815 61.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 71.405 61.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 70.995 61.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 70.585 61.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 70.175 61.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 69.765 61.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 69.355 61.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 68.945 61.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 68.535 61.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 68.125 61.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 22.160 61.170 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 21.730 61.170 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 21.300 61.170 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 20.870 61.170 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 20.440 61.170 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 20.010 61.170 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 19.580 61.170 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 19.150 61.170 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 18.720 61.170 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 18.290 61.170 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.970 17.860 61.170 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.675 91.385 60.995 91.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.675 90.955 60.995 91.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655 90.495 60.975 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655 90.065 60.975 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655 89.635 60.975 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655 89.205 60.975 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655 88.775 60.975 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.655 88.350 60.975 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 82.360 60.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 81.955 60.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 81.550 60.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 81.145 60.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 80.740 60.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 80.335 60.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 79.930 60.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 79.525 60.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 79.120 60.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 78.715 60.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 78.310 60.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 77.905 60.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 77.500 60.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 77.095 60.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 76.690 60.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 76.285 60.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 75.880 60.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 75.475 60.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 75.070 60.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 74.665 60.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 74.260 60.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 73.855 60.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 73.450 60.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 73.045 60.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 72.635 60.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 72.225 60.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 71.815 60.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 71.405 60.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 70.995 60.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 70.585 60.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 70.175 60.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 69.765 60.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 69.355 60.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 68.945 60.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 68.535 60.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.610 68.125 60.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 87.815 60.850 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 87.410 60.850 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 87.005 60.850 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 86.600 60.850 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 86.195 60.850 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 85.795 60.850 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 85.395 60.850 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 84.995 60.850 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 84.595 60.850 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 84.195 60.850 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 83.795 60.850 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 83.395 60.850 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.530 82.995 60.850 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 22.160 60.765 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 21.730 60.765 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 21.300 60.765 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 20.870 60.765 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 20.440 60.765 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 20.010 60.765 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 19.580 60.765 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 19.150 60.765 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 18.720 60.765 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 18.290 60.765 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.565 17.860 60.765 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245 90.495 60.565 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245 90.065 60.565 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245 89.635 60.565 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245 89.205 60.565 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245 88.775 60.565 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.245 88.350 60.565 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 82.360 60.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 81.955 60.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 81.550 60.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 81.145 60.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 80.740 60.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 80.335 60.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 79.930 60.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 79.525 60.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 79.120 60.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 78.715 60.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 78.310 60.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 77.905 60.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 77.500 60.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 77.095 60.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 76.690 60.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 76.285 60.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 75.880 60.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 75.475 60.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 75.070 60.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 74.665 60.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 74.260 60.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 73.855 60.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 73.450 60.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 73.045 60.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 72.635 60.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 72.225 60.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 71.815 60.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 71.405 60.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 70.995 60.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 70.585 60.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 70.175 60.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 69.765 60.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 69.355 60.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 68.945 60.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 68.535 60.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.210 68.125 60.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 87.815 60.440 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 87.410 60.440 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 87.005 60.440 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 86.600 60.440 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 86.195 60.440 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 85.795 60.440 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 85.395 60.440 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 84.995 60.440 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 84.595 60.440 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 84.195 60.440 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 83.795 60.440 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 83.395 60.440 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.120 82.995 60.440 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 22.160 60.360 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 21.730 60.360 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 21.300 60.360 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 20.870 60.360 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 20.440 60.360 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 20.010 60.360 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 19.580 60.360 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 19.150 60.360 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 18.720 60.360 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 18.290 60.360 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.160 17.860 60.360 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.895 91.385 60.215 91.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.895 90.955 60.215 91.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835 90.495 60.155 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835 90.065 60.155 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835 89.635 60.155 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835 89.205 60.155 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835 88.775 60.155 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.835 88.350 60.155 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 82.360 60.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 81.955 60.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 81.550 60.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 81.145 60.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 80.740 60.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 80.335 60.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 79.930 60.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 79.525 60.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 79.120 60.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 78.715 60.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 78.310 60.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 77.905 60.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 77.500 60.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 77.095 60.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 76.690 60.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 76.285 60.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 75.880 60.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 75.475 60.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 75.070 60.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 74.665 60.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 74.260 60.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 73.855 60.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 73.450 60.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 73.045 60.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 72.635 60.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 72.225 60.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 71.815 60.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 71.405 60.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 70.995 60.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 70.585 60.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 70.175 60.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 69.765 60.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 69.355 60.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 68.945 60.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 68.535 60.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.810 68.125 60.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 87.815 60.030 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 87.410 60.030 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 87.005 60.030 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 86.600 60.030 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 86.195 60.030 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 85.795 60.030 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 85.395 60.030 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 84.995 60.030 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 84.595 60.030 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 84.195 60.030 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 83.795 60.030 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 83.395 60.030 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.710 82.995 60.030 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 22.160 59.955 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 21.730 59.955 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 21.300 59.955 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 20.870 59.955 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 20.440 59.955 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 20.010 59.955 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 19.580 59.955 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 19.150 59.955 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 18.720 59.955 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 18.290 59.955 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.755 17.860 59.955 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 90.495 59.745 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 90.065 59.745 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 89.635 59.745 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 89.205 59.745 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 88.775 59.745 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 88.350 59.745 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 82.360 59.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 81.955 59.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 81.550 59.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 81.145 59.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 80.740 59.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 80.335 59.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 79.930 59.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 79.525 59.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 79.120 59.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 78.715 59.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 78.310 59.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 77.905 59.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 77.500 59.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 77.095 59.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 76.690 59.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 76.285 59.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 75.880 59.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 75.475 59.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 75.070 59.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 74.665 59.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 74.260 59.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 73.855 59.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 73.450 59.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 73.045 59.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 72.635 59.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 72.225 59.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 71.815 59.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 71.405 59.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 70.995 59.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 70.585 59.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 70.175 59.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 69.765 59.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 69.355 59.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 68.945 59.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 68.535 59.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.410 68.125 59.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 87.815 59.620 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 87.410 59.620 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 87.005 59.620 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 86.600 59.620 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 86.195 59.620 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 85.795 59.620 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 85.395 59.620 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 84.995 59.620 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 84.595 59.620 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 84.195 59.620 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 83.795 59.620 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 83.395 59.620 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.300 82.995 59.620 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 22.160 59.550 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 21.730 59.550 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 21.300 59.550 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 20.870 59.550 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 20.440 59.550 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 20.010 59.550 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 19.580 59.550 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 19.150 59.550 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 18.720 59.550 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 18.290 59.550 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.350 17.860 59.550 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 90.495 59.335 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 90.065 59.335 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 89.635 59.335 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 89.205 59.335 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 88.775 59.335 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 88.350 59.335 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 82.360 59.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 81.955 59.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 81.550 59.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 81.145 59.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 80.740 59.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 80.335 59.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 79.930 59.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 79.525 59.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 79.120 59.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 78.715 59.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 78.310 59.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 77.905 59.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 77.500 59.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 77.095 59.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 76.690 59.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 76.285 59.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 75.880 59.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 75.475 59.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 75.070 59.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 74.665 59.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 74.260 59.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 73.855 59.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 73.450 59.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 73.045 59.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 72.635 59.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 72.225 59.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 71.815 59.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 71.405 59.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 70.995 59.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 70.585 59.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 70.175 59.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 69.765 59.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 69.355 59.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 68.945 59.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 68.535 59.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.010 68.125 59.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 87.815 59.210 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 87.410 59.210 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 87.005 59.210 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 86.600 59.210 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 86.195 59.210 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 85.795 59.210 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 85.395 59.210 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 84.995 59.210 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 84.595 59.210 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 84.195 59.210 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 83.795 59.210 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 83.395 59.210 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.890 82.995 59.210 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 22.160 59.145 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 21.730 59.145 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 21.300 59.145 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 20.870 59.145 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 20.440 59.145 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 20.010 59.145 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 19.580 59.145 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 19.150 59.145 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 18.720 59.145 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 18.290 59.145 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.945 17.860 59.145 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 82.360 58.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 81.955 58.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 81.550 58.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 81.145 58.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 80.740 58.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 80.335 58.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 79.930 58.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 79.525 58.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 79.120 58.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 78.715 58.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 78.310 58.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 77.905 58.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 77.500 58.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 77.095 58.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 76.690 58.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 76.285 58.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 75.880 58.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 75.475 58.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 75.070 58.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 74.665 58.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 74.260 58.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 73.855 58.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 73.450 58.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 73.045 58.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 72.635 58.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 72.225 58.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 71.815 58.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 71.405 58.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 70.995 58.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 70.585 58.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 70.175 58.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 69.765 58.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 69.355 58.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 68.945 58.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 68.535 58.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 68.125 58.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.515 89.205 58.835 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.515 88.785 58.835 89.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.515 88.370 58.835 88.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 87.815 58.800 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 87.410 58.800 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 87.005 58.800 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 86.600 58.800 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 86.195 58.800 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 85.795 58.800 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 85.395 58.800 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 84.995 58.800 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 84.595 58.800 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 84.195 58.800 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 83.795 58.800 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 83.395 58.800 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.480 82.995 58.800 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 22.160 58.740 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 21.730 58.740 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 21.300 58.740 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 20.870 58.740 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 20.440 58.740 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 20.010 58.740 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 19.580 58.740 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 19.150 58.740 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 18.720 58.740 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 18.290 58.740 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.540 17.860 58.740 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 82.360 58.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 81.955 58.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 81.550 58.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 81.145 58.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 80.740 58.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 80.335 58.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 79.930 58.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 79.525 58.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 79.120 58.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 78.715 58.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 78.310 58.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 77.905 58.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 77.500 58.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 77.095 58.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 76.690 58.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 76.285 58.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 75.880 58.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 75.475 58.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 75.070 58.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 74.665 58.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 74.260 58.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 73.855 58.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 73.450 58.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 73.045 58.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 72.635 58.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 72.225 58.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 71.815 58.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 71.405 58.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 70.995 58.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 70.585 58.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 70.175 58.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 69.765 58.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 69.355 58.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 68.945 58.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 68.535 58.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 68.125 58.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 22.160 58.335 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 21.730 58.335 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 21.300 58.335 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 20.870 58.335 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 20.440 58.335 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 20.010 58.335 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 19.580 58.335 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 19.150 58.335 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 18.720 58.335 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 18.290 58.335 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.135 17.860 58.335 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 87.815 58.390 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 87.410 58.390 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 87.005 58.390 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 86.600 58.390 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 86.195 58.390 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 85.795 58.390 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 85.395 58.390 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 84.995 58.390 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 84.595 58.390 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 84.195 58.390 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 83.795 58.390 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 83.395 58.390 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.070 82.995 58.390 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 82.360 58.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 81.955 58.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 81.550 58.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 81.145 58.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 80.740 58.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 80.335 58.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 79.930 58.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 79.525 58.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 79.120 58.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 78.715 58.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 78.310 58.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 77.905 58.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 77.500 58.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 77.095 58.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 76.690 58.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 76.285 58.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 75.880 58.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 75.475 58.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 75.070 58.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 74.665 58.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 74.260 58.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 73.855 58.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 73.450 58.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 73.045 58.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 72.635 58.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 72.225 58.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 71.815 58.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 71.405 58.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 70.995 58.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 70.585 58.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 70.175 58.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 69.765 58.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 69.355 58.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 68.945 58.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 68.535 58.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.810 68.125 58.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.735 89.205 58.055 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.735 88.785 58.055 89.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.735 88.370 58.055 88.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 22.160 57.930 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 21.730 57.930 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 21.300 57.930 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 20.870 57.930 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 20.440 57.930 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 20.010 57.930 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 19.580 57.930 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 19.150 57.930 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 18.720 57.930 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 18.290 57.930 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.730 17.860 57.930 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 87.815 57.980 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 87.410 57.980 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 87.005 57.980 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 86.600 57.980 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 86.195 57.980 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 85.795 57.980 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 85.395 57.980 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 84.995 57.980 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 84.595 57.980 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 84.195 57.980 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 83.795 57.980 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 83.395 57.980 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.660 82.995 57.980 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 82.360 57.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 81.955 57.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 81.550 57.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 81.145 57.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 80.740 57.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 80.335 57.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 79.930 57.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 79.525 57.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 79.120 57.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 78.715 57.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 78.310 57.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 77.905 57.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 77.500 57.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 77.095 57.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 76.690 57.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 76.285 57.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 75.880 57.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 75.475 57.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 75.070 57.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 74.665 57.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 74.260 57.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 73.855 57.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 73.450 57.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 73.045 57.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 72.635 57.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 72.225 57.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 71.815 57.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 71.405 57.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 70.995 57.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 70.585 57.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 70.175 57.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 69.765 57.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 69.355 57.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 68.945 57.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 68.535 57.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.410 68.125 57.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 22.160 57.525 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 21.730 57.525 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 21.300 57.525 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 20.870 57.525 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 20.440 57.525 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 20.010 57.525 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 19.580 57.525 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 19.150 57.525 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 18.720 57.525 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 18.290 57.525 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.325 17.860 57.525 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 87.815 57.570 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 87.410 57.570 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 87.005 57.570 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 86.600 57.570 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 86.195 57.570 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 85.795 57.570 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 85.395 57.570 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 84.995 57.570 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 84.595 57.570 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 84.195 57.570 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 83.795 57.570 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 83.395 57.570 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.250 82.995 57.570 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 82.360 57.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 81.955 57.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 81.550 57.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 81.145 57.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 80.740 57.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 80.335 57.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 79.930 57.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 79.525 57.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 79.120 57.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 78.715 57.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 78.310 57.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 77.905 57.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 77.500 57.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 77.095 57.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 76.690 57.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 76.285 57.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 75.880 57.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 75.475 57.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 75.070 57.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 74.665 57.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 74.260 57.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 73.855 57.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 73.450 57.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 73.045 57.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 72.635 57.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 72.225 57.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 71.815 57.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 71.405 57.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 70.995 57.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 70.585 57.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 70.175 57.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 69.765 57.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 69.355 57.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 68.945 57.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 68.535 57.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.010 68.125 57.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 22.160 57.120 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 21.730 57.120 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 21.300 57.120 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 20.870 57.120 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 20.440 57.120 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 20.010 57.120 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 19.580 57.120 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 19.150 57.120 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 18.720 57.120 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 18.290 57.120 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.920 17.860 57.120 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 87.815 57.160 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 87.410 57.160 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 87.005 57.160 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 86.600 57.160 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 86.195 57.160 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 85.795 57.160 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 85.395 57.160 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 84.995 57.160 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 84.595 57.160 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 84.195 57.160 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 83.795 57.160 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 83.395 57.160 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.840 82.995 57.160 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 82.360 56.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 81.955 56.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 81.550 56.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 81.145 56.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 80.740 56.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 80.335 56.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 79.930 56.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 79.525 56.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 79.120 56.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 78.715 56.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 78.310 56.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 77.905 56.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 77.500 56.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 77.095 56.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 76.690 56.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 76.285 56.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 75.880 56.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 75.475 56.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 75.070 56.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 74.665 56.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 74.260 56.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 73.855 56.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 73.450 56.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 73.045 56.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 72.635 56.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 72.225 56.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 71.815 56.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 71.405 56.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 70.995 56.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 70.585 56.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 70.175 56.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 69.765 56.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 69.355 56.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 68.945 56.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 68.535 56.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.610 68.125 56.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 22.160 56.715 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 21.730 56.715 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 21.300 56.715 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 20.870 56.715 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 20.440 56.715 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 20.010 56.715 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 19.580 56.715 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 19.150 56.715 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 18.720 56.715 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 18.290 56.715 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.515 17.860 56.715 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 87.815 56.750 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 87.410 56.750 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 87.005 56.750 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 86.600 56.750 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 86.195 56.750 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 85.795 56.750 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 85.395 56.750 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 84.995 56.750 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 84.595 56.750 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 84.195 56.750 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 83.795 56.750 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 83.395 56.750 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.430 82.995 56.750 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 82.360 56.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 81.955 56.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 81.550 56.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 81.145 56.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 80.740 56.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 80.335 56.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 79.930 56.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 79.525 56.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 79.120 56.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 78.715 56.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 78.310 56.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 77.905 56.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 77.500 56.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 77.095 56.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 76.690 56.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 76.285 56.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 75.880 56.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 75.475 56.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 75.070 56.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 74.665 56.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 74.260 56.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 73.855 56.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 73.450 56.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 73.045 56.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 72.635 56.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 72.225 56.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 71.815 56.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 71.405 56.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 70.995 56.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 70.585 56.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 70.175 56.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 69.765 56.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 69.355 56.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 68.945 56.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 68.535 56.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.210 68.125 56.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 22.160 56.310 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 21.730 56.310 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 21.300 56.310 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 20.870 56.310 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 20.440 56.310 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 20.010 56.310 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 19.580 56.310 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 19.150 56.310 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 18.720 56.310 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 18.290 56.310 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.110 17.860 56.310 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.935 86.690 56.255 87.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.935 86.250 56.255 86.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.935 85.815 56.255 86.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 82.360 56.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 81.955 56.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 81.550 56.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 81.145 56.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 80.740 56.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 80.335 56.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 79.930 56.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 79.525 56.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 79.120 56.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 78.715 56.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 78.310 56.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 77.905 56.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 77.500 56.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 77.095 56.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 76.690 56.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 76.285 56.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 75.880 56.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 75.475 56.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 75.070 56.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 74.665 56.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 74.260 56.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 73.855 56.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 73.450 56.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 73.045 56.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 72.635 56.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 72.225 56.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 71.815 56.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 71.405 56.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 70.995 56.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 70.585 56.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 70.175 56.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 69.765 56.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 69.355 56.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 68.945 56.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 68.535 56.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.810 68.125 56.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 85.265 56.065 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 84.800 56.065 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 84.335 56.065 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 83.870 56.065 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 83.410 56.065 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 82.950 56.065 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 22.160 55.905 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 21.730 55.905 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 21.300 55.905 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 20.870 55.905 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 20.440 55.905 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 20.010 55.905 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 19.580 55.905 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 19.150 55.905 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 18.720 55.905 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 18.290 55.905 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.705 17.860 55.905 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 82.360 55.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 81.955 55.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 81.550 55.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 81.145 55.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 80.740 55.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 80.335 55.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 79.930 55.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 79.525 55.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 79.120 55.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 78.715 55.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 78.310 55.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 77.905 55.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 77.500 55.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 77.095 55.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 76.690 55.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 76.285 55.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 75.880 55.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 75.475 55.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 75.070 55.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 74.665 55.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 74.260 55.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 73.855 55.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 73.450 55.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 73.045 55.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 72.635 55.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 72.225 55.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 71.815 55.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 71.405 55.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 70.995 55.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 70.585 55.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 70.175 55.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 69.765 55.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 69.355 55.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 68.945 55.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 68.535 55.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.410 68.125 55.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265 85.265 55.585 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265 84.800 55.585 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265 84.335 55.585 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265 83.870 55.585 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265 83.410 55.585 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.265 82.950 55.585 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 22.160 55.500 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 21.730 55.500 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 21.300 55.500 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 20.870 55.500 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 20.440 55.500 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 20.010 55.500 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 19.580 55.500 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 19.150 55.500 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 18.720 55.500 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 18.290 55.500 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.300 17.860 55.500 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.195 86.690 55.515 87.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.195 86.250 55.515 86.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.195 85.815 55.515 86.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 82.360 55.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 81.955 55.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 81.550 55.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 81.145 55.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 80.740 55.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 80.335 55.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 79.930 55.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 79.525 55.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 79.120 55.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 78.715 55.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 78.310 55.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 77.905 55.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 77.500 55.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 77.095 55.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 76.690 55.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 76.285 55.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 75.880 55.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 75.475 55.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 75.070 55.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 74.665 55.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 74.260 55.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 73.855 55.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 73.450 55.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 73.045 55.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 72.635 55.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 72.225 55.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 71.815 55.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 71.405 55.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 70.995 55.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 70.585 55.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 70.175 55.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 69.765 55.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 69.355 55.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 68.945 55.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 68.535 55.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.010 68.125 55.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 22.160 55.095 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 21.730 55.095 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 21.300 55.095 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 20.870 55.095 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 20.440 55.095 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 20.010 55.095 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 19.580 55.095 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 19.150 55.095 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 18.720 55.095 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 18.290 55.095 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.895 17.860 55.095 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785 85.265 55.105 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785 84.800 55.105 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785 84.335 55.105 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785 83.870 55.105 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785 83.410 55.105 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.785 82.950 55.105 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 82.360 54.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 81.955 54.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 81.550 54.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 81.145 54.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 80.740 54.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 80.335 54.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 79.930 54.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 79.525 54.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 79.120 54.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 78.715 54.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 78.310 54.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 77.905 54.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 77.500 54.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 77.095 54.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 76.690 54.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 76.285 54.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 75.880 54.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 75.475 54.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 75.070 54.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 74.665 54.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 74.260 54.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 73.855 54.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 73.450 54.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 73.045 54.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 72.635 54.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 72.225 54.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 71.815 54.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 71.405 54.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 70.995 54.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 70.585 54.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 70.175 54.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 69.765 54.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 69.355 54.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 68.945 54.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 68.535 54.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.610 68.125 54.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 22.160 54.690 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 21.730 54.690 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 21.300 54.690 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 20.870 54.690 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 20.440 54.690 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 20.010 54.690 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 19.580 54.690 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 19.150 54.690 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 18.720 54.690 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 18.290 54.690 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.490 17.860 54.690 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305 85.265 54.625 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305 84.800 54.625 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305 84.335 54.625 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305 83.870 54.625 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305 83.410 54.625 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.305 82.950 54.625 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 82.360 54.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 81.955 54.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 81.550 54.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 81.145 54.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 80.740 54.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 80.335 54.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 79.930 54.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 79.525 54.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 79.120 54.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 78.715 54.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 78.310 54.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 77.905 54.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 77.500 54.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 77.095 54.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 76.690 54.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 76.285 54.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 75.880 54.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 75.475 54.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 75.070 54.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 74.665 54.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 74.260 54.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 73.855 54.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 73.450 54.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 73.045 54.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 72.635 54.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 72.225 54.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 71.815 54.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 71.405 54.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 70.995 54.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 70.585 54.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 70.175 54.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 69.765 54.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 69.355 54.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 68.945 54.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 68.535 54.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.210 68.125 54.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 22.160 54.285 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 21.730 54.285 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 21.300 54.285 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 20.870 54.285 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 20.440 54.285 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 20.010 54.285 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 19.580 54.285 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 19.150 54.285 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 18.720 54.285 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 18.290 54.285 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.085 17.860 54.285 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825 85.265 54.145 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825 84.800 54.145 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825 84.335 54.145 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825 83.870 54.145 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825 83.410 54.145 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.825 82.950 54.145 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 82.360 54.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 81.955 54.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 81.550 54.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 81.145 54.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 80.740 54.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 80.335 54.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 79.930 54.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 79.525 54.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 79.120 54.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 78.715 54.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 78.310 54.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 77.905 54.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 77.500 54.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 77.095 54.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 76.690 54.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 76.285 54.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 75.880 54.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 75.475 54.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 75.070 54.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 74.665 54.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 74.260 54.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 73.855 54.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 73.450 54.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 73.045 54.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 72.635 54.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 72.225 54.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 71.815 54.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 71.405 54.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 70.995 54.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 70.585 54.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 70.175 54.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 69.765 54.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 69.355 54.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 68.945 54.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 68.535 54.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.810 68.125 54.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 22.160 53.880 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 21.730 53.880 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 21.300 53.880 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 20.870 53.880 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 20.440 53.880 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 20.010 53.880 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 19.580 53.880 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 19.150 53.880 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 18.720 53.880 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 18.290 53.880 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.680 17.860 53.880 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 82.360 53.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 81.955 53.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 81.550 53.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 81.145 53.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 80.740 53.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 80.335 53.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 79.930 53.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 79.525 53.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 79.120 53.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 78.715 53.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 78.310 53.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 77.905 53.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 77.500 53.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 77.095 53.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 76.690 53.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 76.285 53.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 75.880 53.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 75.475 53.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 75.070 53.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 74.665 53.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 74.260 53.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 73.855 53.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 73.450 53.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 73.045 53.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 72.635 53.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 72.225 53.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 71.815 53.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 71.405 53.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 70.995 53.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 70.585 53.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 70.175 53.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 69.765 53.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 69.355 53.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 68.945 53.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 68.535 53.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.410 68.125 53.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.280 83.960 53.600 84.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.280 83.410 53.600 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.280 82.860 53.600 83.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 22.160 53.475 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 21.730 53.475 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 21.300 53.475 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 20.870 53.475 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 20.440 53.475 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 20.010 53.475 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 19.580 53.475 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 19.150 53.475 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 18.720 53.475 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 18.290 53.475 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.275 17.860 53.475 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 82.360 53.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 81.955 53.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 81.550 53.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 81.145 53.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 80.740 53.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 80.335 53.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 79.930 53.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 79.525 53.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 79.120 53.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 78.715 53.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 78.310 53.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 77.905 53.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 77.500 53.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 77.095 53.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 76.690 53.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 76.285 53.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 75.880 53.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 75.475 53.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 75.070 53.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 74.665 53.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 74.260 53.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 73.855 53.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 73.450 53.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 73.045 53.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 72.635 53.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 72.225 53.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 71.815 53.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 71.405 53.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 70.995 53.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 70.585 53.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 70.175 53.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 69.765 53.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 69.355 53.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 68.945 53.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 68.535 53.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.010 68.125 53.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 22.160 53.070 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 21.730 53.070 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 21.300 53.070 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 20.870 53.070 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 20.440 53.070 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 20.010 53.070 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 19.580 53.070 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 19.150 53.070 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 18.720 53.070 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 18.290 53.070 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.870 17.860 53.070 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 82.360 52.810 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 81.955 52.810 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 81.550 52.810 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 81.145 52.810 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 80.740 52.810 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 80.335 52.810 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 79.930 52.810 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 79.525 52.810 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 79.120 52.810 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 78.715 52.810 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 78.310 52.810 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 77.905 52.810 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 77.500 52.810 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 77.095 52.810 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 76.690 52.810 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 76.285 52.810 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 75.880 52.810 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 75.475 52.810 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 75.070 52.810 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 74.665 52.810 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 74.260 52.810 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 73.855 52.810 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 73.450 52.810 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 73.045 52.810 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 72.635 52.810 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 72.225 52.810 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 71.815 52.810 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 71.405 52.810 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 70.995 52.810 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 70.585 52.810 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 70.175 52.810 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 69.765 52.810 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 69.355 52.810 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 68.945 52.810 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 68.535 52.810 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.610 68.125 52.810 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490 83.960 52.810 84.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490 83.410 52.810 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.490 82.860 52.810 83.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 22.160 52.665 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 21.730 52.665 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 21.300 52.665 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 20.870 52.665 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 20.440 52.665 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 20.010 52.665 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 19.580 52.665 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 19.150 52.665 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 18.720 52.665 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 18.290 52.665 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.465 17.860 52.665 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 82.360 52.410 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 81.955 52.410 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 81.550 52.410 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 81.145 52.410 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 80.740 52.410 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 80.335 52.410 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 79.930 52.410 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 79.525 52.410 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 79.120 52.410 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 78.715 52.410 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 78.310 52.410 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 77.905 52.410 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 77.500 52.410 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 77.095 52.410 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 76.690 52.410 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 76.285 52.410 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 75.880 52.410 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 75.475 52.410 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 75.070 52.410 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 74.665 52.410 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 74.260 52.410 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 73.855 52.410 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 73.450 52.410 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 73.045 52.410 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 72.635 52.410 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 72.225 52.410 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 71.815 52.410 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 71.405 52.410 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 70.995 52.410 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 70.585 52.410 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 70.175 52.410 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 69.765 52.410 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 69.355 52.410 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 68.945 52.410 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 68.535 52.410 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.210 68.125 52.410 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 22.160 52.260 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 21.730 52.260 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 21.300 52.260 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 20.870 52.260 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 20.440 52.260 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 20.010 52.260 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 19.580 52.260 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 19.150 52.260 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 18.720 52.260 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 18.290 52.260 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 17.860 52.260 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 82.360 52.010 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 81.955 52.010 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 81.550 52.010 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 81.145 52.010 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 80.740 52.010 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 80.335 52.010 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 79.930 52.010 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 79.525 52.010 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 79.120 52.010 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 78.715 52.010 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 78.310 52.010 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 77.905 52.010 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 77.500 52.010 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 77.095 52.010 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 76.690 52.010 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 76.285 52.010 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 75.880 52.010 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 75.475 52.010 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 75.070 52.010 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 74.665 52.010 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 74.260 52.010 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 73.855 52.010 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 73.450 52.010 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 73.045 52.010 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 72.635 52.010 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 72.225 52.010 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 71.815 52.010 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 71.405 52.010 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 70.995 52.010 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 70.585 52.010 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 70.175 52.010 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 69.765 52.010 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 69.355 52.010 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 68.945 52.010 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 68.535 52.010 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.810 68.125 52.010 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 22.160 51.855 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 21.730 51.855 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 21.300 51.855 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 20.870 51.855 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 20.440 51.855 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 20.010 51.855 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 19.580 51.855 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 19.150 51.855 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 18.720 51.855 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 18.290 51.855 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.655 17.860 51.855 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 82.360 51.610 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 81.955 51.610 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 81.550 51.610 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 81.145 51.610 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 80.740 51.610 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 80.335 51.610 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 79.930 51.610 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 79.525 51.610 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 79.120 51.610 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 78.715 51.610 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 78.310 51.610 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 77.905 51.610 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 77.500 51.610 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 77.095 51.610 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 76.690 51.610 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 76.285 51.610 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 75.880 51.610 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 75.475 51.610 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 75.070 51.610 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 74.665 51.610 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 74.260 51.610 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 73.855 51.610 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 73.450 51.610 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 73.045 51.610 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 72.635 51.610 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 72.225 51.610 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 71.815 51.610 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 71.405 51.610 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 70.995 51.610 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 70.585 51.610 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 70.175 51.610 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 69.765 51.610 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 69.355 51.610 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 68.945 51.610 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 68.535 51.610 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.410 68.125 51.610 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 22.160 51.450 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 21.730 51.450 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 21.300 51.450 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 20.870 51.450 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 20.440 51.450 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 20.010 51.450 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 19.580 51.450 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 19.150 51.450 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 18.720 51.450 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 18.290 51.450 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.250 17.860 51.450 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 82.360 51.210 82.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 81.955 51.210 82.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 81.550 51.210 81.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 81.145 51.210 81.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 80.740 51.210 80.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 80.335 51.210 80.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 79.930 51.210 80.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 79.525 51.210 79.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 79.120 51.210 79.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 78.715 51.210 78.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 78.310 51.210 78.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 77.905 51.210 78.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 77.500 51.210 77.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 77.095 51.210 77.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 76.690 51.210 76.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 76.285 51.210 76.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 75.880 51.210 76.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 75.475 51.210 75.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 75.070 51.210 75.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 74.665 51.210 74.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 74.260 51.210 74.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 73.855 51.210 74.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 73.450 51.210 73.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 73.045 51.210 73.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 72.635 51.210 72.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 72.225 51.210 72.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 71.815 51.210 72.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 71.405 51.210 71.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 70.995 51.210 71.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 70.585 51.210 70.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 70.175 51.210 70.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 69.765 51.210 69.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 69.355 51.210 69.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 68.945 51.210 69.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 68.535 51.210 68.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.010 68.125 51.210 68.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 22.160 51.045 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 21.730 51.045 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 21.300 51.045 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 20.870 51.045 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 20.440 51.045 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 20.010 51.045 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 19.580 51.045 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 19.150 51.045 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 18.720 51.045 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 18.290 51.045 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 17.860 51.045 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 22.160 24.410 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 21.730 24.410 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 21.300 24.410 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 20.870 24.410 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 20.440 24.410 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 20.010 24.410 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 19.580 24.410 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 19.150 24.410 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 18.720 24.410 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 18.290 24.410 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.210 17.860 24.410 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 82.300 24.305 82.620 ;
      LAYER met4 ;
        RECT 23.985 82.300 24.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 81.895 24.305 82.215 ;
      LAYER met4 ;
        RECT 23.985 81.895 24.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 81.490 24.305 81.810 ;
      LAYER met4 ;
        RECT 23.985 81.490 24.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 81.085 24.305 81.405 ;
      LAYER met4 ;
        RECT 23.985 81.085 24.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 80.680 24.305 81.000 ;
      LAYER met4 ;
        RECT 23.985 80.680 24.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 80.275 24.305 80.595 ;
      LAYER met4 ;
        RECT 23.985 80.275 24.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 79.870 24.305 80.190 ;
      LAYER met4 ;
        RECT 23.985 79.870 24.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 79.465 24.305 79.785 ;
      LAYER met4 ;
        RECT 23.985 79.465 24.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 79.060 24.305 79.380 ;
      LAYER met4 ;
        RECT 23.985 79.060 24.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 78.655 24.305 78.975 ;
      LAYER met4 ;
        RECT 23.985 78.655 24.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 78.250 24.305 78.570 ;
      LAYER met4 ;
        RECT 23.985 78.250 24.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 77.845 24.305 78.165 ;
      LAYER met4 ;
        RECT 23.985 77.845 24.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 77.440 24.305 77.760 ;
      LAYER met4 ;
        RECT 23.985 77.440 24.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 77.035 24.305 77.355 ;
      LAYER met4 ;
        RECT 23.985 77.035 24.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 76.630 24.305 76.950 ;
      LAYER met4 ;
        RECT 23.985 76.630 24.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 76.225 24.305 76.545 ;
      LAYER met4 ;
        RECT 23.985 76.225 24.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 75.820 24.305 76.140 ;
      LAYER met4 ;
        RECT 23.985 75.820 24.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 75.415 24.305 75.735 ;
      LAYER met4 ;
        RECT 23.985 75.415 24.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 75.010 24.305 75.330 ;
      LAYER met4 ;
        RECT 23.985 75.010 24.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 74.605 24.305 74.925 ;
      LAYER met4 ;
        RECT 23.985 74.605 24.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 74.200 24.305 74.520 ;
      LAYER met4 ;
        RECT 23.985 74.200 24.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 73.795 24.305 74.115 ;
      LAYER met4 ;
        RECT 23.985 73.795 24.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 73.390 24.305 73.710 ;
      LAYER met4 ;
        RECT 23.985 73.390 24.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 72.985 24.305 73.305 ;
      LAYER met4 ;
        RECT 23.985 72.985 24.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 72.575 24.305 72.895 ;
      LAYER met4 ;
        RECT 23.985 72.575 24.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 72.165 24.305 72.485 ;
      LAYER met4 ;
        RECT 23.985 72.165 24.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 71.755 24.305 72.075 ;
      LAYER met4 ;
        RECT 23.985 71.755 24.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 71.345 24.305 71.665 ;
      LAYER met4 ;
        RECT 23.985 71.345 24.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 70.935 24.305 71.255 ;
      LAYER met4 ;
        RECT 23.985 70.935 24.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 70.525 24.305 70.845 ;
      LAYER met4 ;
        RECT 23.985 70.525 24.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 70.115 24.305 70.435 ;
      LAYER met4 ;
        RECT 23.985 70.115 24.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 69.705 24.305 70.025 ;
      LAYER met4 ;
        RECT 23.985 69.705 24.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 69.295 24.305 69.615 ;
      LAYER met4 ;
        RECT 23.985 69.295 24.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 68.885 24.305 69.205 ;
      LAYER met4 ;
        RECT 23.985 68.885 24.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 68.475 24.305 68.795 ;
      LAYER met4 ;
        RECT 23.985 68.475 24.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.985 68.065 24.305 68.385 ;
      LAYER met4 ;
        RECT 23.985 68.065 24.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 22.160 24.000 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 21.730 24.000 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 21.300 24.000 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 20.870 24.000 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 20.440 24.000 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 20.010 24.000 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 19.580 24.000 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 19.150 24.000 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 18.720 24.000 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 18.290 24.000 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.800 17.860 24.000 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 82.300 23.905 82.620 ;
      LAYER met4 ;
        RECT 23.585 82.300 23.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 81.895 23.905 82.215 ;
      LAYER met4 ;
        RECT 23.585 81.895 23.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 81.490 23.905 81.810 ;
      LAYER met4 ;
        RECT 23.585 81.490 23.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 81.085 23.905 81.405 ;
      LAYER met4 ;
        RECT 23.585 81.085 23.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 80.680 23.905 81.000 ;
      LAYER met4 ;
        RECT 23.585 80.680 23.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 80.275 23.905 80.595 ;
      LAYER met4 ;
        RECT 23.585 80.275 23.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 79.870 23.905 80.190 ;
      LAYER met4 ;
        RECT 23.585 79.870 23.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 79.465 23.905 79.785 ;
      LAYER met4 ;
        RECT 23.585 79.465 23.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 79.060 23.905 79.380 ;
      LAYER met4 ;
        RECT 23.585 79.060 23.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 78.655 23.905 78.975 ;
      LAYER met4 ;
        RECT 23.585 78.655 23.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 78.250 23.905 78.570 ;
      LAYER met4 ;
        RECT 23.585 78.250 23.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 77.845 23.905 78.165 ;
      LAYER met4 ;
        RECT 23.585 77.845 23.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 77.440 23.905 77.760 ;
      LAYER met4 ;
        RECT 23.585 77.440 23.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 77.035 23.905 77.355 ;
      LAYER met4 ;
        RECT 23.585 77.035 23.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 76.630 23.905 76.950 ;
      LAYER met4 ;
        RECT 23.585 76.630 23.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 76.225 23.905 76.545 ;
      LAYER met4 ;
        RECT 23.585 76.225 23.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 75.820 23.905 76.140 ;
      LAYER met4 ;
        RECT 23.585 75.820 23.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 75.415 23.905 75.735 ;
      LAYER met4 ;
        RECT 23.585 75.415 23.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 75.010 23.905 75.330 ;
      LAYER met4 ;
        RECT 23.585 75.010 23.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 74.605 23.905 74.925 ;
      LAYER met4 ;
        RECT 23.585 74.605 23.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 74.200 23.905 74.520 ;
      LAYER met4 ;
        RECT 23.585 74.200 23.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 73.795 23.905 74.115 ;
      LAYER met4 ;
        RECT 23.585 73.795 23.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 73.390 23.905 73.710 ;
      LAYER met4 ;
        RECT 23.585 73.390 23.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 72.985 23.905 73.305 ;
      LAYER met4 ;
        RECT 23.585 72.985 23.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 72.575 23.905 72.895 ;
      LAYER met4 ;
        RECT 23.585 72.575 23.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 72.165 23.905 72.485 ;
      LAYER met4 ;
        RECT 23.585 72.165 23.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 71.755 23.905 72.075 ;
      LAYER met4 ;
        RECT 23.585 71.755 23.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 71.345 23.905 71.665 ;
      LAYER met4 ;
        RECT 23.585 71.345 23.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 70.935 23.905 71.255 ;
      LAYER met4 ;
        RECT 23.585 70.935 23.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 70.525 23.905 70.845 ;
      LAYER met4 ;
        RECT 23.585 70.525 23.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 70.115 23.905 70.435 ;
      LAYER met4 ;
        RECT 23.585 70.115 23.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 69.705 23.905 70.025 ;
      LAYER met4 ;
        RECT 23.585 69.705 23.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 69.295 23.905 69.615 ;
      LAYER met4 ;
        RECT 23.585 69.295 23.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 68.885 23.905 69.205 ;
      LAYER met4 ;
        RECT 23.585 68.885 23.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 68.475 23.905 68.795 ;
      LAYER met4 ;
        RECT 23.585 68.475 23.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.585 68.065 23.905 68.385 ;
      LAYER met4 ;
        RECT 23.585 68.065 23.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 22.160 23.590 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 21.730 23.590 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 21.300 23.590 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 20.870 23.590 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 20.440 23.590 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 20.010 23.590 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 19.580 23.590 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 19.150 23.590 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 18.720 23.590 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 18.290 23.590 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.390 17.860 23.590 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 82.300 23.505 82.620 ;
      LAYER met4 ;
        RECT 23.185 82.300 23.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 81.895 23.505 82.215 ;
      LAYER met4 ;
        RECT 23.185 81.895 23.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 81.490 23.505 81.810 ;
      LAYER met4 ;
        RECT 23.185 81.490 23.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 81.085 23.505 81.405 ;
      LAYER met4 ;
        RECT 23.185 81.085 23.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 80.680 23.505 81.000 ;
      LAYER met4 ;
        RECT 23.185 80.680 23.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 80.275 23.505 80.595 ;
      LAYER met4 ;
        RECT 23.185 80.275 23.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 79.870 23.505 80.190 ;
      LAYER met4 ;
        RECT 23.185 79.870 23.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 79.465 23.505 79.785 ;
      LAYER met4 ;
        RECT 23.185 79.465 23.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 79.060 23.505 79.380 ;
      LAYER met4 ;
        RECT 23.185 79.060 23.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 78.655 23.505 78.975 ;
      LAYER met4 ;
        RECT 23.185 78.655 23.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 78.250 23.505 78.570 ;
      LAYER met4 ;
        RECT 23.185 78.250 23.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 77.845 23.505 78.165 ;
      LAYER met4 ;
        RECT 23.185 77.845 23.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 77.440 23.505 77.760 ;
      LAYER met4 ;
        RECT 23.185 77.440 23.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 77.035 23.505 77.355 ;
      LAYER met4 ;
        RECT 23.185 77.035 23.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 76.630 23.505 76.950 ;
      LAYER met4 ;
        RECT 23.185 76.630 23.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 76.225 23.505 76.545 ;
      LAYER met4 ;
        RECT 23.185 76.225 23.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 75.820 23.505 76.140 ;
      LAYER met4 ;
        RECT 23.185 75.820 23.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 75.415 23.505 75.735 ;
      LAYER met4 ;
        RECT 23.185 75.415 23.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 75.010 23.505 75.330 ;
      LAYER met4 ;
        RECT 23.185 75.010 23.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 74.605 23.505 74.925 ;
      LAYER met4 ;
        RECT 23.185 74.605 23.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 74.200 23.505 74.520 ;
      LAYER met4 ;
        RECT 23.185 74.200 23.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 73.795 23.505 74.115 ;
      LAYER met4 ;
        RECT 23.185 73.795 23.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 73.390 23.505 73.710 ;
      LAYER met4 ;
        RECT 23.185 73.390 23.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 72.985 23.505 73.305 ;
      LAYER met4 ;
        RECT 23.185 72.985 23.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 72.575 23.505 72.895 ;
      LAYER met4 ;
        RECT 23.185 72.575 23.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 72.165 23.505 72.485 ;
      LAYER met4 ;
        RECT 23.185 72.165 23.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 71.755 23.505 72.075 ;
      LAYER met4 ;
        RECT 23.185 71.755 23.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 71.345 23.505 71.665 ;
      LAYER met4 ;
        RECT 23.185 71.345 23.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 70.935 23.505 71.255 ;
      LAYER met4 ;
        RECT 23.185 70.935 23.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 70.525 23.505 70.845 ;
      LAYER met4 ;
        RECT 23.185 70.525 23.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 70.115 23.505 70.435 ;
      LAYER met4 ;
        RECT 23.185 70.115 23.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 69.705 23.505 70.025 ;
      LAYER met4 ;
        RECT 23.185 69.705 23.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 69.295 23.505 69.615 ;
      LAYER met4 ;
        RECT 23.185 69.295 23.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 68.885 23.505 69.205 ;
      LAYER met4 ;
        RECT 23.185 68.885 23.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 68.475 23.505 68.795 ;
      LAYER met4 ;
        RECT 23.185 68.475 23.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.185 68.065 23.505 68.385 ;
      LAYER met4 ;
        RECT 23.185 68.065 23.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 22.160 23.180 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 21.730 23.180 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 21.300 23.180 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 20.870 23.180 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 20.440 23.180 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 20.010 23.180 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 19.580 23.180 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 19.150 23.180 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 18.720 23.180 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 18.290 23.180 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.980 17.860 23.180 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 82.300 23.105 82.620 ;
      LAYER met4 ;
        RECT 22.785 82.300 23.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 81.895 23.105 82.215 ;
      LAYER met4 ;
        RECT 22.785 81.895 23.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 81.490 23.105 81.810 ;
      LAYER met4 ;
        RECT 22.785 81.490 23.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 81.085 23.105 81.405 ;
      LAYER met4 ;
        RECT 22.785 81.085 23.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 80.680 23.105 81.000 ;
      LAYER met4 ;
        RECT 22.785 80.680 23.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 80.275 23.105 80.595 ;
      LAYER met4 ;
        RECT 22.785 80.275 23.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 79.870 23.105 80.190 ;
      LAYER met4 ;
        RECT 22.785 79.870 23.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 79.465 23.105 79.785 ;
      LAYER met4 ;
        RECT 22.785 79.465 23.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 79.060 23.105 79.380 ;
      LAYER met4 ;
        RECT 22.785 79.060 23.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 78.655 23.105 78.975 ;
      LAYER met4 ;
        RECT 22.785 78.655 23.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 78.250 23.105 78.570 ;
      LAYER met4 ;
        RECT 22.785 78.250 23.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 77.845 23.105 78.165 ;
      LAYER met4 ;
        RECT 22.785 77.845 23.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 77.440 23.105 77.760 ;
      LAYER met4 ;
        RECT 22.785 77.440 23.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 77.035 23.105 77.355 ;
      LAYER met4 ;
        RECT 22.785 77.035 23.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 76.630 23.105 76.950 ;
      LAYER met4 ;
        RECT 22.785 76.630 23.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 76.225 23.105 76.545 ;
      LAYER met4 ;
        RECT 22.785 76.225 23.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 75.820 23.105 76.140 ;
      LAYER met4 ;
        RECT 22.785 75.820 23.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 75.415 23.105 75.735 ;
      LAYER met4 ;
        RECT 22.785 75.415 23.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 75.010 23.105 75.330 ;
      LAYER met4 ;
        RECT 22.785 75.010 23.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 74.605 23.105 74.925 ;
      LAYER met4 ;
        RECT 22.785 74.605 23.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 74.200 23.105 74.520 ;
      LAYER met4 ;
        RECT 22.785 74.200 23.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 73.795 23.105 74.115 ;
      LAYER met4 ;
        RECT 22.785 73.795 23.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 73.390 23.105 73.710 ;
      LAYER met4 ;
        RECT 22.785 73.390 23.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 72.985 23.105 73.305 ;
      LAYER met4 ;
        RECT 22.785 72.985 23.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 72.575 23.105 72.895 ;
      LAYER met4 ;
        RECT 22.785 72.575 23.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 72.165 23.105 72.485 ;
      LAYER met4 ;
        RECT 22.785 72.165 23.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 71.755 23.105 72.075 ;
      LAYER met4 ;
        RECT 22.785 71.755 23.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 71.345 23.105 71.665 ;
      LAYER met4 ;
        RECT 22.785 71.345 23.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 70.935 23.105 71.255 ;
      LAYER met4 ;
        RECT 22.785 70.935 23.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 70.525 23.105 70.845 ;
      LAYER met4 ;
        RECT 22.785 70.525 23.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 70.115 23.105 70.435 ;
      LAYER met4 ;
        RECT 22.785 70.115 23.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 69.705 23.105 70.025 ;
      LAYER met4 ;
        RECT 22.785 69.705 23.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 69.295 23.105 69.615 ;
      LAYER met4 ;
        RECT 22.785 69.295 23.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 68.885 23.105 69.205 ;
      LAYER met4 ;
        RECT 22.785 68.885 23.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 68.475 23.105 68.795 ;
      LAYER met4 ;
        RECT 22.785 68.475 23.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.785 68.065 23.105 68.385 ;
      LAYER met4 ;
        RECT 22.785 68.065 23.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 22.160 22.770 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 21.730 22.770 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 21.300 22.770 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 20.870 22.770 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 20.440 22.770 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 20.010 22.770 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 19.580 22.770 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 19.150 22.770 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 18.720 22.770 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 18.290 22.770 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.570 17.860 22.770 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 83.960 22.765 84.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 83.410 22.765 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 82.860 22.765 83.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 82.300 22.705 82.620 ;
      LAYER met4 ;
        RECT 22.385 82.300 22.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 81.895 22.705 82.215 ;
      LAYER met4 ;
        RECT 22.385 81.895 22.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 81.490 22.705 81.810 ;
      LAYER met4 ;
        RECT 22.385 81.490 22.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 81.085 22.705 81.405 ;
      LAYER met4 ;
        RECT 22.385 81.085 22.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 80.680 22.705 81.000 ;
      LAYER met4 ;
        RECT 22.385 80.680 22.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 80.275 22.705 80.595 ;
      LAYER met4 ;
        RECT 22.385 80.275 22.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 79.870 22.705 80.190 ;
      LAYER met4 ;
        RECT 22.385 79.870 22.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 79.465 22.705 79.785 ;
      LAYER met4 ;
        RECT 22.385 79.465 22.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 79.060 22.705 79.380 ;
      LAYER met4 ;
        RECT 22.385 79.060 22.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 78.655 22.705 78.975 ;
      LAYER met4 ;
        RECT 22.385 78.655 22.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 78.250 22.705 78.570 ;
      LAYER met4 ;
        RECT 22.385 78.250 22.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 77.845 22.705 78.165 ;
      LAYER met4 ;
        RECT 22.385 77.845 22.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 77.440 22.705 77.760 ;
      LAYER met4 ;
        RECT 22.385 77.440 22.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 77.035 22.705 77.355 ;
      LAYER met4 ;
        RECT 22.385 77.035 22.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 76.630 22.705 76.950 ;
      LAYER met4 ;
        RECT 22.385 76.630 22.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 76.225 22.705 76.545 ;
      LAYER met4 ;
        RECT 22.385 76.225 22.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 75.820 22.705 76.140 ;
      LAYER met4 ;
        RECT 22.385 75.820 22.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 75.415 22.705 75.735 ;
      LAYER met4 ;
        RECT 22.385 75.415 22.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 75.010 22.705 75.330 ;
      LAYER met4 ;
        RECT 22.385 75.010 22.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 74.605 22.705 74.925 ;
      LAYER met4 ;
        RECT 22.385 74.605 22.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 74.200 22.705 74.520 ;
      LAYER met4 ;
        RECT 22.385 74.200 22.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 73.795 22.705 74.115 ;
      LAYER met4 ;
        RECT 22.385 73.795 22.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 73.390 22.705 73.710 ;
      LAYER met4 ;
        RECT 22.385 73.390 22.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 72.985 22.705 73.305 ;
      LAYER met4 ;
        RECT 22.385 72.985 22.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 72.575 22.705 72.895 ;
      LAYER met4 ;
        RECT 22.385 72.575 22.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 72.165 22.705 72.485 ;
      LAYER met4 ;
        RECT 22.385 72.165 22.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 71.755 22.705 72.075 ;
      LAYER met4 ;
        RECT 22.385 71.755 22.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 71.345 22.705 71.665 ;
      LAYER met4 ;
        RECT 22.385 71.345 22.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 70.935 22.705 71.255 ;
      LAYER met4 ;
        RECT 22.385 70.935 22.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 70.525 22.705 70.845 ;
      LAYER met4 ;
        RECT 22.385 70.525 22.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 70.115 22.705 70.435 ;
      LAYER met4 ;
        RECT 22.385 70.115 22.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 69.705 22.705 70.025 ;
      LAYER met4 ;
        RECT 22.385 69.705 22.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 69.295 22.705 69.615 ;
      LAYER met4 ;
        RECT 22.385 69.295 22.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 68.885 22.705 69.205 ;
      LAYER met4 ;
        RECT 22.385 68.885 22.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 68.475 22.705 68.795 ;
      LAYER met4 ;
        RECT 22.385 68.475 22.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.385 68.065 22.705 68.385 ;
      LAYER met4 ;
        RECT 22.385 68.065 22.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 22.160 22.360 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 21.730 22.360 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 21.300 22.360 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 20.870 22.360 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 20.440 22.360 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 20.010 22.360 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 19.580 22.360 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 19.150 22.360 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 18.720 22.360 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 18.290 22.360 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.160 17.860 22.360 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 82.300 22.305 82.620 ;
      LAYER met4 ;
        RECT 21.985 82.300 22.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 81.895 22.305 82.215 ;
      LAYER met4 ;
        RECT 21.985 81.895 22.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 81.490 22.305 81.810 ;
      LAYER met4 ;
        RECT 21.985 81.490 22.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 81.085 22.305 81.405 ;
      LAYER met4 ;
        RECT 21.985 81.085 22.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 80.680 22.305 81.000 ;
      LAYER met4 ;
        RECT 21.985 80.680 22.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 80.275 22.305 80.595 ;
      LAYER met4 ;
        RECT 21.985 80.275 22.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 79.870 22.305 80.190 ;
      LAYER met4 ;
        RECT 21.985 79.870 22.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 79.465 22.305 79.785 ;
      LAYER met4 ;
        RECT 21.985 79.465 22.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 79.060 22.305 79.380 ;
      LAYER met4 ;
        RECT 21.985 79.060 22.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 78.655 22.305 78.975 ;
      LAYER met4 ;
        RECT 21.985 78.655 22.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 78.250 22.305 78.570 ;
      LAYER met4 ;
        RECT 21.985 78.250 22.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 77.845 22.305 78.165 ;
      LAYER met4 ;
        RECT 21.985 77.845 22.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 77.440 22.305 77.760 ;
      LAYER met4 ;
        RECT 21.985 77.440 22.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 77.035 22.305 77.355 ;
      LAYER met4 ;
        RECT 21.985 77.035 22.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 76.630 22.305 76.950 ;
      LAYER met4 ;
        RECT 21.985 76.630 22.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 76.225 22.305 76.545 ;
      LAYER met4 ;
        RECT 21.985 76.225 22.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 75.820 22.305 76.140 ;
      LAYER met4 ;
        RECT 21.985 75.820 22.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 75.415 22.305 75.735 ;
      LAYER met4 ;
        RECT 21.985 75.415 22.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 75.010 22.305 75.330 ;
      LAYER met4 ;
        RECT 21.985 75.010 22.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 74.605 22.305 74.925 ;
      LAYER met4 ;
        RECT 21.985 74.605 22.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 74.200 22.305 74.520 ;
      LAYER met4 ;
        RECT 21.985 74.200 22.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 73.795 22.305 74.115 ;
      LAYER met4 ;
        RECT 21.985 73.795 22.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 73.390 22.305 73.710 ;
      LAYER met4 ;
        RECT 21.985 73.390 22.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 72.985 22.305 73.305 ;
      LAYER met4 ;
        RECT 21.985 72.985 22.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 72.575 22.305 72.895 ;
      LAYER met4 ;
        RECT 21.985 72.575 22.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 72.165 22.305 72.485 ;
      LAYER met4 ;
        RECT 21.985 72.165 22.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 71.755 22.305 72.075 ;
      LAYER met4 ;
        RECT 21.985 71.755 22.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 71.345 22.305 71.665 ;
      LAYER met4 ;
        RECT 21.985 71.345 22.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 70.935 22.305 71.255 ;
      LAYER met4 ;
        RECT 21.985 70.935 22.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 70.525 22.305 70.845 ;
      LAYER met4 ;
        RECT 21.985 70.525 22.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 70.115 22.305 70.435 ;
      LAYER met4 ;
        RECT 21.985 70.115 22.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 69.705 22.305 70.025 ;
      LAYER met4 ;
        RECT 21.985 69.705 22.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 69.295 22.305 69.615 ;
      LAYER met4 ;
        RECT 21.985 69.295 22.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 68.885 22.305 69.205 ;
      LAYER met4 ;
        RECT 21.985 68.885 22.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 68.475 22.305 68.795 ;
      LAYER met4 ;
        RECT 21.985 68.475 22.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.985 68.065 22.305 68.385 ;
      LAYER met4 ;
        RECT 21.985 68.065 22.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 22.160 21.950 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 21.730 21.950 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 21.300 21.950 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 20.870 21.950 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 20.440 21.950 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 20.010 21.950 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 19.580 21.950 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 19.150 21.950 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 18.720 21.950 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 18.290 21.950 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 17.860 21.950 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.655 83.960 21.975 84.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.655 83.410 21.975 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.655 82.860 21.975 83.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 82.300 21.905 82.620 ;
      LAYER met4 ;
        RECT 21.585 82.300 21.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 81.895 21.905 82.215 ;
      LAYER met4 ;
        RECT 21.585 81.895 21.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 81.490 21.905 81.810 ;
      LAYER met4 ;
        RECT 21.585 81.490 21.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 81.085 21.905 81.405 ;
      LAYER met4 ;
        RECT 21.585 81.085 21.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 80.680 21.905 81.000 ;
      LAYER met4 ;
        RECT 21.585 80.680 21.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 80.275 21.905 80.595 ;
      LAYER met4 ;
        RECT 21.585 80.275 21.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 79.870 21.905 80.190 ;
      LAYER met4 ;
        RECT 21.585 79.870 21.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 79.465 21.905 79.785 ;
      LAYER met4 ;
        RECT 21.585 79.465 21.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 79.060 21.905 79.380 ;
      LAYER met4 ;
        RECT 21.585 79.060 21.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 78.655 21.905 78.975 ;
      LAYER met4 ;
        RECT 21.585 78.655 21.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 78.250 21.905 78.570 ;
      LAYER met4 ;
        RECT 21.585 78.250 21.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 77.845 21.905 78.165 ;
      LAYER met4 ;
        RECT 21.585 77.845 21.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 77.440 21.905 77.760 ;
      LAYER met4 ;
        RECT 21.585 77.440 21.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 77.035 21.905 77.355 ;
      LAYER met4 ;
        RECT 21.585 77.035 21.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 76.630 21.905 76.950 ;
      LAYER met4 ;
        RECT 21.585 76.630 21.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 76.225 21.905 76.545 ;
      LAYER met4 ;
        RECT 21.585 76.225 21.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 75.820 21.905 76.140 ;
      LAYER met4 ;
        RECT 21.585 75.820 21.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 75.415 21.905 75.735 ;
      LAYER met4 ;
        RECT 21.585 75.415 21.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 75.010 21.905 75.330 ;
      LAYER met4 ;
        RECT 21.585 75.010 21.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 74.605 21.905 74.925 ;
      LAYER met4 ;
        RECT 21.585 74.605 21.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 74.200 21.905 74.520 ;
      LAYER met4 ;
        RECT 21.585 74.200 21.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 73.795 21.905 74.115 ;
      LAYER met4 ;
        RECT 21.585 73.795 21.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 73.390 21.905 73.710 ;
      LAYER met4 ;
        RECT 21.585 73.390 21.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 72.985 21.905 73.305 ;
      LAYER met4 ;
        RECT 21.585 72.985 21.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 72.575 21.905 72.895 ;
      LAYER met4 ;
        RECT 21.585 72.575 21.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 72.165 21.905 72.485 ;
      LAYER met4 ;
        RECT 21.585 72.165 21.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 71.755 21.905 72.075 ;
      LAYER met4 ;
        RECT 21.585 71.755 21.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 71.345 21.905 71.665 ;
      LAYER met4 ;
        RECT 21.585 71.345 21.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 70.935 21.905 71.255 ;
      LAYER met4 ;
        RECT 21.585 70.935 21.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 70.525 21.905 70.845 ;
      LAYER met4 ;
        RECT 21.585 70.525 21.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 70.115 21.905 70.435 ;
      LAYER met4 ;
        RECT 21.585 70.115 21.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 69.705 21.905 70.025 ;
      LAYER met4 ;
        RECT 21.585 69.705 21.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 69.295 21.905 69.615 ;
      LAYER met4 ;
        RECT 21.585 69.295 21.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 68.885 21.905 69.205 ;
      LAYER met4 ;
        RECT 21.585 68.885 21.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 68.475 21.905 68.795 ;
      LAYER met4 ;
        RECT 21.585 68.475 21.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.585 68.065 21.905 68.385 ;
      LAYER met4 ;
        RECT 21.585 68.065 21.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 22.160 21.545 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 21.730 21.545 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 21.300 21.545 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 20.870 21.545 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 20.440 21.545 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 20.010 21.545 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 19.580 21.545 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 19.150 21.545 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 18.720 21.545 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 18.290 21.545 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.345 17.860 21.545 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 82.300 21.505 82.620 ;
      LAYER met4 ;
        RECT 21.185 82.300 21.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 81.895 21.505 82.215 ;
      LAYER met4 ;
        RECT 21.185 81.895 21.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 81.490 21.505 81.810 ;
      LAYER met4 ;
        RECT 21.185 81.490 21.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 81.085 21.505 81.405 ;
      LAYER met4 ;
        RECT 21.185 81.085 21.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 80.680 21.505 81.000 ;
      LAYER met4 ;
        RECT 21.185 80.680 21.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 80.275 21.505 80.595 ;
      LAYER met4 ;
        RECT 21.185 80.275 21.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 79.870 21.505 80.190 ;
      LAYER met4 ;
        RECT 21.185 79.870 21.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 79.465 21.505 79.785 ;
      LAYER met4 ;
        RECT 21.185 79.465 21.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 79.060 21.505 79.380 ;
      LAYER met4 ;
        RECT 21.185 79.060 21.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 78.655 21.505 78.975 ;
      LAYER met4 ;
        RECT 21.185 78.655 21.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 78.250 21.505 78.570 ;
      LAYER met4 ;
        RECT 21.185 78.250 21.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 77.845 21.505 78.165 ;
      LAYER met4 ;
        RECT 21.185 77.845 21.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 77.440 21.505 77.760 ;
      LAYER met4 ;
        RECT 21.185 77.440 21.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 77.035 21.505 77.355 ;
      LAYER met4 ;
        RECT 21.185 77.035 21.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 76.630 21.505 76.950 ;
      LAYER met4 ;
        RECT 21.185 76.630 21.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 76.225 21.505 76.545 ;
      LAYER met4 ;
        RECT 21.185 76.225 21.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 75.820 21.505 76.140 ;
      LAYER met4 ;
        RECT 21.185 75.820 21.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 75.415 21.505 75.735 ;
      LAYER met4 ;
        RECT 21.185 75.415 21.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 75.010 21.505 75.330 ;
      LAYER met4 ;
        RECT 21.185 75.010 21.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 74.605 21.505 74.925 ;
      LAYER met4 ;
        RECT 21.185 74.605 21.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 74.200 21.505 74.520 ;
      LAYER met4 ;
        RECT 21.185 74.200 21.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 73.795 21.505 74.115 ;
      LAYER met4 ;
        RECT 21.185 73.795 21.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 73.390 21.505 73.710 ;
      LAYER met4 ;
        RECT 21.185 73.390 21.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 72.985 21.505 73.305 ;
      LAYER met4 ;
        RECT 21.185 72.985 21.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 72.575 21.505 72.895 ;
      LAYER met4 ;
        RECT 21.185 72.575 21.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 72.165 21.505 72.485 ;
      LAYER met4 ;
        RECT 21.185 72.165 21.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 71.755 21.505 72.075 ;
      LAYER met4 ;
        RECT 21.185 71.755 21.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 71.345 21.505 71.665 ;
      LAYER met4 ;
        RECT 21.185 71.345 21.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 70.935 21.505 71.255 ;
      LAYER met4 ;
        RECT 21.185 70.935 21.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 70.525 21.505 70.845 ;
      LAYER met4 ;
        RECT 21.185 70.525 21.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 70.115 21.505 70.435 ;
      LAYER met4 ;
        RECT 21.185 70.115 21.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 69.705 21.505 70.025 ;
      LAYER met4 ;
        RECT 21.185 69.705 21.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 69.295 21.505 69.615 ;
      LAYER met4 ;
        RECT 21.185 69.295 21.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 68.885 21.505 69.205 ;
      LAYER met4 ;
        RECT 21.185 68.885 21.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 68.475 21.505 68.795 ;
      LAYER met4 ;
        RECT 21.185 68.475 21.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.185 68.065 21.505 68.385 ;
      LAYER met4 ;
        RECT 21.185 68.065 21.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110 85.265 21.430 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110 84.800 21.430 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110 84.335 21.430 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110 83.870 21.430 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110 83.410 21.430 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.110 82.950 21.430 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 22.160 21.140 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 21.730 21.140 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 21.300 21.140 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 20.870 21.140 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 20.440 21.140 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 20.010 21.140 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 19.580 21.140 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 19.150 21.140 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 18.720 21.140 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 18.290 21.140 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.940 17.860 21.140 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 82.300 21.105 82.620 ;
      LAYER met4 ;
        RECT 20.785 82.300 21.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 81.895 21.105 82.215 ;
      LAYER met4 ;
        RECT 20.785 81.895 21.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 81.490 21.105 81.810 ;
      LAYER met4 ;
        RECT 20.785 81.490 21.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 81.085 21.105 81.405 ;
      LAYER met4 ;
        RECT 20.785 81.085 21.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 80.680 21.105 81.000 ;
      LAYER met4 ;
        RECT 20.785 80.680 21.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 80.275 21.105 80.595 ;
      LAYER met4 ;
        RECT 20.785 80.275 21.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 79.870 21.105 80.190 ;
      LAYER met4 ;
        RECT 20.785 79.870 21.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 79.465 21.105 79.785 ;
      LAYER met4 ;
        RECT 20.785 79.465 21.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 79.060 21.105 79.380 ;
      LAYER met4 ;
        RECT 20.785 79.060 21.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 78.655 21.105 78.975 ;
      LAYER met4 ;
        RECT 20.785 78.655 21.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 78.250 21.105 78.570 ;
      LAYER met4 ;
        RECT 20.785 78.250 21.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 77.845 21.105 78.165 ;
      LAYER met4 ;
        RECT 20.785 77.845 21.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 77.440 21.105 77.760 ;
      LAYER met4 ;
        RECT 20.785 77.440 21.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 77.035 21.105 77.355 ;
      LAYER met4 ;
        RECT 20.785 77.035 21.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 76.630 21.105 76.950 ;
      LAYER met4 ;
        RECT 20.785 76.630 21.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 76.225 21.105 76.545 ;
      LAYER met4 ;
        RECT 20.785 76.225 21.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 75.820 21.105 76.140 ;
      LAYER met4 ;
        RECT 20.785 75.820 21.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 75.415 21.105 75.735 ;
      LAYER met4 ;
        RECT 20.785 75.415 21.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 75.010 21.105 75.330 ;
      LAYER met4 ;
        RECT 20.785 75.010 21.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 74.605 21.105 74.925 ;
      LAYER met4 ;
        RECT 20.785 74.605 21.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 74.200 21.105 74.520 ;
      LAYER met4 ;
        RECT 20.785 74.200 21.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 73.795 21.105 74.115 ;
      LAYER met4 ;
        RECT 20.785 73.795 21.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 73.390 21.105 73.710 ;
      LAYER met4 ;
        RECT 20.785 73.390 21.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 72.985 21.105 73.305 ;
      LAYER met4 ;
        RECT 20.785 72.985 21.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 72.575 21.105 72.895 ;
      LAYER met4 ;
        RECT 20.785 72.575 21.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 72.165 21.105 72.485 ;
      LAYER met4 ;
        RECT 20.785 72.165 21.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 71.755 21.105 72.075 ;
      LAYER met4 ;
        RECT 20.785 71.755 21.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 71.345 21.105 71.665 ;
      LAYER met4 ;
        RECT 20.785 71.345 21.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 70.935 21.105 71.255 ;
      LAYER met4 ;
        RECT 20.785 70.935 21.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 70.525 21.105 70.845 ;
      LAYER met4 ;
        RECT 20.785 70.525 21.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 70.115 21.105 70.435 ;
      LAYER met4 ;
        RECT 20.785 70.115 21.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 69.705 21.105 70.025 ;
      LAYER met4 ;
        RECT 20.785 69.705 21.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 69.295 21.105 69.615 ;
      LAYER met4 ;
        RECT 20.785 69.295 21.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 68.885 21.105 69.205 ;
      LAYER met4 ;
        RECT 20.785 68.885 21.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 68.475 21.105 68.795 ;
      LAYER met4 ;
        RECT 20.785 68.475 21.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.785 68.065 21.105 68.385 ;
      LAYER met4 ;
        RECT 20.785 68.065 21.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630 85.265 20.950 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630 84.800 20.950 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630 84.335 20.950 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630 83.870 20.950 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630 83.410 20.950 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.630 82.950 20.950 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 22.160 20.735 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 21.730 20.735 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 21.300 20.735 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 20.870 20.735 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 20.440 20.735 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 20.010 20.735 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 19.580 20.735 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 19.150 20.735 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 18.720 20.735 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 18.290 20.735 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.535 17.860 20.735 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 82.300 20.705 82.620 ;
      LAYER met4 ;
        RECT 20.385 82.300 20.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 81.895 20.705 82.215 ;
      LAYER met4 ;
        RECT 20.385 81.895 20.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 81.490 20.705 81.810 ;
      LAYER met4 ;
        RECT 20.385 81.490 20.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 81.085 20.705 81.405 ;
      LAYER met4 ;
        RECT 20.385 81.085 20.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 80.680 20.705 81.000 ;
      LAYER met4 ;
        RECT 20.385 80.680 20.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 80.275 20.705 80.595 ;
      LAYER met4 ;
        RECT 20.385 80.275 20.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 79.870 20.705 80.190 ;
      LAYER met4 ;
        RECT 20.385 79.870 20.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 79.465 20.705 79.785 ;
      LAYER met4 ;
        RECT 20.385 79.465 20.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 79.060 20.705 79.380 ;
      LAYER met4 ;
        RECT 20.385 79.060 20.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 78.655 20.705 78.975 ;
      LAYER met4 ;
        RECT 20.385 78.655 20.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 78.250 20.705 78.570 ;
      LAYER met4 ;
        RECT 20.385 78.250 20.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 77.845 20.705 78.165 ;
      LAYER met4 ;
        RECT 20.385 77.845 20.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 77.440 20.705 77.760 ;
      LAYER met4 ;
        RECT 20.385 77.440 20.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 77.035 20.705 77.355 ;
      LAYER met4 ;
        RECT 20.385 77.035 20.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 76.630 20.705 76.950 ;
      LAYER met4 ;
        RECT 20.385 76.630 20.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 76.225 20.705 76.545 ;
      LAYER met4 ;
        RECT 20.385 76.225 20.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 75.820 20.705 76.140 ;
      LAYER met4 ;
        RECT 20.385 75.820 20.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 75.415 20.705 75.735 ;
      LAYER met4 ;
        RECT 20.385 75.415 20.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 75.010 20.705 75.330 ;
      LAYER met4 ;
        RECT 20.385 75.010 20.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 74.605 20.705 74.925 ;
      LAYER met4 ;
        RECT 20.385 74.605 20.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 74.200 20.705 74.520 ;
      LAYER met4 ;
        RECT 20.385 74.200 20.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 73.795 20.705 74.115 ;
      LAYER met4 ;
        RECT 20.385 73.795 20.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 73.390 20.705 73.710 ;
      LAYER met4 ;
        RECT 20.385 73.390 20.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 72.985 20.705 73.305 ;
      LAYER met4 ;
        RECT 20.385 72.985 20.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 72.575 20.705 72.895 ;
      LAYER met4 ;
        RECT 20.385 72.575 20.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 72.165 20.705 72.485 ;
      LAYER met4 ;
        RECT 20.385 72.165 20.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 71.755 20.705 72.075 ;
      LAYER met4 ;
        RECT 20.385 71.755 20.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 71.345 20.705 71.665 ;
      LAYER met4 ;
        RECT 20.385 71.345 20.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 70.935 20.705 71.255 ;
      LAYER met4 ;
        RECT 20.385 70.935 20.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 70.525 20.705 70.845 ;
      LAYER met4 ;
        RECT 20.385 70.525 20.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 70.115 20.705 70.435 ;
      LAYER met4 ;
        RECT 20.385 70.115 20.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 69.705 20.705 70.025 ;
      LAYER met4 ;
        RECT 20.385 69.705 20.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 69.295 20.705 69.615 ;
      LAYER met4 ;
        RECT 20.385 69.295 20.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 68.885 20.705 69.205 ;
      LAYER met4 ;
        RECT 20.385 68.885 20.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 68.475 20.705 68.795 ;
      LAYER met4 ;
        RECT 20.385 68.475 20.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.385 68.065 20.705 68.385 ;
      LAYER met4 ;
        RECT 20.385 68.065 20.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 85.265 20.470 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 84.800 20.470 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 84.335 20.470 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 83.870 20.470 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 83.410 20.470 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 82.950 20.470 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 22.160 20.330 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 21.730 20.330 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 21.300 20.330 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 20.870 20.330 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 20.440 20.330 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 20.010 20.330 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 19.580 20.330 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 19.150 20.330 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 18.720 20.330 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 18.290 20.330 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.130 17.860 20.330 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 82.300 20.305 82.620 ;
      LAYER met4 ;
        RECT 19.985 82.300 20.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 81.895 20.305 82.215 ;
      LAYER met4 ;
        RECT 19.985 81.895 20.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 81.490 20.305 81.810 ;
      LAYER met4 ;
        RECT 19.985 81.490 20.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 81.085 20.305 81.405 ;
      LAYER met4 ;
        RECT 19.985 81.085 20.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 80.680 20.305 81.000 ;
      LAYER met4 ;
        RECT 19.985 80.680 20.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 80.275 20.305 80.595 ;
      LAYER met4 ;
        RECT 19.985 80.275 20.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 79.870 20.305 80.190 ;
      LAYER met4 ;
        RECT 19.985 79.870 20.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 79.465 20.305 79.785 ;
      LAYER met4 ;
        RECT 19.985 79.465 20.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 79.060 20.305 79.380 ;
      LAYER met4 ;
        RECT 19.985 79.060 20.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 78.655 20.305 78.975 ;
      LAYER met4 ;
        RECT 19.985 78.655 20.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 78.250 20.305 78.570 ;
      LAYER met4 ;
        RECT 19.985 78.250 20.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 77.845 20.305 78.165 ;
      LAYER met4 ;
        RECT 19.985 77.845 20.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 77.440 20.305 77.760 ;
      LAYER met4 ;
        RECT 19.985 77.440 20.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 77.035 20.305 77.355 ;
      LAYER met4 ;
        RECT 19.985 77.035 20.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 76.630 20.305 76.950 ;
      LAYER met4 ;
        RECT 19.985 76.630 20.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 76.225 20.305 76.545 ;
      LAYER met4 ;
        RECT 19.985 76.225 20.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 75.820 20.305 76.140 ;
      LAYER met4 ;
        RECT 19.985 75.820 20.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 75.415 20.305 75.735 ;
      LAYER met4 ;
        RECT 19.985 75.415 20.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 75.010 20.305 75.330 ;
      LAYER met4 ;
        RECT 19.985 75.010 20.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 74.605 20.305 74.925 ;
      LAYER met4 ;
        RECT 19.985 74.605 20.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 74.200 20.305 74.520 ;
      LAYER met4 ;
        RECT 19.985 74.200 20.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 73.795 20.305 74.115 ;
      LAYER met4 ;
        RECT 19.985 73.795 20.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 73.390 20.305 73.710 ;
      LAYER met4 ;
        RECT 19.985 73.390 20.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 72.985 20.305 73.305 ;
      LAYER met4 ;
        RECT 19.985 72.985 20.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 72.575 20.305 72.895 ;
      LAYER met4 ;
        RECT 19.985 72.575 20.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 72.165 20.305 72.485 ;
      LAYER met4 ;
        RECT 19.985 72.165 20.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 71.755 20.305 72.075 ;
      LAYER met4 ;
        RECT 19.985 71.755 20.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 71.345 20.305 71.665 ;
      LAYER met4 ;
        RECT 19.985 71.345 20.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 70.935 20.305 71.255 ;
      LAYER met4 ;
        RECT 19.985 70.935 20.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 70.525 20.305 70.845 ;
      LAYER met4 ;
        RECT 19.985 70.525 20.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 70.115 20.305 70.435 ;
      LAYER met4 ;
        RECT 19.985 70.115 20.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 69.705 20.305 70.025 ;
      LAYER met4 ;
        RECT 19.985 69.705 20.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 69.295 20.305 69.615 ;
      LAYER met4 ;
        RECT 19.985 69.295 20.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 68.885 20.305 69.205 ;
      LAYER met4 ;
        RECT 19.985 68.885 20.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 68.475 20.305 68.795 ;
      LAYER met4 ;
        RECT 19.985 68.475 20.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.985 68.065 20.305 68.385 ;
      LAYER met4 ;
        RECT 19.985 68.065 20.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.740 86.690 20.060 87.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.740 86.250 20.060 86.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.740 85.815 20.060 86.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670 85.265 19.990 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670 84.800 19.990 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670 84.335 19.990 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670 83.870 19.990 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670 83.410 19.990 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.670 82.950 19.990 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 22.160 19.925 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 21.730 19.925 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 21.300 19.925 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 20.870 19.925 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 20.440 19.925 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 20.010 19.925 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 19.580 19.925 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 19.150 19.925 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 18.720 19.925 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 18.290 19.925 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.725 17.860 19.925 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 82.300 19.905 82.620 ;
      LAYER met4 ;
        RECT 19.585 82.300 19.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 81.895 19.905 82.215 ;
      LAYER met4 ;
        RECT 19.585 81.895 19.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 81.490 19.905 81.810 ;
      LAYER met4 ;
        RECT 19.585 81.490 19.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 81.085 19.905 81.405 ;
      LAYER met4 ;
        RECT 19.585 81.085 19.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 80.680 19.905 81.000 ;
      LAYER met4 ;
        RECT 19.585 80.680 19.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 80.275 19.905 80.595 ;
      LAYER met4 ;
        RECT 19.585 80.275 19.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 79.870 19.905 80.190 ;
      LAYER met4 ;
        RECT 19.585 79.870 19.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 79.465 19.905 79.785 ;
      LAYER met4 ;
        RECT 19.585 79.465 19.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 79.060 19.905 79.380 ;
      LAYER met4 ;
        RECT 19.585 79.060 19.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 78.655 19.905 78.975 ;
      LAYER met4 ;
        RECT 19.585 78.655 19.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 78.250 19.905 78.570 ;
      LAYER met4 ;
        RECT 19.585 78.250 19.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 77.845 19.905 78.165 ;
      LAYER met4 ;
        RECT 19.585 77.845 19.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 77.440 19.905 77.760 ;
      LAYER met4 ;
        RECT 19.585 77.440 19.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 77.035 19.905 77.355 ;
      LAYER met4 ;
        RECT 19.585 77.035 19.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 76.630 19.905 76.950 ;
      LAYER met4 ;
        RECT 19.585 76.630 19.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 76.225 19.905 76.545 ;
      LAYER met4 ;
        RECT 19.585 76.225 19.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 75.820 19.905 76.140 ;
      LAYER met4 ;
        RECT 19.585 75.820 19.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 75.415 19.905 75.735 ;
      LAYER met4 ;
        RECT 19.585 75.415 19.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 75.010 19.905 75.330 ;
      LAYER met4 ;
        RECT 19.585 75.010 19.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 74.605 19.905 74.925 ;
      LAYER met4 ;
        RECT 19.585 74.605 19.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 74.200 19.905 74.520 ;
      LAYER met4 ;
        RECT 19.585 74.200 19.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 73.795 19.905 74.115 ;
      LAYER met4 ;
        RECT 19.585 73.795 19.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 73.390 19.905 73.710 ;
      LAYER met4 ;
        RECT 19.585 73.390 19.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 72.985 19.905 73.305 ;
      LAYER met4 ;
        RECT 19.585 72.985 19.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 72.575 19.905 72.895 ;
      LAYER met4 ;
        RECT 19.585 72.575 19.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 72.165 19.905 72.485 ;
      LAYER met4 ;
        RECT 19.585 72.165 19.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 71.755 19.905 72.075 ;
      LAYER met4 ;
        RECT 19.585 71.755 19.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 71.345 19.905 71.665 ;
      LAYER met4 ;
        RECT 19.585 71.345 19.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 70.935 19.905 71.255 ;
      LAYER met4 ;
        RECT 19.585 70.935 19.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 70.525 19.905 70.845 ;
      LAYER met4 ;
        RECT 19.585 70.525 19.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 70.115 19.905 70.435 ;
      LAYER met4 ;
        RECT 19.585 70.115 19.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 69.705 19.905 70.025 ;
      LAYER met4 ;
        RECT 19.585 69.705 19.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 69.295 19.905 69.615 ;
      LAYER met4 ;
        RECT 19.585 69.295 19.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 68.885 19.905 69.205 ;
      LAYER met4 ;
        RECT 19.585 68.885 19.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 68.475 19.905 68.795 ;
      LAYER met4 ;
        RECT 19.585 68.475 19.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.585 68.065 19.905 68.385 ;
      LAYER met4 ;
        RECT 19.585 68.065 19.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 22.160 19.520 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 21.730 19.520 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 21.300 19.520 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 20.870 19.520 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 20.440 19.520 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 20.010 19.520 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 19.580 19.520 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 19.150 19.520 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 18.720 19.520 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 18.290 19.520 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.320 17.860 19.520 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 85.265 19.510 85.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 84.800 19.510 85.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 84.335 19.510 84.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 83.870 19.510 84.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 83.410 19.510 83.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 82.950 19.510 83.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 82.300 19.505 82.620 ;
      LAYER met4 ;
        RECT 19.185 82.300 19.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 81.895 19.505 82.215 ;
      LAYER met4 ;
        RECT 19.185 81.895 19.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 81.490 19.505 81.810 ;
      LAYER met4 ;
        RECT 19.185 81.490 19.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 81.085 19.505 81.405 ;
      LAYER met4 ;
        RECT 19.185 81.085 19.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 80.680 19.505 81.000 ;
      LAYER met4 ;
        RECT 19.185 80.680 19.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 80.275 19.505 80.595 ;
      LAYER met4 ;
        RECT 19.185 80.275 19.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 79.870 19.505 80.190 ;
      LAYER met4 ;
        RECT 19.185 79.870 19.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 79.465 19.505 79.785 ;
      LAYER met4 ;
        RECT 19.185 79.465 19.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 79.060 19.505 79.380 ;
      LAYER met4 ;
        RECT 19.185 79.060 19.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 78.655 19.505 78.975 ;
      LAYER met4 ;
        RECT 19.185 78.655 19.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 78.250 19.505 78.570 ;
      LAYER met4 ;
        RECT 19.185 78.250 19.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 77.845 19.505 78.165 ;
      LAYER met4 ;
        RECT 19.185 77.845 19.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 77.440 19.505 77.760 ;
      LAYER met4 ;
        RECT 19.185 77.440 19.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 77.035 19.505 77.355 ;
      LAYER met4 ;
        RECT 19.185 77.035 19.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 76.630 19.505 76.950 ;
      LAYER met4 ;
        RECT 19.185 76.630 19.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 76.225 19.505 76.545 ;
      LAYER met4 ;
        RECT 19.185 76.225 19.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 75.820 19.505 76.140 ;
      LAYER met4 ;
        RECT 19.185 75.820 19.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 75.415 19.505 75.735 ;
      LAYER met4 ;
        RECT 19.185 75.415 19.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 75.010 19.505 75.330 ;
      LAYER met4 ;
        RECT 19.185 75.010 19.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 74.605 19.505 74.925 ;
      LAYER met4 ;
        RECT 19.185 74.605 19.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 74.200 19.505 74.520 ;
      LAYER met4 ;
        RECT 19.185 74.200 19.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 73.795 19.505 74.115 ;
      LAYER met4 ;
        RECT 19.185 73.795 19.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 73.390 19.505 73.710 ;
      LAYER met4 ;
        RECT 19.185 73.390 19.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 72.985 19.505 73.305 ;
      LAYER met4 ;
        RECT 19.185 72.985 19.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 72.575 19.505 72.895 ;
      LAYER met4 ;
        RECT 19.185 72.575 19.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 72.165 19.505 72.485 ;
      LAYER met4 ;
        RECT 19.185 72.165 19.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 71.755 19.505 72.075 ;
      LAYER met4 ;
        RECT 19.185 71.755 19.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 71.345 19.505 71.665 ;
      LAYER met4 ;
        RECT 19.185 71.345 19.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 70.935 19.505 71.255 ;
      LAYER met4 ;
        RECT 19.185 70.935 19.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 70.525 19.505 70.845 ;
      LAYER met4 ;
        RECT 19.185 70.525 19.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 70.115 19.505 70.435 ;
      LAYER met4 ;
        RECT 19.185 70.115 19.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 69.705 19.505 70.025 ;
      LAYER met4 ;
        RECT 19.185 69.705 19.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 69.295 19.505 69.615 ;
      LAYER met4 ;
        RECT 19.185 69.295 19.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 68.885 19.505 69.205 ;
      LAYER met4 ;
        RECT 19.185 68.885 19.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 68.475 19.505 68.795 ;
      LAYER met4 ;
        RECT 19.185 68.475 19.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 68.065 19.505 68.385 ;
      LAYER met4 ;
        RECT 19.185 68.065 19.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.000 86.690 19.320 87.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.000 86.250 19.320 86.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.000 85.815 19.320 86.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 22.160 19.115 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 21.730 19.115 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 21.300 19.115 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 20.870 19.115 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 20.440 19.115 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 20.010 19.115 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 19.580 19.115 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 19.150 19.115 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 18.720 19.115 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 18.290 19.115 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.915 17.860 19.115 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 82.300 19.105 82.620 ;
      LAYER met4 ;
        RECT 18.785 82.300 19.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 81.895 19.105 82.215 ;
      LAYER met4 ;
        RECT 18.785 81.895 19.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 81.490 19.105 81.810 ;
      LAYER met4 ;
        RECT 18.785 81.490 19.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 81.085 19.105 81.405 ;
      LAYER met4 ;
        RECT 18.785 81.085 19.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 80.680 19.105 81.000 ;
      LAYER met4 ;
        RECT 18.785 80.680 19.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 80.275 19.105 80.595 ;
      LAYER met4 ;
        RECT 18.785 80.275 19.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 79.870 19.105 80.190 ;
      LAYER met4 ;
        RECT 18.785 79.870 19.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 79.465 19.105 79.785 ;
      LAYER met4 ;
        RECT 18.785 79.465 19.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 79.060 19.105 79.380 ;
      LAYER met4 ;
        RECT 18.785 79.060 19.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 78.655 19.105 78.975 ;
      LAYER met4 ;
        RECT 18.785 78.655 19.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 78.250 19.105 78.570 ;
      LAYER met4 ;
        RECT 18.785 78.250 19.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 77.845 19.105 78.165 ;
      LAYER met4 ;
        RECT 18.785 77.845 19.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 77.440 19.105 77.760 ;
      LAYER met4 ;
        RECT 18.785 77.440 19.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 77.035 19.105 77.355 ;
      LAYER met4 ;
        RECT 18.785 77.035 19.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 76.630 19.105 76.950 ;
      LAYER met4 ;
        RECT 18.785 76.630 19.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 76.225 19.105 76.545 ;
      LAYER met4 ;
        RECT 18.785 76.225 19.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 75.820 19.105 76.140 ;
      LAYER met4 ;
        RECT 18.785 75.820 19.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 75.415 19.105 75.735 ;
      LAYER met4 ;
        RECT 18.785 75.415 19.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 75.010 19.105 75.330 ;
      LAYER met4 ;
        RECT 18.785 75.010 19.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 74.605 19.105 74.925 ;
      LAYER met4 ;
        RECT 18.785 74.605 19.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 74.200 19.105 74.520 ;
      LAYER met4 ;
        RECT 18.785 74.200 19.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 73.795 19.105 74.115 ;
      LAYER met4 ;
        RECT 18.785 73.795 19.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 73.390 19.105 73.710 ;
      LAYER met4 ;
        RECT 18.785 73.390 19.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 72.985 19.105 73.305 ;
      LAYER met4 ;
        RECT 18.785 72.985 19.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 72.575 19.105 72.895 ;
      LAYER met4 ;
        RECT 18.785 72.575 19.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 72.165 19.105 72.485 ;
      LAYER met4 ;
        RECT 18.785 72.165 19.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 71.755 19.105 72.075 ;
      LAYER met4 ;
        RECT 18.785 71.755 19.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 71.345 19.105 71.665 ;
      LAYER met4 ;
        RECT 18.785 71.345 19.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 70.935 19.105 71.255 ;
      LAYER met4 ;
        RECT 18.785 70.935 19.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 70.525 19.105 70.845 ;
      LAYER met4 ;
        RECT 18.785 70.525 19.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 70.115 19.105 70.435 ;
      LAYER met4 ;
        RECT 18.785 70.115 19.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 69.705 19.105 70.025 ;
      LAYER met4 ;
        RECT 18.785 69.705 19.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 69.295 19.105 69.615 ;
      LAYER met4 ;
        RECT 18.785 69.295 19.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 68.885 19.105 69.205 ;
      LAYER met4 ;
        RECT 18.785 68.885 19.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 68.475 19.105 68.795 ;
      LAYER met4 ;
        RECT 18.785 68.475 19.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 68.065 19.105 68.385 ;
      LAYER met4 ;
        RECT 18.785 68.065 19.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 87.815 18.825 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 87.410 18.825 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 87.005 18.825 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 86.600 18.825 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 86.195 18.825 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 85.795 18.825 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 85.395 18.825 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 84.995 18.825 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 84.595 18.825 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 84.195 18.825 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 83.795 18.825 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 83.395 18.825 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.505 82.995 18.825 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 22.160 18.710 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 21.730 18.710 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 21.300 18.710 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 20.870 18.710 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 20.440 18.710 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 20.010 18.710 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 19.580 18.710 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 19.150 18.710 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 18.720 18.710 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 18.290 18.710 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.510 17.860 18.710 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 82.300 18.705 82.620 ;
      LAYER met4 ;
        RECT 18.385 82.300 18.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 81.895 18.705 82.215 ;
      LAYER met4 ;
        RECT 18.385 81.895 18.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 81.490 18.705 81.810 ;
      LAYER met4 ;
        RECT 18.385 81.490 18.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 81.085 18.705 81.405 ;
      LAYER met4 ;
        RECT 18.385 81.085 18.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 80.680 18.705 81.000 ;
      LAYER met4 ;
        RECT 18.385 80.680 18.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 80.275 18.705 80.595 ;
      LAYER met4 ;
        RECT 18.385 80.275 18.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 79.870 18.705 80.190 ;
      LAYER met4 ;
        RECT 18.385 79.870 18.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 79.465 18.705 79.785 ;
      LAYER met4 ;
        RECT 18.385 79.465 18.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 79.060 18.705 79.380 ;
      LAYER met4 ;
        RECT 18.385 79.060 18.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 78.655 18.705 78.975 ;
      LAYER met4 ;
        RECT 18.385 78.655 18.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 78.250 18.705 78.570 ;
      LAYER met4 ;
        RECT 18.385 78.250 18.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 77.845 18.705 78.165 ;
      LAYER met4 ;
        RECT 18.385 77.845 18.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 77.440 18.705 77.760 ;
      LAYER met4 ;
        RECT 18.385 77.440 18.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 77.035 18.705 77.355 ;
      LAYER met4 ;
        RECT 18.385 77.035 18.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 76.630 18.705 76.950 ;
      LAYER met4 ;
        RECT 18.385 76.630 18.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 76.225 18.705 76.545 ;
      LAYER met4 ;
        RECT 18.385 76.225 18.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 75.820 18.705 76.140 ;
      LAYER met4 ;
        RECT 18.385 75.820 18.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 75.415 18.705 75.735 ;
      LAYER met4 ;
        RECT 18.385 75.415 18.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 75.010 18.705 75.330 ;
      LAYER met4 ;
        RECT 18.385 75.010 18.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 74.605 18.705 74.925 ;
      LAYER met4 ;
        RECT 18.385 74.605 18.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 74.200 18.705 74.520 ;
      LAYER met4 ;
        RECT 18.385 74.200 18.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 73.795 18.705 74.115 ;
      LAYER met4 ;
        RECT 18.385 73.795 18.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 73.390 18.705 73.710 ;
      LAYER met4 ;
        RECT 18.385 73.390 18.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 72.985 18.705 73.305 ;
      LAYER met4 ;
        RECT 18.385 72.985 18.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 72.575 18.705 72.895 ;
      LAYER met4 ;
        RECT 18.385 72.575 18.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 72.165 18.705 72.485 ;
      LAYER met4 ;
        RECT 18.385 72.165 18.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 71.755 18.705 72.075 ;
      LAYER met4 ;
        RECT 18.385 71.755 18.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 71.345 18.705 71.665 ;
      LAYER met4 ;
        RECT 18.385 71.345 18.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 70.935 18.705 71.255 ;
      LAYER met4 ;
        RECT 18.385 70.935 18.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 70.525 18.705 70.845 ;
      LAYER met4 ;
        RECT 18.385 70.525 18.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 70.115 18.705 70.435 ;
      LAYER met4 ;
        RECT 18.385 70.115 18.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 69.705 18.705 70.025 ;
      LAYER met4 ;
        RECT 18.385 69.705 18.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 69.295 18.705 69.615 ;
      LAYER met4 ;
        RECT 18.385 69.295 18.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 68.885 18.705 69.205 ;
      LAYER met4 ;
        RECT 18.385 68.885 18.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 68.475 18.705 68.795 ;
      LAYER met4 ;
        RECT 18.385 68.475 18.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.385 68.065 18.705 68.385 ;
      LAYER met4 ;
        RECT 18.385 68.065 18.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 87.815 18.415 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 87.410 18.415 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 87.005 18.415 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 86.600 18.415 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 86.195 18.415 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 85.795 18.415 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 85.395 18.415 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 84.995 18.415 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 84.595 18.415 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 84.195 18.415 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 83.795 18.415 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 83.395 18.415 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.095 82.995 18.415 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 22.160 18.305 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 21.730 18.305 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 21.300 18.305 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 20.870 18.305 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 20.440 18.305 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 20.010 18.305 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 19.580 18.305 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 19.150 18.305 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 18.720 18.305 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 18.290 18.305 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.105 17.860 18.305 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 82.300 18.305 82.620 ;
      LAYER met4 ;
        RECT 17.985 82.300 18.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 81.895 18.305 82.215 ;
      LAYER met4 ;
        RECT 17.985 81.895 18.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 81.490 18.305 81.810 ;
      LAYER met4 ;
        RECT 17.985 81.490 18.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 81.085 18.305 81.405 ;
      LAYER met4 ;
        RECT 17.985 81.085 18.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 80.680 18.305 81.000 ;
      LAYER met4 ;
        RECT 17.985 80.680 18.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 80.275 18.305 80.595 ;
      LAYER met4 ;
        RECT 17.985 80.275 18.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 79.870 18.305 80.190 ;
      LAYER met4 ;
        RECT 17.985 79.870 18.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 79.465 18.305 79.785 ;
      LAYER met4 ;
        RECT 17.985 79.465 18.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 79.060 18.305 79.380 ;
      LAYER met4 ;
        RECT 17.985 79.060 18.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 78.655 18.305 78.975 ;
      LAYER met4 ;
        RECT 17.985 78.655 18.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 78.250 18.305 78.570 ;
      LAYER met4 ;
        RECT 17.985 78.250 18.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 77.845 18.305 78.165 ;
      LAYER met4 ;
        RECT 17.985 77.845 18.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 77.440 18.305 77.760 ;
      LAYER met4 ;
        RECT 17.985 77.440 18.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 77.035 18.305 77.355 ;
      LAYER met4 ;
        RECT 17.985 77.035 18.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 76.630 18.305 76.950 ;
      LAYER met4 ;
        RECT 17.985 76.630 18.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 76.225 18.305 76.545 ;
      LAYER met4 ;
        RECT 17.985 76.225 18.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 75.820 18.305 76.140 ;
      LAYER met4 ;
        RECT 17.985 75.820 18.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 75.415 18.305 75.735 ;
      LAYER met4 ;
        RECT 17.985 75.415 18.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 75.010 18.305 75.330 ;
      LAYER met4 ;
        RECT 17.985 75.010 18.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 74.605 18.305 74.925 ;
      LAYER met4 ;
        RECT 17.985 74.605 18.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 74.200 18.305 74.520 ;
      LAYER met4 ;
        RECT 17.985 74.200 18.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 73.795 18.305 74.115 ;
      LAYER met4 ;
        RECT 17.985 73.795 18.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 73.390 18.305 73.710 ;
      LAYER met4 ;
        RECT 17.985 73.390 18.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 72.985 18.305 73.305 ;
      LAYER met4 ;
        RECT 17.985 72.985 18.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 72.575 18.305 72.895 ;
      LAYER met4 ;
        RECT 17.985 72.575 18.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 72.165 18.305 72.485 ;
      LAYER met4 ;
        RECT 17.985 72.165 18.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 71.755 18.305 72.075 ;
      LAYER met4 ;
        RECT 17.985 71.755 18.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 71.345 18.305 71.665 ;
      LAYER met4 ;
        RECT 17.985 71.345 18.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 70.935 18.305 71.255 ;
      LAYER met4 ;
        RECT 17.985 70.935 18.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 70.525 18.305 70.845 ;
      LAYER met4 ;
        RECT 17.985 70.525 18.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 70.115 18.305 70.435 ;
      LAYER met4 ;
        RECT 17.985 70.115 18.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 69.705 18.305 70.025 ;
      LAYER met4 ;
        RECT 17.985 69.705 18.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 69.295 18.305 69.615 ;
      LAYER met4 ;
        RECT 17.985 69.295 18.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 68.885 18.305 69.205 ;
      LAYER met4 ;
        RECT 17.985 68.885 18.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 68.475 18.305 68.795 ;
      LAYER met4 ;
        RECT 17.985 68.475 18.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.985 68.065 18.305 68.385 ;
      LAYER met4 ;
        RECT 17.985 68.065 18.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 87.815 18.005 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 87.410 18.005 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 87.005 18.005 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 86.600 18.005 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 86.195 18.005 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 85.795 18.005 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 85.395 18.005 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 84.995 18.005 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 84.595 18.005 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 84.195 18.005 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 83.795 18.005 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 83.395 18.005 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 82.995 18.005 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 22.160 17.900 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 21.730 17.900 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 21.300 17.900 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 20.870 17.900 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 20.440 17.900 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 20.010 17.900 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 19.580 17.900 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 19.150 17.900 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 18.720 17.900 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 18.290 17.900 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.700 17.860 17.900 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 82.300 17.905 82.620 ;
      LAYER met4 ;
        RECT 17.585 82.300 17.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 81.895 17.905 82.215 ;
      LAYER met4 ;
        RECT 17.585 81.895 17.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 81.490 17.905 81.810 ;
      LAYER met4 ;
        RECT 17.585 81.490 17.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 81.085 17.905 81.405 ;
      LAYER met4 ;
        RECT 17.585 81.085 17.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 80.680 17.905 81.000 ;
      LAYER met4 ;
        RECT 17.585 80.680 17.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 80.275 17.905 80.595 ;
      LAYER met4 ;
        RECT 17.585 80.275 17.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 79.870 17.905 80.190 ;
      LAYER met4 ;
        RECT 17.585 79.870 17.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 79.465 17.905 79.785 ;
      LAYER met4 ;
        RECT 17.585 79.465 17.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 79.060 17.905 79.380 ;
      LAYER met4 ;
        RECT 17.585 79.060 17.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 78.655 17.905 78.975 ;
      LAYER met4 ;
        RECT 17.585 78.655 17.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 78.250 17.905 78.570 ;
      LAYER met4 ;
        RECT 17.585 78.250 17.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 77.845 17.905 78.165 ;
      LAYER met4 ;
        RECT 17.585 77.845 17.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 77.440 17.905 77.760 ;
      LAYER met4 ;
        RECT 17.585 77.440 17.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 77.035 17.905 77.355 ;
      LAYER met4 ;
        RECT 17.585 77.035 17.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 76.630 17.905 76.950 ;
      LAYER met4 ;
        RECT 17.585 76.630 17.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 76.225 17.905 76.545 ;
      LAYER met4 ;
        RECT 17.585 76.225 17.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 75.820 17.905 76.140 ;
      LAYER met4 ;
        RECT 17.585 75.820 17.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 75.415 17.905 75.735 ;
      LAYER met4 ;
        RECT 17.585 75.415 17.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 75.010 17.905 75.330 ;
      LAYER met4 ;
        RECT 17.585 75.010 17.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 74.605 17.905 74.925 ;
      LAYER met4 ;
        RECT 17.585 74.605 17.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 74.200 17.905 74.520 ;
      LAYER met4 ;
        RECT 17.585 74.200 17.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 73.795 17.905 74.115 ;
      LAYER met4 ;
        RECT 17.585 73.795 17.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 73.390 17.905 73.710 ;
      LAYER met4 ;
        RECT 17.585 73.390 17.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 72.985 17.905 73.305 ;
      LAYER met4 ;
        RECT 17.585 72.985 17.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 72.575 17.905 72.895 ;
      LAYER met4 ;
        RECT 17.585 72.575 17.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 72.165 17.905 72.485 ;
      LAYER met4 ;
        RECT 17.585 72.165 17.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 71.755 17.905 72.075 ;
      LAYER met4 ;
        RECT 17.585 71.755 17.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 71.345 17.905 71.665 ;
      LAYER met4 ;
        RECT 17.585 71.345 17.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 70.935 17.905 71.255 ;
      LAYER met4 ;
        RECT 17.585 70.935 17.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 70.525 17.905 70.845 ;
      LAYER met4 ;
        RECT 17.585 70.525 17.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 70.115 17.905 70.435 ;
      LAYER met4 ;
        RECT 17.585 70.115 17.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 69.705 17.905 70.025 ;
      LAYER met4 ;
        RECT 17.585 69.705 17.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 69.295 17.905 69.615 ;
      LAYER met4 ;
        RECT 17.585 69.295 17.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 68.885 17.905 69.205 ;
      LAYER met4 ;
        RECT 17.585 68.885 17.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 68.475 17.905 68.795 ;
      LAYER met4 ;
        RECT 17.585 68.475 17.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.585 68.065 17.905 68.385 ;
      LAYER met4 ;
        RECT 17.585 68.065 17.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 87.815 17.595 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 87.410 17.595 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 87.005 17.595 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 86.600 17.595 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 86.195 17.595 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 85.795 17.595 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 85.395 17.595 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 84.995 17.595 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 84.595 17.595 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 84.195 17.595 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 83.795 17.595 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 83.395 17.595 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.275 82.995 17.595 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 22.160 17.495 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 21.730 17.495 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 21.300 17.495 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 20.870 17.495 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 20.440 17.495 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 20.010 17.495 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 19.580 17.495 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 19.150 17.495 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 18.720 17.495 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 18.290 17.495 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 17.860 17.495 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 89.205 17.520 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 88.785 17.520 89.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 88.370 17.520 88.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 82.300 17.505 82.620 ;
      LAYER met4 ;
        RECT 17.185 82.300 17.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 81.895 17.505 82.215 ;
      LAYER met4 ;
        RECT 17.185 81.895 17.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 81.490 17.505 81.810 ;
      LAYER met4 ;
        RECT 17.185 81.490 17.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 81.085 17.505 81.405 ;
      LAYER met4 ;
        RECT 17.185 81.085 17.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 80.680 17.505 81.000 ;
      LAYER met4 ;
        RECT 17.185 80.680 17.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 80.275 17.505 80.595 ;
      LAYER met4 ;
        RECT 17.185 80.275 17.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 79.870 17.505 80.190 ;
      LAYER met4 ;
        RECT 17.185 79.870 17.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 79.465 17.505 79.785 ;
      LAYER met4 ;
        RECT 17.185 79.465 17.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 79.060 17.505 79.380 ;
      LAYER met4 ;
        RECT 17.185 79.060 17.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 78.655 17.505 78.975 ;
      LAYER met4 ;
        RECT 17.185 78.655 17.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 78.250 17.505 78.570 ;
      LAYER met4 ;
        RECT 17.185 78.250 17.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 77.845 17.505 78.165 ;
      LAYER met4 ;
        RECT 17.185 77.845 17.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 77.440 17.505 77.760 ;
      LAYER met4 ;
        RECT 17.185 77.440 17.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 77.035 17.505 77.355 ;
      LAYER met4 ;
        RECT 17.185 77.035 17.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 76.630 17.505 76.950 ;
      LAYER met4 ;
        RECT 17.185 76.630 17.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 76.225 17.505 76.545 ;
      LAYER met4 ;
        RECT 17.185 76.225 17.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 75.820 17.505 76.140 ;
      LAYER met4 ;
        RECT 17.185 75.820 17.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 75.415 17.505 75.735 ;
      LAYER met4 ;
        RECT 17.185 75.415 17.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 75.010 17.505 75.330 ;
      LAYER met4 ;
        RECT 17.185 75.010 17.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 74.605 17.505 74.925 ;
      LAYER met4 ;
        RECT 17.185 74.605 17.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 74.200 17.505 74.520 ;
      LAYER met4 ;
        RECT 17.185 74.200 17.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 73.795 17.505 74.115 ;
      LAYER met4 ;
        RECT 17.185 73.795 17.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 73.390 17.505 73.710 ;
      LAYER met4 ;
        RECT 17.185 73.390 17.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 72.985 17.505 73.305 ;
      LAYER met4 ;
        RECT 17.185 72.985 17.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 72.575 17.505 72.895 ;
      LAYER met4 ;
        RECT 17.185 72.575 17.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 72.165 17.505 72.485 ;
      LAYER met4 ;
        RECT 17.185 72.165 17.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 71.755 17.505 72.075 ;
      LAYER met4 ;
        RECT 17.185 71.755 17.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 71.345 17.505 71.665 ;
      LAYER met4 ;
        RECT 17.185 71.345 17.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 70.935 17.505 71.255 ;
      LAYER met4 ;
        RECT 17.185 70.935 17.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 70.525 17.505 70.845 ;
      LAYER met4 ;
        RECT 17.185 70.525 17.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 70.115 17.505 70.435 ;
      LAYER met4 ;
        RECT 17.185 70.115 17.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 69.705 17.505 70.025 ;
      LAYER met4 ;
        RECT 17.185 69.705 17.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 69.295 17.505 69.615 ;
      LAYER met4 ;
        RECT 17.185 69.295 17.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 68.885 17.505 69.205 ;
      LAYER met4 ;
        RECT 17.185 68.885 17.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 68.475 17.505 68.795 ;
      LAYER met4 ;
        RECT 17.185 68.475 17.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.185 68.065 17.505 68.385 ;
      LAYER met4 ;
        RECT 17.185 68.065 17.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 87.815 17.185 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 87.410 17.185 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 87.005 17.185 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 86.600 17.185 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 86.195 17.185 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 85.795 17.185 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 85.395 17.185 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 84.995 17.185 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 84.595 17.185 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 84.195 17.185 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 83.795 17.185 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 83.395 17.185 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.865 82.995 17.185 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 22.160 17.090 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 21.730 17.090 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 21.300 17.090 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 20.870 17.090 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 20.440 17.090 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 20.010 17.090 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 19.580 17.090 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 19.150 17.090 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 18.720 17.090 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 18.290 17.090 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.890 17.860 17.090 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 82.300 17.105 82.620 ;
      LAYER met4 ;
        RECT 16.785 82.300 17.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 81.895 17.105 82.215 ;
      LAYER met4 ;
        RECT 16.785 81.895 17.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 81.490 17.105 81.810 ;
      LAYER met4 ;
        RECT 16.785 81.490 17.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 81.085 17.105 81.405 ;
      LAYER met4 ;
        RECT 16.785 81.085 17.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 80.680 17.105 81.000 ;
      LAYER met4 ;
        RECT 16.785 80.680 17.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 80.275 17.105 80.595 ;
      LAYER met4 ;
        RECT 16.785 80.275 17.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 79.870 17.105 80.190 ;
      LAYER met4 ;
        RECT 16.785 79.870 17.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 79.465 17.105 79.785 ;
      LAYER met4 ;
        RECT 16.785 79.465 17.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 79.060 17.105 79.380 ;
      LAYER met4 ;
        RECT 16.785 79.060 17.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 78.655 17.105 78.975 ;
      LAYER met4 ;
        RECT 16.785 78.655 17.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 78.250 17.105 78.570 ;
      LAYER met4 ;
        RECT 16.785 78.250 17.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 77.845 17.105 78.165 ;
      LAYER met4 ;
        RECT 16.785 77.845 17.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 77.440 17.105 77.760 ;
      LAYER met4 ;
        RECT 16.785 77.440 17.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 77.035 17.105 77.355 ;
      LAYER met4 ;
        RECT 16.785 77.035 17.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 76.630 17.105 76.950 ;
      LAYER met4 ;
        RECT 16.785 76.630 17.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 76.225 17.105 76.545 ;
      LAYER met4 ;
        RECT 16.785 76.225 17.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 75.820 17.105 76.140 ;
      LAYER met4 ;
        RECT 16.785 75.820 17.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 75.415 17.105 75.735 ;
      LAYER met4 ;
        RECT 16.785 75.415 17.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 75.010 17.105 75.330 ;
      LAYER met4 ;
        RECT 16.785 75.010 17.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 74.605 17.105 74.925 ;
      LAYER met4 ;
        RECT 16.785 74.605 17.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 74.200 17.105 74.520 ;
      LAYER met4 ;
        RECT 16.785 74.200 17.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 73.795 17.105 74.115 ;
      LAYER met4 ;
        RECT 16.785 73.795 17.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 73.390 17.105 73.710 ;
      LAYER met4 ;
        RECT 16.785 73.390 17.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 72.985 17.105 73.305 ;
      LAYER met4 ;
        RECT 16.785 72.985 17.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 72.575 17.105 72.895 ;
      LAYER met4 ;
        RECT 16.785 72.575 17.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 72.165 17.105 72.485 ;
      LAYER met4 ;
        RECT 16.785 72.165 17.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 71.755 17.105 72.075 ;
      LAYER met4 ;
        RECT 16.785 71.755 17.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 71.345 17.105 71.665 ;
      LAYER met4 ;
        RECT 16.785 71.345 17.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 70.935 17.105 71.255 ;
      LAYER met4 ;
        RECT 16.785 70.935 17.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 70.525 17.105 70.845 ;
      LAYER met4 ;
        RECT 16.785 70.525 17.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 70.115 17.105 70.435 ;
      LAYER met4 ;
        RECT 16.785 70.115 17.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 69.705 17.105 70.025 ;
      LAYER met4 ;
        RECT 16.785 69.705 17.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 69.295 17.105 69.615 ;
      LAYER met4 ;
        RECT 16.785 69.295 17.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 68.885 17.105 69.205 ;
      LAYER met4 ;
        RECT 16.785 68.885 17.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 68.475 17.105 68.795 ;
      LAYER met4 ;
        RECT 16.785 68.475 17.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.785 68.065 17.105 68.385 ;
      LAYER met4 ;
        RECT 16.785 68.065 17.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 87.815 16.775 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 87.410 16.775 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 87.005 16.775 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 86.600 16.775 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 86.195 16.775 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 85.795 16.775 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 85.395 16.775 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 84.995 16.775 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 84.595 16.775 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 84.195 16.775 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 83.795 16.775 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 83.395 16.775 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.455 82.995 16.775 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 22.160 16.685 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 21.730 16.685 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 21.300 16.685 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 20.870 16.685 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 20.440 16.685 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 20.010 16.685 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 19.580 16.685 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 19.150 16.685 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 18.720 16.685 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 18.290 16.685 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.485 17.860 16.685 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.420 89.205 16.740 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.420 88.785 16.740 89.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.420 88.370 16.740 88.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 82.300 16.705 82.620 ;
      LAYER met4 ;
        RECT 16.385 82.300 16.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 81.895 16.705 82.215 ;
      LAYER met4 ;
        RECT 16.385 81.895 16.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 81.490 16.705 81.810 ;
      LAYER met4 ;
        RECT 16.385 81.490 16.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 81.085 16.705 81.405 ;
      LAYER met4 ;
        RECT 16.385 81.085 16.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 80.680 16.705 81.000 ;
      LAYER met4 ;
        RECT 16.385 80.680 16.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 80.275 16.705 80.595 ;
      LAYER met4 ;
        RECT 16.385 80.275 16.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 79.870 16.705 80.190 ;
      LAYER met4 ;
        RECT 16.385 79.870 16.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 79.465 16.705 79.785 ;
      LAYER met4 ;
        RECT 16.385 79.465 16.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 79.060 16.705 79.380 ;
      LAYER met4 ;
        RECT 16.385 79.060 16.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 78.655 16.705 78.975 ;
      LAYER met4 ;
        RECT 16.385 78.655 16.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 78.250 16.705 78.570 ;
      LAYER met4 ;
        RECT 16.385 78.250 16.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 77.845 16.705 78.165 ;
      LAYER met4 ;
        RECT 16.385 77.845 16.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 77.440 16.705 77.760 ;
      LAYER met4 ;
        RECT 16.385 77.440 16.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 77.035 16.705 77.355 ;
      LAYER met4 ;
        RECT 16.385 77.035 16.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 76.630 16.705 76.950 ;
      LAYER met4 ;
        RECT 16.385 76.630 16.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 76.225 16.705 76.545 ;
      LAYER met4 ;
        RECT 16.385 76.225 16.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 75.820 16.705 76.140 ;
      LAYER met4 ;
        RECT 16.385 75.820 16.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 75.415 16.705 75.735 ;
      LAYER met4 ;
        RECT 16.385 75.415 16.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 75.010 16.705 75.330 ;
      LAYER met4 ;
        RECT 16.385 75.010 16.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 74.605 16.705 74.925 ;
      LAYER met4 ;
        RECT 16.385 74.605 16.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 74.200 16.705 74.520 ;
      LAYER met4 ;
        RECT 16.385 74.200 16.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 73.795 16.705 74.115 ;
      LAYER met4 ;
        RECT 16.385 73.795 16.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 73.390 16.705 73.710 ;
      LAYER met4 ;
        RECT 16.385 73.390 16.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 72.985 16.705 73.305 ;
      LAYER met4 ;
        RECT 16.385 72.985 16.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 72.575 16.705 72.895 ;
      LAYER met4 ;
        RECT 16.385 72.575 16.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 72.165 16.705 72.485 ;
      LAYER met4 ;
        RECT 16.385 72.165 16.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 71.755 16.705 72.075 ;
      LAYER met4 ;
        RECT 16.385 71.755 16.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 71.345 16.705 71.665 ;
      LAYER met4 ;
        RECT 16.385 71.345 16.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 70.935 16.705 71.255 ;
      LAYER met4 ;
        RECT 16.385 70.935 16.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 70.525 16.705 70.845 ;
      LAYER met4 ;
        RECT 16.385 70.525 16.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 70.115 16.705 70.435 ;
      LAYER met4 ;
        RECT 16.385 70.115 16.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 69.705 16.705 70.025 ;
      LAYER met4 ;
        RECT 16.385 69.705 16.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 69.295 16.705 69.615 ;
      LAYER met4 ;
        RECT 16.385 69.295 16.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 68.885 16.705 69.205 ;
      LAYER met4 ;
        RECT 16.385 68.885 16.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 68.475 16.705 68.795 ;
      LAYER met4 ;
        RECT 16.385 68.475 16.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.385 68.065 16.705 68.385 ;
      LAYER met4 ;
        RECT 16.385 68.065 16.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 87.815 16.365 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 87.410 16.365 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 87.005 16.365 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 86.600 16.365 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 86.195 16.365 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 85.795 16.365 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 85.395 16.365 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 84.995 16.365 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 84.595 16.365 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 84.195 16.365 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 83.795 16.365 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 83.395 16.365 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 82.995 16.365 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 22.160 16.280 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 21.730 16.280 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 21.300 16.280 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 20.870 16.280 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 20.440 16.280 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 20.010 16.280 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 19.580 16.280 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 19.150 16.280 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 18.720 16.280 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 18.290 16.280 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.080 17.860 16.280 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 82.300 16.305 82.620 ;
      LAYER met4 ;
        RECT 15.985 82.300 16.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 81.895 16.305 82.215 ;
      LAYER met4 ;
        RECT 15.985 81.895 16.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 81.490 16.305 81.810 ;
      LAYER met4 ;
        RECT 15.985 81.490 16.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 81.085 16.305 81.405 ;
      LAYER met4 ;
        RECT 15.985 81.085 16.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 80.680 16.305 81.000 ;
      LAYER met4 ;
        RECT 15.985 80.680 16.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 80.275 16.305 80.595 ;
      LAYER met4 ;
        RECT 15.985 80.275 16.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 79.870 16.305 80.190 ;
      LAYER met4 ;
        RECT 15.985 79.870 16.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 79.465 16.305 79.785 ;
      LAYER met4 ;
        RECT 15.985 79.465 16.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 79.060 16.305 79.380 ;
      LAYER met4 ;
        RECT 15.985 79.060 16.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 78.655 16.305 78.975 ;
      LAYER met4 ;
        RECT 15.985 78.655 16.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 78.250 16.305 78.570 ;
      LAYER met4 ;
        RECT 15.985 78.250 16.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 77.845 16.305 78.165 ;
      LAYER met4 ;
        RECT 15.985 77.845 16.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 77.440 16.305 77.760 ;
      LAYER met4 ;
        RECT 15.985 77.440 16.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 77.035 16.305 77.355 ;
      LAYER met4 ;
        RECT 15.985 77.035 16.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 76.630 16.305 76.950 ;
      LAYER met4 ;
        RECT 15.985 76.630 16.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 76.225 16.305 76.545 ;
      LAYER met4 ;
        RECT 15.985 76.225 16.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 75.820 16.305 76.140 ;
      LAYER met4 ;
        RECT 15.985 75.820 16.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 75.415 16.305 75.735 ;
      LAYER met4 ;
        RECT 15.985 75.415 16.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 75.010 16.305 75.330 ;
      LAYER met4 ;
        RECT 15.985 75.010 16.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 74.605 16.305 74.925 ;
      LAYER met4 ;
        RECT 15.985 74.605 16.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 74.200 16.305 74.520 ;
      LAYER met4 ;
        RECT 15.985 74.200 16.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 73.795 16.305 74.115 ;
      LAYER met4 ;
        RECT 15.985 73.795 16.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 73.390 16.305 73.710 ;
      LAYER met4 ;
        RECT 15.985 73.390 16.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 72.985 16.305 73.305 ;
      LAYER met4 ;
        RECT 15.985 72.985 16.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 72.575 16.305 72.895 ;
      LAYER met4 ;
        RECT 15.985 72.575 16.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 72.165 16.305 72.485 ;
      LAYER met4 ;
        RECT 15.985 72.165 16.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 71.755 16.305 72.075 ;
      LAYER met4 ;
        RECT 15.985 71.755 16.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 71.345 16.305 71.665 ;
      LAYER met4 ;
        RECT 15.985 71.345 16.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 70.935 16.305 71.255 ;
      LAYER met4 ;
        RECT 15.985 70.935 16.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 70.525 16.305 70.845 ;
      LAYER met4 ;
        RECT 15.985 70.525 16.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 70.115 16.305 70.435 ;
      LAYER met4 ;
        RECT 15.985 70.115 16.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 69.705 16.305 70.025 ;
      LAYER met4 ;
        RECT 15.985 69.705 16.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 69.295 16.305 69.615 ;
      LAYER met4 ;
        RECT 15.985 69.295 16.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 68.885 16.305 69.205 ;
      LAYER met4 ;
        RECT 15.985 68.885 16.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 68.475 16.305 68.795 ;
      LAYER met4 ;
        RECT 15.985 68.475 16.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 68.065 16.305 68.385 ;
      LAYER met4 ;
        RECT 15.985 68.065 16.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920 90.495 16.240 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920 90.065 16.240 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920 89.635 16.240 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920 89.205 16.240 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920 88.775 16.240 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.920 88.350 16.240 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 87.815 15.955 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 87.410 15.955 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 87.005 15.955 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 86.600 15.955 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 86.195 15.955 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 85.795 15.955 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 85.395 15.955 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 84.995 15.955 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 84.595 15.955 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 84.195 15.955 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 83.795 15.955 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 83.395 15.955 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.635 82.995 15.955 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 22.160 15.875 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 21.730 15.875 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 21.300 15.875 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 20.870 15.875 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 20.440 15.875 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 20.010 15.875 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 19.580 15.875 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 19.150 15.875 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 18.720 15.875 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 18.290 15.875 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.675 17.860 15.875 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 82.300 15.905 82.620 ;
      LAYER met4 ;
        RECT 15.585 82.300 15.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 81.895 15.905 82.215 ;
      LAYER met4 ;
        RECT 15.585 81.895 15.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 81.490 15.905 81.810 ;
      LAYER met4 ;
        RECT 15.585 81.490 15.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 81.085 15.905 81.405 ;
      LAYER met4 ;
        RECT 15.585 81.085 15.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 80.680 15.905 81.000 ;
      LAYER met4 ;
        RECT 15.585 80.680 15.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 80.275 15.905 80.595 ;
      LAYER met4 ;
        RECT 15.585 80.275 15.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 79.870 15.905 80.190 ;
      LAYER met4 ;
        RECT 15.585 79.870 15.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 79.465 15.905 79.785 ;
      LAYER met4 ;
        RECT 15.585 79.465 15.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 79.060 15.905 79.380 ;
      LAYER met4 ;
        RECT 15.585 79.060 15.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 78.655 15.905 78.975 ;
      LAYER met4 ;
        RECT 15.585 78.655 15.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 78.250 15.905 78.570 ;
      LAYER met4 ;
        RECT 15.585 78.250 15.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 77.845 15.905 78.165 ;
      LAYER met4 ;
        RECT 15.585 77.845 15.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 77.440 15.905 77.760 ;
      LAYER met4 ;
        RECT 15.585 77.440 15.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 77.035 15.905 77.355 ;
      LAYER met4 ;
        RECT 15.585 77.035 15.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 76.630 15.905 76.950 ;
      LAYER met4 ;
        RECT 15.585 76.630 15.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 76.225 15.905 76.545 ;
      LAYER met4 ;
        RECT 15.585 76.225 15.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 75.820 15.905 76.140 ;
      LAYER met4 ;
        RECT 15.585 75.820 15.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 75.415 15.905 75.735 ;
      LAYER met4 ;
        RECT 15.585 75.415 15.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 75.010 15.905 75.330 ;
      LAYER met4 ;
        RECT 15.585 75.010 15.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 74.605 15.905 74.925 ;
      LAYER met4 ;
        RECT 15.585 74.605 15.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 74.200 15.905 74.520 ;
      LAYER met4 ;
        RECT 15.585 74.200 15.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 73.795 15.905 74.115 ;
      LAYER met4 ;
        RECT 15.585 73.795 15.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 73.390 15.905 73.710 ;
      LAYER met4 ;
        RECT 15.585 73.390 15.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 72.985 15.905 73.305 ;
      LAYER met4 ;
        RECT 15.585 72.985 15.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 72.575 15.905 72.895 ;
      LAYER met4 ;
        RECT 15.585 72.575 15.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 72.165 15.905 72.485 ;
      LAYER met4 ;
        RECT 15.585 72.165 15.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 71.755 15.905 72.075 ;
      LAYER met4 ;
        RECT 15.585 71.755 15.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 71.345 15.905 71.665 ;
      LAYER met4 ;
        RECT 15.585 71.345 15.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 70.935 15.905 71.255 ;
      LAYER met4 ;
        RECT 15.585 70.935 15.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 70.525 15.905 70.845 ;
      LAYER met4 ;
        RECT 15.585 70.525 15.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 70.115 15.905 70.435 ;
      LAYER met4 ;
        RECT 15.585 70.115 15.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 69.705 15.905 70.025 ;
      LAYER met4 ;
        RECT 15.585 69.705 15.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 69.295 15.905 69.615 ;
      LAYER met4 ;
        RECT 15.585 69.295 15.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 68.885 15.905 69.205 ;
      LAYER met4 ;
        RECT 15.585 68.885 15.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 68.475 15.905 68.795 ;
      LAYER met4 ;
        RECT 15.585 68.475 15.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.585 68.065 15.905 68.385 ;
      LAYER met4 ;
        RECT 15.585 68.065 15.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510 90.495 15.830 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510 90.065 15.830 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510 89.635 15.830 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510 89.205 15.830 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510 88.775 15.830 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.510 88.350 15.830 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 87.815 15.545 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 87.410 15.545 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 87.005 15.545 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 86.600 15.545 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 86.195 15.545 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 85.795 15.545 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 85.395 15.545 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 84.995 15.545 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 84.595 15.545 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 84.195 15.545 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 83.795 15.545 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 83.395 15.545 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.225 82.995 15.545 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 22.160 15.470 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 21.730 15.470 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 21.300 15.470 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 20.870 15.470 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 20.440 15.470 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 20.010 15.470 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 19.580 15.470 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 19.150 15.470 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 18.720 15.470 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 18.290 15.470 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.270 17.860 15.470 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 82.300 15.505 82.620 ;
      LAYER met4 ;
        RECT 15.185 82.300 15.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 81.895 15.505 82.215 ;
      LAYER met4 ;
        RECT 15.185 81.895 15.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 81.490 15.505 81.810 ;
      LAYER met4 ;
        RECT 15.185 81.490 15.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 81.085 15.505 81.405 ;
      LAYER met4 ;
        RECT 15.185 81.085 15.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 80.680 15.505 81.000 ;
      LAYER met4 ;
        RECT 15.185 80.680 15.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 80.275 15.505 80.595 ;
      LAYER met4 ;
        RECT 15.185 80.275 15.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 79.870 15.505 80.190 ;
      LAYER met4 ;
        RECT 15.185 79.870 15.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 79.465 15.505 79.785 ;
      LAYER met4 ;
        RECT 15.185 79.465 15.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 79.060 15.505 79.380 ;
      LAYER met4 ;
        RECT 15.185 79.060 15.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 78.655 15.505 78.975 ;
      LAYER met4 ;
        RECT 15.185 78.655 15.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 78.250 15.505 78.570 ;
      LAYER met4 ;
        RECT 15.185 78.250 15.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 77.845 15.505 78.165 ;
      LAYER met4 ;
        RECT 15.185 77.845 15.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 77.440 15.505 77.760 ;
      LAYER met4 ;
        RECT 15.185 77.440 15.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 77.035 15.505 77.355 ;
      LAYER met4 ;
        RECT 15.185 77.035 15.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 76.630 15.505 76.950 ;
      LAYER met4 ;
        RECT 15.185 76.630 15.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 76.225 15.505 76.545 ;
      LAYER met4 ;
        RECT 15.185 76.225 15.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 75.820 15.505 76.140 ;
      LAYER met4 ;
        RECT 15.185 75.820 15.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 75.415 15.505 75.735 ;
      LAYER met4 ;
        RECT 15.185 75.415 15.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 75.010 15.505 75.330 ;
      LAYER met4 ;
        RECT 15.185 75.010 15.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 74.605 15.505 74.925 ;
      LAYER met4 ;
        RECT 15.185 74.605 15.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 74.200 15.505 74.520 ;
      LAYER met4 ;
        RECT 15.185 74.200 15.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 73.795 15.505 74.115 ;
      LAYER met4 ;
        RECT 15.185 73.795 15.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 73.390 15.505 73.710 ;
      LAYER met4 ;
        RECT 15.185 73.390 15.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 72.985 15.505 73.305 ;
      LAYER met4 ;
        RECT 15.185 72.985 15.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 72.575 15.505 72.895 ;
      LAYER met4 ;
        RECT 15.185 72.575 15.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 72.165 15.505 72.485 ;
      LAYER met4 ;
        RECT 15.185 72.165 15.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 71.755 15.505 72.075 ;
      LAYER met4 ;
        RECT 15.185 71.755 15.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 71.345 15.505 71.665 ;
      LAYER met4 ;
        RECT 15.185 71.345 15.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 70.935 15.505 71.255 ;
      LAYER met4 ;
        RECT 15.185 70.935 15.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 70.525 15.505 70.845 ;
      LAYER met4 ;
        RECT 15.185 70.525 15.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 70.115 15.505 70.435 ;
      LAYER met4 ;
        RECT 15.185 70.115 15.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 69.705 15.505 70.025 ;
      LAYER met4 ;
        RECT 15.185 69.705 15.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 69.295 15.505 69.615 ;
      LAYER met4 ;
        RECT 15.185 69.295 15.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 68.885 15.505 69.205 ;
      LAYER met4 ;
        RECT 15.185 68.885 15.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 68.475 15.505 68.795 ;
      LAYER met4 ;
        RECT 15.185 68.475 15.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.185 68.065 15.505 68.385 ;
      LAYER met4 ;
        RECT 15.185 68.065 15.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100 90.495 15.420 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100 90.065 15.420 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100 89.635 15.420 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100 89.205 15.420 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100 88.775 15.420 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.100 88.350 15.420 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.040 91.385 15.360 91.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.040 90.955 15.360 91.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 87.815 15.135 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 87.410 15.135 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 87.005 15.135 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 86.600 15.135 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 86.195 15.135 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 85.795 15.135 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 85.395 15.135 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 84.995 15.135 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 84.595 15.135 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 84.195 15.135 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 83.795 15.135 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 83.395 15.135 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.815 82.995 15.135 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 22.160 15.065 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 21.730 15.065 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 21.300 15.065 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 20.870 15.065 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 20.440 15.065 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 20.010 15.065 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 19.580 15.065 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 19.150 15.065 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 18.720 15.065 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 18.290 15.065 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.865 17.860 15.065 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 82.300 15.105 82.620 ;
      LAYER met4 ;
        RECT 14.785 82.300 15.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 81.895 15.105 82.215 ;
      LAYER met4 ;
        RECT 14.785 81.895 15.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 81.490 15.105 81.810 ;
      LAYER met4 ;
        RECT 14.785 81.490 15.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 81.085 15.105 81.405 ;
      LAYER met4 ;
        RECT 14.785 81.085 15.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 80.680 15.105 81.000 ;
      LAYER met4 ;
        RECT 14.785 80.680 15.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 80.275 15.105 80.595 ;
      LAYER met4 ;
        RECT 14.785 80.275 15.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 79.870 15.105 80.190 ;
      LAYER met4 ;
        RECT 14.785 79.870 15.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 79.465 15.105 79.785 ;
      LAYER met4 ;
        RECT 14.785 79.465 15.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 79.060 15.105 79.380 ;
      LAYER met4 ;
        RECT 14.785 79.060 15.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 78.655 15.105 78.975 ;
      LAYER met4 ;
        RECT 14.785 78.655 15.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 78.250 15.105 78.570 ;
      LAYER met4 ;
        RECT 14.785 78.250 15.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 77.845 15.105 78.165 ;
      LAYER met4 ;
        RECT 14.785 77.845 15.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 77.440 15.105 77.760 ;
      LAYER met4 ;
        RECT 14.785 77.440 15.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 77.035 15.105 77.355 ;
      LAYER met4 ;
        RECT 14.785 77.035 15.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 76.630 15.105 76.950 ;
      LAYER met4 ;
        RECT 14.785 76.630 15.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 76.225 15.105 76.545 ;
      LAYER met4 ;
        RECT 14.785 76.225 15.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 75.820 15.105 76.140 ;
      LAYER met4 ;
        RECT 14.785 75.820 15.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 75.415 15.105 75.735 ;
      LAYER met4 ;
        RECT 14.785 75.415 15.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 75.010 15.105 75.330 ;
      LAYER met4 ;
        RECT 14.785 75.010 15.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 74.605 15.105 74.925 ;
      LAYER met4 ;
        RECT 14.785 74.605 15.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 74.200 15.105 74.520 ;
      LAYER met4 ;
        RECT 14.785 74.200 15.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 73.795 15.105 74.115 ;
      LAYER met4 ;
        RECT 14.785 73.795 15.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 73.390 15.105 73.710 ;
      LAYER met4 ;
        RECT 14.785 73.390 15.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 72.985 15.105 73.305 ;
      LAYER met4 ;
        RECT 14.785 72.985 15.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 72.575 15.105 72.895 ;
      LAYER met4 ;
        RECT 14.785 72.575 15.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 72.165 15.105 72.485 ;
      LAYER met4 ;
        RECT 14.785 72.165 15.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 71.755 15.105 72.075 ;
      LAYER met4 ;
        RECT 14.785 71.755 15.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 71.345 15.105 71.665 ;
      LAYER met4 ;
        RECT 14.785 71.345 15.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 70.935 15.105 71.255 ;
      LAYER met4 ;
        RECT 14.785 70.935 15.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 70.525 15.105 70.845 ;
      LAYER met4 ;
        RECT 14.785 70.525 15.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 70.115 15.105 70.435 ;
      LAYER met4 ;
        RECT 14.785 70.115 15.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 69.705 15.105 70.025 ;
      LAYER met4 ;
        RECT 14.785 69.705 15.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 69.295 15.105 69.615 ;
      LAYER met4 ;
        RECT 14.785 69.295 15.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 68.885 15.105 69.205 ;
      LAYER met4 ;
        RECT 14.785 68.885 15.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 68.475 15.105 68.795 ;
      LAYER met4 ;
        RECT 14.785 68.475 15.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.785 68.065 15.105 68.385 ;
      LAYER met4 ;
        RECT 14.785 68.065 15.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690 90.495 15.010 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690 90.065 15.010 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690 89.635 15.010 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690 89.205 15.010 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690 88.775 15.010 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.690 88.350 15.010 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 87.815 14.725 88.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 87.410 14.725 87.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 87.005 14.725 87.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 86.600 14.725 86.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 86.195 14.725 86.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 85.795 14.725 86.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 85.395 14.725 85.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 84.995 14.725 85.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 84.595 14.725 84.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 84.195 14.725 84.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 83.795 14.725 84.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 83.395 14.725 83.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.405 82.995 14.725 83.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 22.160 14.660 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 21.730 14.660 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 21.300 14.660 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 20.870 14.660 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 20.440 14.660 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 20.010 14.660 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 19.580 14.660 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 19.150 14.660 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 18.720 14.660 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 18.290 14.660 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.460 17.860 14.660 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 82.300 14.705 82.620 ;
      LAYER met4 ;
        RECT 14.385 82.300 14.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 81.895 14.705 82.215 ;
      LAYER met4 ;
        RECT 14.385 81.895 14.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 81.490 14.705 81.810 ;
      LAYER met4 ;
        RECT 14.385 81.490 14.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 81.085 14.705 81.405 ;
      LAYER met4 ;
        RECT 14.385 81.085 14.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 80.680 14.705 81.000 ;
      LAYER met4 ;
        RECT 14.385 80.680 14.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 80.275 14.705 80.595 ;
      LAYER met4 ;
        RECT 14.385 80.275 14.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 79.870 14.705 80.190 ;
      LAYER met4 ;
        RECT 14.385 79.870 14.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 79.465 14.705 79.785 ;
      LAYER met4 ;
        RECT 14.385 79.465 14.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 79.060 14.705 79.380 ;
      LAYER met4 ;
        RECT 14.385 79.060 14.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 78.655 14.705 78.975 ;
      LAYER met4 ;
        RECT 14.385 78.655 14.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 78.250 14.705 78.570 ;
      LAYER met4 ;
        RECT 14.385 78.250 14.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 77.845 14.705 78.165 ;
      LAYER met4 ;
        RECT 14.385 77.845 14.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 77.440 14.705 77.760 ;
      LAYER met4 ;
        RECT 14.385 77.440 14.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 77.035 14.705 77.355 ;
      LAYER met4 ;
        RECT 14.385 77.035 14.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 76.630 14.705 76.950 ;
      LAYER met4 ;
        RECT 14.385 76.630 14.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 76.225 14.705 76.545 ;
      LAYER met4 ;
        RECT 14.385 76.225 14.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 75.820 14.705 76.140 ;
      LAYER met4 ;
        RECT 14.385 75.820 14.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 75.415 14.705 75.735 ;
      LAYER met4 ;
        RECT 14.385 75.415 14.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 75.010 14.705 75.330 ;
      LAYER met4 ;
        RECT 14.385 75.010 14.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 74.605 14.705 74.925 ;
      LAYER met4 ;
        RECT 14.385 74.605 14.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 74.200 14.705 74.520 ;
      LAYER met4 ;
        RECT 14.385 74.200 14.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 73.795 14.705 74.115 ;
      LAYER met4 ;
        RECT 14.385 73.795 14.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 73.390 14.705 73.710 ;
      LAYER met4 ;
        RECT 14.385 73.390 14.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 72.985 14.705 73.305 ;
      LAYER met4 ;
        RECT 14.385 72.985 14.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 72.575 14.705 72.895 ;
      LAYER met4 ;
        RECT 14.385 72.575 14.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 72.165 14.705 72.485 ;
      LAYER met4 ;
        RECT 14.385 72.165 14.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 71.755 14.705 72.075 ;
      LAYER met4 ;
        RECT 14.385 71.755 14.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 71.345 14.705 71.665 ;
      LAYER met4 ;
        RECT 14.385 71.345 14.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 70.935 14.705 71.255 ;
      LAYER met4 ;
        RECT 14.385 70.935 14.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 70.525 14.705 70.845 ;
      LAYER met4 ;
        RECT 14.385 70.525 14.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 70.115 14.705 70.435 ;
      LAYER met4 ;
        RECT 14.385 70.115 14.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 69.705 14.705 70.025 ;
      LAYER met4 ;
        RECT 14.385 69.705 14.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 69.295 14.705 69.615 ;
      LAYER met4 ;
        RECT 14.385 69.295 14.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 68.885 14.705 69.205 ;
      LAYER met4 ;
        RECT 14.385 68.885 14.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 68.475 14.705 68.795 ;
      LAYER met4 ;
        RECT 14.385 68.475 14.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 68.065 14.705 68.385 ;
      LAYER met4 ;
        RECT 14.385 68.065 14.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280 90.495 14.600 90.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280 90.065 14.600 90.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280 89.635 14.600 89.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280 89.205 14.600 89.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280 88.775 14.600 89.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.280 88.350 14.600 88.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.260 91.385 14.580 91.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.260 90.955 14.580 91.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 22.160 14.255 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 21.730 14.255 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 21.300 14.255 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 20.870 14.255 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 20.440 14.255 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 20.010 14.255 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 19.580 14.255 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 19.150 14.255 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 18.720 14.255 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 18.290 14.255 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.055 17.860 14.255 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 82.300 14.305 82.620 ;
      LAYER met4 ;
        RECT 13.985 82.300 14.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 81.895 14.305 82.215 ;
      LAYER met4 ;
        RECT 13.985 81.895 14.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 81.490 14.305 81.810 ;
      LAYER met4 ;
        RECT 13.985 81.490 14.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 81.085 14.305 81.405 ;
      LAYER met4 ;
        RECT 13.985 81.085 14.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 80.680 14.305 81.000 ;
      LAYER met4 ;
        RECT 13.985 80.680 14.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 80.275 14.305 80.595 ;
      LAYER met4 ;
        RECT 13.985 80.275 14.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 79.870 14.305 80.190 ;
      LAYER met4 ;
        RECT 13.985 79.870 14.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 79.465 14.305 79.785 ;
      LAYER met4 ;
        RECT 13.985 79.465 14.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 79.060 14.305 79.380 ;
      LAYER met4 ;
        RECT 13.985 79.060 14.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 78.655 14.305 78.975 ;
      LAYER met4 ;
        RECT 13.985 78.655 14.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 78.250 14.305 78.570 ;
      LAYER met4 ;
        RECT 13.985 78.250 14.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 77.845 14.305 78.165 ;
      LAYER met4 ;
        RECT 13.985 77.845 14.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 77.440 14.305 77.760 ;
      LAYER met4 ;
        RECT 13.985 77.440 14.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 77.035 14.305 77.355 ;
      LAYER met4 ;
        RECT 13.985 77.035 14.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 76.630 14.305 76.950 ;
      LAYER met4 ;
        RECT 13.985 76.630 14.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 76.225 14.305 76.545 ;
      LAYER met4 ;
        RECT 13.985 76.225 14.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 75.820 14.305 76.140 ;
      LAYER met4 ;
        RECT 13.985 75.820 14.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 75.415 14.305 75.735 ;
      LAYER met4 ;
        RECT 13.985 75.415 14.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 75.010 14.305 75.330 ;
      LAYER met4 ;
        RECT 13.985 75.010 14.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 74.605 14.305 74.925 ;
      LAYER met4 ;
        RECT 13.985 74.605 14.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 74.200 14.305 74.520 ;
      LAYER met4 ;
        RECT 13.985 74.200 14.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 73.795 14.305 74.115 ;
      LAYER met4 ;
        RECT 13.985 73.795 14.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 73.390 14.305 73.710 ;
      LAYER met4 ;
        RECT 13.985 73.390 14.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 72.985 14.305 73.305 ;
      LAYER met4 ;
        RECT 13.985 72.985 14.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 72.575 14.305 72.895 ;
      LAYER met4 ;
        RECT 13.985 72.575 14.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 72.165 14.305 72.485 ;
      LAYER met4 ;
        RECT 13.985 72.165 14.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 71.755 14.305 72.075 ;
      LAYER met4 ;
        RECT 13.985 71.755 14.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 71.345 14.305 71.665 ;
      LAYER met4 ;
        RECT 13.985 71.345 14.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 70.935 14.305 71.255 ;
      LAYER met4 ;
        RECT 13.985 70.935 14.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 70.525 14.305 70.845 ;
      LAYER met4 ;
        RECT 13.985 70.525 14.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 70.115 14.305 70.435 ;
      LAYER met4 ;
        RECT 13.985 70.115 14.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 69.705 14.305 70.025 ;
      LAYER met4 ;
        RECT 13.985 69.705 14.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 69.295 14.305 69.615 ;
      LAYER met4 ;
        RECT 13.985 69.295 14.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 68.885 14.305 69.205 ;
      LAYER met4 ;
        RECT 13.985 68.885 14.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 68.475 14.305 68.795 ;
      LAYER met4 ;
        RECT 13.985 68.475 14.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 68.065 14.305 68.385 ;
      LAYER met4 ;
        RECT 13.985 68.065 14.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 92.635 14.100 92.955 ;
      LAYER met4 ;
        RECT 13.780 92.635 14.100 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 92.225 14.100 92.545 ;
      LAYER met4 ;
        RECT 13.780 92.225 14.100 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 91.815 14.100 92.135 ;
      LAYER met4 ;
        RECT 13.780 91.815 14.100 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 91.405 14.100 91.725 ;
      LAYER met4 ;
        RECT 13.780 91.405 14.100 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 90.995 14.100 91.315 ;
      LAYER met4 ;
        RECT 13.780 90.995 14.100 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 90.585 14.100 90.905 ;
      LAYER met4 ;
        RECT 13.780 90.585 14.100 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 90.175 14.100 90.495 ;
      LAYER met4 ;
        RECT 13.780 90.175 14.100 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 89.765 14.100 90.085 ;
      LAYER met4 ;
        RECT 13.780 89.765 14.100 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 89.355 14.100 89.675 ;
      LAYER met4 ;
        RECT 13.780 89.355 14.100 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 88.945 14.100 89.265 ;
      LAYER met4 ;
        RECT 13.780 88.945 14.100 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 88.535 14.100 88.855 ;
      LAYER met4 ;
        RECT 13.780 88.535 14.100 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 88.125 14.100 88.445 ;
      LAYER met4 ;
        RECT 13.780 88.125 14.100 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 87.715 14.100 88.035 ;
      LAYER met4 ;
        RECT 13.780 87.715 14.100 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 87.305 14.100 87.625 ;
      LAYER met4 ;
        RECT 13.780 87.305 14.100 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 86.895 14.100 87.215 ;
      LAYER met4 ;
        RECT 13.780 86.895 14.100 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 86.485 14.100 86.805 ;
      LAYER met4 ;
        RECT 13.780 86.485 14.100 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 86.075 14.100 86.395 ;
      LAYER met4 ;
        RECT 13.780 86.075 14.100 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 85.665 14.100 85.985 ;
      LAYER met4 ;
        RECT 13.780 85.665 14.100 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 85.255 14.100 85.575 ;
      LAYER met4 ;
        RECT 13.780 85.255 14.100 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 84.845 14.100 85.165 ;
      LAYER met4 ;
        RECT 13.780 84.845 14.100 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 84.435 14.100 84.755 ;
      LAYER met4 ;
        RECT 13.780 84.435 14.100 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 84.025 14.100 84.345 ;
      LAYER met4 ;
        RECT 13.780 84.025 14.100 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 83.615 14.100 83.935 ;
      LAYER met4 ;
        RECT 13.780 83.615 14.100 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 83.205 14.100 83.525 ;
      LAYER met4 ;
        RECT 13.780 83.205 14.100 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.780 82.795 14.100 83.115 ;
      LAYER met4 ;
        RECT 13.780 82.795 14.100 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 22.160 13.850 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 21.730 13.850 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 21.300 13.850 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 20.870 13.850 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 20.440 13.850 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 20.010 13.850 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 19.580 13.850 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 19.150 13.850 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 18.720 13.850 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 18.290 13.850 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.650 17.860 13.850 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 82.300 13.905 82.620 ;
      LAYER met4 ;
        RECT 13.585 82.300 13.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 81.895 13.905 82.215 ;
      LAYER met4 ;
        RECT 13.585 81.895 13.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 81.490 13.905 81.810 ;
      LAYER met4 ;
        RECT 13.585 81.490 13.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 81.085 13.905 81.405 ;
      LAYER met4 ;
        RECT 13.585 81.085 13.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 80.680 13.905 81.000 ;
      LAYER met4 ;
        RECT 13.585 80.680 13.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 80.275 13.905 80.595 ;
      LAYER met4 ;
        RECT 13.585 80.275 13.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 79.870 13.905 80.190 ;
      LAYER met4 ;
        RECT 13.585 79.870 13.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 79.465 13.905 79.785 ;
      LAYER met4 ;
        RECT 13.585 79.465 13.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 79.060 13.905 79.380 ;
      LAYER met4 ;
        RECT 13.585 79.060 13.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 78.655 13.905 78.975 ;
      LAYER met4 ;
        RECT 13.585 78.655 13.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 78.250 13.905 78.570 ;
      LAYER met4 ;
        RECT 13.585 78.250 13.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 77.845 13.905 78.165 ;
      LAYER met4 ;
        RECT 13.585 77.845 13.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 77.440 13.905 77.760 ;
      LAYER met4 ;
        RECT 13.585 77.440 13.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 77.035 13.905 77.355 ;
      LAYER met4 ;
        RECT 13.585 77.035 13.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 76.630 13.905 76.950 ;
      LAYER met4 ;
        RECT 13.585 76.630 13.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 76.225 13.905 76.545 ;
      LAYER met4 ;
        RECT 13.585 76.225 13.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 75.820 13.905 76.140 ;
      LAYER met4 ;
        RECT 13.585 75.820 13.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 75.415 13.905 75.735 ;
      LAYER met4 ;
        RECT 13.585 75.415 13.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 75.010 13.905 75.330 ;
      LAYER met4 ;
        RECT 13.585 75.010 13.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 74.605 13.905 74.925 ;
      LAYER met4 ;
        RECT 13.585 74.605 13.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 74.200 13.905 74.520 ;
      LAYER met4 ;
        RECT 13.585 74.200 13.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 73.795 13.905 74.115 ;
      LAYER met4 ;
        RECT 13.585 73.795 13.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 73.390 13.905 73.710 ;
      LAYER met4 ;
        RECT 13.585 73.390 13.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 72.985 13.905 73.305 ;
      LAYER met4 ;
        RECT 13.585 72.985 13.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 72.575 13.905 72.895 ;
      LAYER met4 ;
        RECT 13.585 72.575 13.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 72.165 13.905 72.485 ;
      LAYER met4 ;
        RECT 13.585 72.165 13.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 71.755 13.905 72.075 ;
      LAYER met4 ;
        RECT 13.585 71.755 13.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 71.345 13.905 71.665 ;
      LAYER met4 ;
        RECT 13.585 71.345 13.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 70.935 13.905 71.255 ;
      LAYER met4 ;
        RECT 13.585 70.935 13.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 70.525 13.905 70.845 ;
      LAYER met4 ;
        RECT 13.585 70.525 13.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 70.115 13.905 70.435 ;
      LAYER met4 ;
        RECT 13.585 70.115 13.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 69.705 13.905 70.025 ;
      LAYER met4 ;
        RECT 13.585 69.705 13.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 69.295 13.905 69.615 ;
      LAYER met4 ;
        RECT 13.585 69.295 13.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 68.885 13.905 69.205 ;
      LAYER met4 ;
        RECT 13.585 68.885 13.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 68.475 13.905 68.795 ;
      LAYER met4 ;
        RECT 13.585 68.475 13.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.585 68.065 13.905 68.385 ;
      LAYER met4 ;
        RECT 13.585 68.065 13.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 92.635 13.695 92.955 ;
      LAYER met4 ;
        RECT 13.375 92.635 13.695 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 92.225 13.695 92.545 ;
      LAYER met4 ;
        RECT 13.375 92.225 13.695 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 91.815 13.695 92.135 ;
      LAYER met4 ;
        RECT 13.375 91.815 13.695 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 91.405 13.695 91.725 ;
      LAYER met4 ;
        RECT 13.375 91.405 13.695 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 90.995 13.695 91.315 ;
      LAYER met4 ;
        RECT 13.375 90.995 13.695 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 90.585 13.695 90.905 ;
      LAYER met4 ;
        RECT 13.375 90.585 13.695 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 90.175 13.695 90.495 ;
      LAYER met4 ;
        RECT 13.375 90.175 13.695 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 89.765 13.695 90.085 ;
      LAYER met4 ;
        RECT 13.375 89.765 13.695 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 89.355 13.695 89.675 ;
      LAYER met4 ;
        RECT 13.375 89.355 13.695 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 88.945 13.695 89.265 ;
      LAYER met4 ;
        RECT 13.375 88.945 13.695 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 88.535 13.695 88.855 ;
      LAYER met4 ;
        RECT 13.375 88.535 13.695 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 88.125 13.695 88.445 ;
      LAYER met4 ;
        RECT 13.375 88.125 13.695 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 87.715 13.695 88.035 ;
      LAYER met4 ;
        RECT 13.375 87.715 13.695 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 87.305 13.695 87.625 ;
      LAYER met4 ;
        RECT 13.375 87.305 13.695 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 86.895 13.695 87.215 ;
      LAYER met4 ;
        RECT 13.375 86.895 13.695 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 86.485 13.695 86.805 ;
      LAYER met4 ;
        RECT 13.375 86.485 13.695 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 86.075 13.695 86.395 ;
      LAYER met4 ;
        RECT 13.375 86.075 13.695 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 85.665 13.695 85.985 ;
      LAYER met4 ;
        RECT 13.375 85.665 13.695 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 85.255 13.695 85.575 ;
      LAYER met4 ;
        RECT 13.375 85.255 13.695 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 84.845 13.695 85.165 ;
      LAYER met4 ;
        RECT 13.375 84.845 13.695 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 84.435 13.695 84.755 ;
      LAYER met4 ;
        RECT 13.375 84.435 13.695 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 84.025 13.695 84.345 ;
      LAYER met4 ;
        RECT 13.375 84.025 13.695 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 83.615 13.695 83.935 ;
      LAYER met4 ;
        RECT 13.375 83.615 13.695 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 83.205 13.695 83.525 ;
      LAYER met4 ;
        RECT 13.375 83.205 13.695 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.375 82.795 13.695 83.115 ;
      LAYER met4 ;
        RECT 13.375 82.795 13.695 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 82.300 13.505 82.620 ;
      LAYER met4 ;
        RECT 13.185 82.300 13.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 81.895 13.505 82.215 ;
      LAYER met4 ;
        RECT 13.185 81.895 13.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 81.490 13.505 81.810 ;
      LAYER met4 ;
        RECT 13.185 81.490 13.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 81.085 13.505 81.405 ;
      LAYER met4 ;
        RECT 13.185 81.085 13.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 80.680 13.505 81.000 ;
      LAYER met4 ;
        RECT 13.185 80.680 13.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 80.275 13.505 80.595 ;
      LAYER met4 ;
        RECT 13.185 80.275 13.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 79.870 13.505 80.190 ;
      LAYER met4 ;
        RECT 13.185 79.870 13.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 79.465 13.505 79.785 ;
      LAYER met4 ;
        RECT 13.185 79.465 13.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 79.060 13.505 79.380 ;
      LAYER met4 ;
        RECT 13.185 79.060 13.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 78.655 13.505 78.975 ;
      LAYER met4 ;
        RECT 13.185 78.655 13.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 78.250 13.505 78.570 ;
      LAYER met4 ;
        RECT 13.185 78.250 13.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 77.845 13.505 78.165 ;
      LAYER met4 ;
        RECT 13.185 77.845 13.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 77.440 13.505 77.760 ;
      LAYER met4 ;
        RECT 13.185 77.440 13.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 77.035 13.505 77.355 ;
      LAYER met4 ;
        RECT 13.185 77.035 13.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 76.630 13.505 76.950 ;
      LAYER met4 ;
        RECT 13.185 76.630 13.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 76.225 13.505 76.545 ;
      LAYER met4 ;
        RECT 13.185 76.225 13.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 75.820 13.505 76.140 ;
      LAYER met4 ;
        RECT 13.185 75.820 13.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 75.415 13.505 75.735 ;
      LAYER met4 ;
        RECT 13.185 75.415 13.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 75.010 13.505 75.330 ;
      LAYER met4 ;
        RECT 13.185 75.010 13.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 74.605 13.505 74.925 ;
      LAYER met4 ;
        RECT 13.185 74.605 13.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 74.200 13.505 74.520 ;
      LAYER met4 ;
        RECT 13.185 74.200 13.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 73.795 13.505 74.115 ;
      LAYER met4 ;
        RECT 13.185 73.795 13.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 73.390 13.505 73.710 ;
      LAYER met4 ;
        RECT 13.185 73.390 13.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 72.985 13.505 73.305 ;
      LAYER met4 ;
        RECT 13.185 72.985 13.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 72.575 13.505 72.895 ;
      LAYER met4 ;
        RECT 13.185 72.575 13.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 72.165 13.505 72.485 ;
      LAYER met4 ;
        RECT 13.185 72.165 13.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 71.755 13.505 72.075 ;
      LAYER met4 ;
        RECT 13.185 71.755 13.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 71.345 13.505 71.665 ;
      LAYER met4 ;
        RECT 13.185 71.345 13.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 70.935 13.505 71.255 ;
      LAYER met4 ;
        RECT 13.185 70.935 13.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 70.525 13.505 70.845 ;
      LAYER met4 ;
        RECT 13.185 70.525 13.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 70.115 13.505 70.435 ;
      LAYER met4 ;
        RECT 13.185 70.115 13.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 69.705 13.505 70.025 ;
      LAYER met4 ;
        RECT 13.185 69.705 13.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 69.295 13.505 69.615 ;
      LAYER met4 ;
        RECT 13.185 69.295 13.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 68.885 13.505 69.205 ;
      LAYER met4 ;
        RECT 13.185 68.885 13.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 68.475 13.505 68.795 ;
      LAYER met4 ;
        RECT 13.185 68.475 13.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.185 68.065 13.505 68.385 ;
      LAYER met4 ;
        RECT 13.185 68.065 13.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 22.160 13.445 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 21.730 13.445 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 21.300 13.445 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 20.870 13.445 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 20.440 13.445 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 20.010 13.445 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 19.580 13.445 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 19.150 13.445 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 18.720 13.445 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 18.290 13.445 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.245 17.860 13.445 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 92.635 13.290 92.955 ;
      LAYER met4 ;
        RECT 12.970 92.635 13.290 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 92.225 13.290 92.545 ;
      LAYER met4 ;
        RECT 12.970 92.225 13.290 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 91.815 13.290 92.135 ;
      LAYER met4 ;
        RECT 12.970 91.815 13.290 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 91.405 13.290 91.725 ;
      LAYER met4 ;
        RECT 12.970 91.405 13.290 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 90.995 13.290 91.315 ;
      LAYER met4 ;
        RECT 12.970 90.995 13.290 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 90.585 13.290 90.905 ;
      LAYER met4 ;
        RECT 12.970 90.585 13.290 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 90.175 13.290 90.495 ;
      LAYER met4 ;
        RECT 12.970 90.175 13.290 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 89.765 13.290 90.085 ;
      LAYER met4 ;
        RECT 12.970 89.765 13.290 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 89.355 13.290 89.675 ;
      LAYER met4 ;
        RECT 12.970 89.355 13.290 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 88.945 13.290 89.265 ;
      LAYER met4 ;
        RECT 12.970 88.945 13.290 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 88.535 13.290 88.855 ;
      LAYER met4 ;
        RECT 12.970 88.535 13.290 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 88.125 13.290 88.445 ;
      LAYER met4 ;
        RECT 12.970 88.125 13.290 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 87.715 13.290 88.035 ;
      LAYER met4 ;
        RECT 12.970 87.715 13.290 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 87.305 13.290 87.625 ;
      LAYER met4 ;
        RECT 12.970 87.305 13.290 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 86.895 13.290 87.215 ;
      LAYER met4 ;
        RECT 12.970 86.895 13.290 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 86.485 13.290 86.805 ;
      LAYER met4 ;
        RECT 12.970 86.485 13.290 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 86.075 13.290 86.395 ;
      LAYER met4 ;
        RECT 12.970 86.075 13.290 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 85.665 13.290 85.985 ;
      LAYER met4 ;
        RECT 12.970 85.665 13.290 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 85.255 13.290 85.575 ;
      LAYER met4 ;
        RECT 12.970 85.255 13.290 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 84.845 13.290 85.165 ;
      LAYER met4 ;
        RECT 12.970 84.845 13.290 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 84.435 13.290 84.755 ;
      LAYER met4 ;
        RECT 12.970 84.435 13.290 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 84.025 13.290 84.345 ;
      LAYER met4 ;
        RECT 12.970 84.025 13.290 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 83.615 13.290 83.935 ;
      LAYER met4 ;
        RECT 12.970 83.615 13.290 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 83.205 13.290 83.525 ;
      LAYER met4 ;
        RECT 12.970 83.205 13.290 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.970 82.795 13.290 83.115 ;
      LAYER met4 ;
        RECT 12.970 82.795 13.290 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 82.300 13.105 82.620 ;
      LAYER met4 ;
        RECT 12.785 82.300 13.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 81.895 13.105 82.215 ;
      LAYER met4 ;
        RECT 12.785 81.895 13.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 81.490 13.105 81.810 ;
      LAYER met4 ;
        RECT 12.785 81.490 13.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 81.085 13.105 81.405 ;
      LAYER met4 ;
        RECT 12.785 81.085 13.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 80.680 13.105 81.000 ;
      LAYER met4 ;
        RECT 12.785 80.680 13.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 80.275 13.105 80.595 ;
      LAYER met4 ;
        RECT 12.785 80.275 13.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 79.870 13.105 80.190 ;
      LAYER met4 ;
        RECT 12.785 79.870 13.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 79.465 13.105 79.785 ;
      LAYER met4 ;
        RECT 12.785 79.465 13.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 79.060 13.105 79.380 ;
      LAYER met4 ;
        RECT 12.785 79.060 13.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 78.655 13.105 78.975 ;
      LAYER met4 ;
        RECT 12.785 78.655 13.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 78.250 13.105 78.570 ;
      LAYER met4 ;
        RECT 12.785 78.250 13.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 77.845 13.105 78.165 ;
      LAYER met4 ;
        RECT 12.785 77.845 13.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 77.440 13.105 77.760 ;
      LAYER met4 ;
        RECT 12.785 77.440 13.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 77.035 13.105 77.355 ;
      LAYER met4 ;
        RECT 12.785 77.035 13.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 76.630 13.105 76.950 ;
      LAYER met4 ;
        RECT 12.785 76.630 13.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 76.225 13.105 76.545 ;
      LAYER met4 ;
        RECT 12.785 76.225 13.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 75.820 13.105 76.140 ;
      LAYER met4 ;
        RECT 12.785 75.820 13.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 75.415 13.105 75.735 ;
      LAYER met4 ;
        RECT 12.785 75.415 13.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 75.010 13.105 75.330 ;
      LAYER met4 ;
        RECT 12.785 75.010 13.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 74.605 13.105 74.925 ;
      LAYER met4 ;
        RECT 12.785 74.605 13.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 74.200 13.105 74.520 ;
      LAYER met4 ;
        RECT 12.785 74.200 13.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 73.795 13.105 74.115 ;
      LAYER met4 ;
        RECT 12.785 73.795 13.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 73.390 13.105 73.710 ;
      LAYER met4 ;
        RECT 12.785 73.390 13.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 72.985 13.105 73.305 ;
      LAYER met4 ;
        RECT 12.785 72.985 13.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 72.575 13.105 72.895 ;
      LAYER met4 ;
        RECT 12.785 72.575 13.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 72.165 13.105 72.485 ;
      LAYER met4 ;
        RECT 12.785 72.165 13.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 71.755 13.105 72.075 ;
      LAYER met4 ;
        RECT 12.785 71.755 13.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 71.345 13.105 71.665 ;
      LAYER met4 ;
        RECT 12.785 71.345 13.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 70.935 13.105 71.255 ;
      LAYER met4 ;
        RECT 12.785 70.935 13.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 70.525 13.105 70.845 ;
      LAYER met4 ;
        RECT 12.785 70.525 13.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 70.115 13.105 70.435 ;
      LAYER met4 ;
        RECT 12.785 70.115 13.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 69.705 13.105 70.025 ;
      LAYER met4 ;
        RECT 12.785 69.705 13.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 69.295 13.105 69.615 ;
      LAYER met4 ;
        RECT 12.785 69.295 13.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 68.885 13.105 69.205 ;
      LAYER met4 ;
        RECT 12.785 68.885 13.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 68.475 13.105 68.795 ;
      LAYER met4 ;
        RECT 12.785 68.475 13.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.785 68.065 13.105 68.385 ;
      LAYER met4 ;
        RECT 12.785 68.065 13.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 22.160 13.040 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 21.730 13.040 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 21.300 13.040 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 20.870 13.040 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 20.440 13.040 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 20.010 13.040 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 19.580 13.040 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 19.150 13.040 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 18.720 13.040 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 18.290 13.040 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.840 17.860 13.040 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 92.635 12.885 92.955 ;
      LAYER met4 ;
        RECT 12.565 92.635 12.885 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 92.225 12.885 92.545 ;
      LAYER met4 ;
        RECT 12.565 92.225 12.885 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 91.815 12.885 92.135 ;
      LAYER met4 ;
        RECT 12.565 91.815 12.885 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 91.405 12.885 91.725 ;
      LAYER met4 ;
        RECT 12.565 91.405 12.885 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 90.995 12.885 91.315 ;
      LAYER met4 ;
        RECT 12.565 90.995 12.885 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 90.585 12.885 90.905 ;
      LAYER met4 ;
        RECT 12.565 90.585 12.885 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 90.175 12.885 90.495 ;
      LAYER met4 ;
        RECT 12.565 90.175 12.885 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 89.765 12.885 90.085 ;
      LAYER met4 ;
        RECT 12.565 89.765 12.885 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 89.355 12.885 89.675 ;
      LAYER met4 ;
        RECT 12.565 89.355 12.885 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 88.945 12.885 89.265 ;
      LAYER met4 ;
        RECT 12.565 88.945 12.885 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 88.535 12.885 88.855 ;
      LAYER met4 ;
        RECT 12.565 88.535 12.885 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 88.125 12.885 88.445 ;
      LAYER met4 ;
        RECT 12.565 88.125 12.885 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 87.715 12.885 88.035 ;
      LAYER met4 ;
        RECT 12.565 87.715 12.885 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 87.305 12.885 87.625 ;
      LAYER met4 ;
        RECT 12.565 87.305 12.885 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 86.895 12.885 87.215 ;
      LAYER met4 ;
        RECT 12.565 86.895 12.885 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 86.485 12.885 86.805 ;
      LAYER met4 ;
        RECT 12.565 86.485 12.885 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 86.075 12.885 86.395 ;
      LAYER met4 ;
        RECT 12.565 86.075 12.885 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 85.665 12.885 85.985 ;
      LAYER met4 ;
        RECT 12.565 85.665 12.885 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 85.255 12.885 85.575 ;
      LAYER met4 ;
        RECT 12.565 85.255 12.885 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 84.845 12.885 85.165 ;
      LAYER met4 ;
        RECT 12.565 84.845 12.885 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 84.435 12.885 84.755 ;
      LAYER met4 ;
        RECT 12.565 84.435 12.885 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 84.025 12.885 84.345 ;
      LAYER met4 ;
        RECT 12.565 84.025 12.885 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 83.615 12.885 83.935 ;
      LAYER met4 ;
        RECT 12.565 83.615 12.885 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 83.205 12.885 83.525 ;
      LAYER met4 ;
        RECT 12.565 83.205 12.885 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.565 82.795 12.885 83.115 ;
      LAYER met4 ;
        RECT 12.565 82.795 12.885 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 82.300 12.705 82.620 ;
      LAYER met4 ;
        RECT 12.385 82.300 12.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 81.895 12.705 82.215 ;
      LAYER met4 ;
        RECT 12.385 81.895 12.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 81.490 12.705 81.810 ;
      LAYER met4 ;
        RECT 12.385 81.490 12.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 81.085 12.705 81.405 ;
      LAYER met4 ;
        RECT 12.385 81.085 12.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 80.680 12.705 81.000 ;
      LAYER met4 ;
        RECT 12.385 80.680 12.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 80.275 12.705 80.595 ;
      LAYER met4 ;
        RECT 12.385 80.275 12.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 79.870 12.705 80.190 ;
      LAYER met4 ;
        RECT 12.385 79.870 12.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 79.465 12.705 79.785 ;
      LAYER met4 ;
        RECT 12.385 79.465 12.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 79.060 12.705 79.380 ;
      LAYER met4 ;
        RECT 12.385 79.060 12.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 78.655 12.705 78.975 ;
      LAYER met4 ;
        RECT 12.385 78.655 12.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 78.250 12.705 78.570 ;
      LAYER met4 ;
        RECT 12.385 78.250 12.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 77.845 12.705 78.165 ;
      LAYER met4 ;
        RECT 12.385 77.845 12.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 77.440 12.705 77.760 ;
      LAYER met4 ;
        RECT 12.385 77.440 12.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 77.035 12.705 77.355 ;
      LAYER met4 ;
        RECT 12.385 77.035 12.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 76.630 12.705 76.950 ;
      LAYER met4 ;
        RECT 12.385 76.630 12.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 76.225 12.705 76.545 ;
      LAYER met4 ;
        RECT 12.385 76.225 12.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 75.820 12.705 76.140 ;
      LAYER met4 ;
        RECT 12.385 75.820 12.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 75.415 12.705 75.735 ;
      LAYER met4 ;
        RECT 12.385 75.415 12.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 75.010 12.705 75.330 ;
      LAYER met4 ;
        RECT 12.385 75.010 12.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 74.605 12.705 74.925 ;
      LAYER met4 ;
        RECT 12.385 74.605 12.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 74.200 12.705 74.520 ;
      LAYER met4 ;
        RECT 12.385 74.200 12.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 73.795 12.705 74.115 ;
      LAYER met4 ;
        RECT 12.385 73.795 12.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 73.390 12.705 73.710 ;
      LAYER met4 ;
        RECT 12.385 73.390 12.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 72.985 12.705 73.305 ;
      LAYER met4 ;
        RECT 12.385 72.985 12.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 72.575 12.705 72.895 ;
      LAYER met4 ;
        RECT 12.385 72.575 12.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 72.165 12.705 72.485 ;
      LAYER met4 ;
        RECT 12.385 72.165 12.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 71.755 12.705 72.075 ;
      LAYER met4 ;
        RECT 12.385 71.755 12.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 71.345 12.705 71.665 ;
      LAYER met4 ;
        RECT 12.385 71.345 12.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 70.935 12.705 71.255 ;
      LAYER met4 ;
        RECT 12.385 70.935 12.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 70.525 12.705 70.845 ;
      LAYER met4 ;
        RECT 12.385 70.525 12.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 70.115 12.705 70.435 ;
      LAYER met4 ;
        RECT 12.385 70.115 12.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 69.705 12.705 70.025 ;
      LAYER met4 ;
        RECT 12.385 69.705 12.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 69.295 12.705 69.615 ;
      LAYER met4 ;
        RECT 12.385 69.295 12.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 68.885 12.705 69.205 ;
      LAYER met4 ;
        RECT 12.385 68.885 12.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 68.475 12.705 68.795 ;
      LAYER met4 ;
        RECT 12.385 68.475 12.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.385 68.065 12.705 68.385 ;
      LAYER met4 ;
        RECT 12.385 68.065 12.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 22.160 12.635 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 21.730 12.635 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 21.300 12.635 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 20.870 12.635 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 20.440 12.635 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 20.010 12.635 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 19.580 12.635 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 19.150 12.635 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 18.720 12.635 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 18.290 12.635 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.435 17.860 12.635 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 92.635 12.475 92.955 ;
      LAYER met4 ;
        RECT 12.155 92.635 12.475 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 92.225 12.475 92.545 ;
      LAYER met4 ;
        RECT 12.155 92.225 12.475 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 91.815 12.475 92.135 ;
      LAYER met4 ;
        RECT 12.155 91.815 12.475 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 91.405 12.475 91.725 ;
      LAYER met4 ;
        RECT 12.155 91.405 12.475 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 90.995 12.475 91.315 ;
      LAYER met4 ;
        RECT 12.155 90.995 12.475 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 90.585 12.475 90.905 ;
      LAYER met4 ;
        RECT 12.155 90.585 12.475 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 90.175 12.475 90.495 ;
      LAYER met4 ;
        RECT 12.155 90.175 12.475 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 89.765 12.475 90.085 ;
      LAYER met4 ;
        RECT 12.155 89.765 12.475 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 89.355 12.475 89.675 ;
      LAYER met4 ;
        RECT 12.155 89.355 12.475 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 88.945 12.475 89.265 ;
      LAYER met4 ;
        RECT 12.155 88.945 12.475 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 88.535 12.475 88.855 ;
      LAYER met4 ;
        RECT 12.155 88.535 12.475 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 88.125 12.475 88.445 ;
      LAYER met4 ;
        RECT 12.155 88.125 12.475 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 87.715 12.475 88.035 ;
      LAYER met4 ;
        RECT 12.155 87.715 12.475 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 87.305 12.475 87.625 ;
      LAYER met4 ;
        RECT 12.155 87.305 12.475 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 86.895 12.475 87.215 ;
      LAYER met4 ;
        RECT 12.155 86.895 12.475 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 86.485 12.475 86.805 ;
      LAYER met4 ;
        RECT 12.155 86.485 12.475 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 86.075 12.475 86.395 ;
      LAYER met4 ;
        RECT 12.155 86.075 12.475 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 85.665 12.475 85.985 ;
      LAYER met4 ;
        RECT 12.155 85.665 12.475 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 85.255 12.475 85.575 ;
      LAYER met4 ;
        RECT 12.155 85.255 12.475 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 84.845 12.475 85.165 ;
      LAYER met4 ;
        RECT 12.155 84.845 12.475 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 84.435 12.475 84.755 ;
      LAYER met4 ;
        RECT 12.155 84.435 12.475 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 84.025 12.475 84.345 ;
      LAYER met4 ;
        RECT 12.155 84.025 12.475 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 83.615 12.475 83.935 ;
      LAYER met4 ;
        RECT 12.155 83.615 12.475 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 83.205 12.475 83.525 ;
      LAYER met4 ;
        RECT 12.155 83.205 12.475 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 82.795 12.475 83.115 ;
      LAYER met4 ;
        RECT 12.155 82.795 12.475 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 82.300 12.305 82.620 ;
      LAYER met4 ;
        RECT 11.985 82.300 12.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 81.895 12.305 82.215 ;
      LAYER met4 ;
        RECT 11.985 81.895 12.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 81.490 12.305 81.810 ;
      LAYER met4 ;
        RECT 11.985 81.490 12.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 81.085 12.305 81.405 ;
      LAYER met4 ;
        RECT 11.985 81.085 12.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 80.680 12.305 81.000 ;
      LAYER met4 ;
        RECT 11.985 80.680 12.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 80.275 12.305 80.595 ;
      LAYER met4 ;
        RECT 11.985 80.275 12.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 79.870 12.305 80.190 ;
      LAYER met4 ;
        RECT 11.985 79.870 12.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 79.465 12.305 79.785 ;
      LAYER met4 ;
        RECT 11.985 79.465 12.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 79.060 12.305 79.380 ;
      LAYER met4 ;
        RECT 11.985 79.060 12.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 78.655 12.305 78.975 ;
      LAYER met4 ;
        RECT 11.985 78.655 12.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 78.250 12.305 78.570 ;
      LAYER met4 ;
        RECT 11.985 78.250 12.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 77.845 12.305 78.165 ;
      LAYER met4 ;
        RECT 11.985 77.845 12.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 77.440 12.305 77.760 ;
      LAYER met4 ;
        RECT 11.985 77.440 12.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 77.035 12.305 77.355 ;
      LAYER met4 ;
        RECT 11.985 77.035 12.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 76.630 12.305 76.950 ;
      LAYER met4 ;
        RECT 11.985 76.630 12.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 76.225 12.305 76.545 ;
      LAYER met4 ;
        RECT 11.985 76.225 12.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 75.820 12.305 76.140 ;
      LAYER met4 ;
        RECT 11.985 75.820 12.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 75.415 12.305 75.735 ;
      LAYER met4 ;
        RECT 11.985 75.415 12.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 75.010 12.305 75.330 ;
      LAYER met4 ;
        RECT 11.985 75.010 12.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 74.605 12.305 74.925 ;
      LAYER met4 ;
        RECT 11.985 74.605 12.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 74.200 12.305 74.520 ;
      LAYER met4 ;
        RECT 11.985 74.200 12.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 73.795 12.305 74.115 ;
      LAYER met4 ;
        RECT 11.985 73.795 12.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 73.390 12.305 73.710 ;
      LAYER met4 ;
        RECT 11.985 73.390 12.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 72.985 12.305 73.305 ;
      LAYER met4 ;
        RECT 11.985 72.985 12.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 72.575 12.305 72.895 ;
      LAYER met4 ;
        RECT 11.985 72.575 12.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 72.165 12.305 72.485 ;
      LAYER met4 ;
        RECT 11.985 72.165 12.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 71.755 12.305 72.075 ;
      LAYER met4 ;
        RECT 11.985 71.755 12.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 71.345 12.305 71.665 ;
      LAYER met4 ;
        RECT 11.985 71.345 12.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 70.935 12.305 71.255 ;
      LAYER met4 ;
        RECT 11.985 70.935 12.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 70.525 12.305 70.845 ;
      LAYER met4 ;
        RECT 11.985 70.525 12.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 70.115 12.305 70.435 ;
      LAYER met4 ;
        RECT 11.985 70.115 12.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 69.705 12.305 70.025 ;
      LAYER met4 ;
        RECT 11.985 69.705 12.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 69.295 12.305 69.615 ;
      LAYER met4 ;
        RECT 11.985 69.295 12.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 68.885 12.305 69.205 ;
      LAYER met4 ;
        RECT 11.985 68.885 12.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 68.475 12.305 68.795 ;
      LAYER met4 ;
        RECT 11.985 68.475 12.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.985 68.065 12.305 68.385 ;
      LAYER met4 ;
        RECT 11.985 68.065 12.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 22.160 12.230 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 21.730 12.230 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 21.300 12.230 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 20.870 12.230 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 20.440 12.230 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 20.010 12.230 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 19.580 12.230 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 19.150 12.230 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 18.720 12.230 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 18.290 12.230 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.030 17.860 12.230 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 92.635 12.065 92.955 ;
      LAYER met4 ;
        RECT 11.745 92.635 12.065 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 92.225 12.065 92.545 ;
      LAYER met4 ;
        RECT 11.745 92.225 12.065 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 91.815 12.065 92.135 ;
      LAYER met4 ;
        RECT 11.745 91.815 12.065 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 91.405 12.065 91.725 ;
      LAYER met4 ;
        RECT 11.745 91.405 12.065 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 90.995 12.065 91.315 ;
      LAYER met4 ;
        RECT 11.745 90.995 12.065 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 90.585 12.065 90.905 ;
      LAYER met4 ;
        RECT 11.745 90.585 12.065 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 90.175 12.065 90.495 ;
      LAYER met4 ;
        RECT 11.745 90.175 12.065 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 89.765 12.065 90.085 ;
      LAYER met4 ;
        RECT 11.745 89.765 12.065 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 89.355 12.065 89.675 ;
      LAYER met4 ;
        RECT 11.745 89.355 12.065 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 88.945 12.065 89.265 ;
      LAYER met4 ;
        RECT 11.745 88.945 12.065 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 88.535 12.065 88.855 ;
      LAYER met4 ;
        RECT 11.745 88.535 12.065 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 88.125 12.065 88.445 ;
      LAYER met4 ;
        RECT 11.745 88.125 12.065 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 87.715 12.065 88.035 ;
      LAYER met4 ;
        RECT 11.745 87.715 12.065 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 87.305 12.065 87.625 ;
      LAYER met4 ;
        RECT 11.745 87.305 12.065 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 86.895 12.065 87.215 ;
      LAYER met4 ;
        RECT 11.745 86.895 12.065 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 86.485 12.065 86.805 ;
      LAYER met4 ;
        RECT 11.745 86.485 12.065 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 86.075 12.065 86.395 ;
      LAYER met4 ;
        RECT 11.745 86.075 12.065 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 85.665 12.065 85.985 ;
      LAYER met4 ;
        RECT 11.745 85.665 12.065 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 85.255 12.065 85.575 ;
      LAYER met4 ;
        RECT 11.745 85.255 12.065 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 84.845 12.065 85.165 ;
      LAYER met4 ;
        RECT 11.745 84.845 12.065 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 84.435 12.065 84.755 ;
      LAYER met4 ;
        RECT 11.745 84.435 12.065 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 84.025 12.065 84.345 ;
      LAYER met4 ;
        RECT 11.745 84.025 12.065 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 83.615 12.065 83.935 ;
      LAYER met4 ;
        RECT 11.745 83.615 12.065 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 83.205 12.065 83.525 ;
      LAYER met4 ;
        RECT 11.745 83.205 12.065 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.745 82.795 12.065 83.115 ;
      LAYER met4 ;
        RECT 11.745 82.795 12.065 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 82.300 11.905 82.620 ;
      LAYER met4 ;
        RECT 11.585 82.300 11.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 81.895 11.905 82.215 ;
      LAYER met4 ;
        RECT 11.585 81.895 11.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 81.490 11.905 81.810 ;
      LAYER met4 ;
        RECT 11.585 81.490 11.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 81.085 11.905 81.405 ;
      LAYER met4 ;
        RECT 11.585 81.085 11.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 80.680 11.905 81.000 ;
      LAYER met4 ;
        RECT 11.585 80.680 11.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 80.275 11.905 80.595 ;
      LAYER met4 ;
        RECT 11.585 80.275 11.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 79.870 11.905 80.190 ;
      LAYER met4 ;
        RECT 11.585 79.870 11.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 79.465 11.905 79.785 ;
      LAYER met4 ;
        RECT 11.585 79.465 11.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 79.060 11.905 79.380 ;
      LAYER met4 ;
        RECT 11.585 79.060 11.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 78.655 11.905 78.975 ;
      LAYER met4 ;
        RECT 11.585 78.655 11.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 78.250 11.905 78.570 ;
      LAYER met4 ;
        RECT 11.585 78.250 11.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 77.845 11.905 78.165 ;
      LAYER met4 ;
        RECT 11.585 77.845 11.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 77.440 11.905 77.760 ;
      LAYER met4 ;
        RECT 11.585 77.440 11.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 77.035 11.905 77.355 ;
      LAYER met4 ;
        RECT 11.585 77.035 11.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 76.630 11.905 76.950 ;
      LAYER met4 ;
        RECT 11.585 76.630 11.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 76.225 11.905 76.545 ;
      LAYER met4 ;
        RECT 11.585 76.225 11.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 75.820 11.905 76.140 ;
      LAYER met4 ;
        RECT 11.585 75.820 11.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 75.415 11.905 75.735 ;
      LAYER met4 ;
        RECT 11.585 75.415 11.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 75.010 11.905 75.330 ;
      LAYER met4 ;
        RECT 11.585 75.010 11.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 74.605 11.905 74.925 ;
      LAYER met4 ;
        RECT 11.585 74.605 11.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 74.200 11.905 74.520 ;
      LAYER met4 ;
        RECT 11.585 74.200 11.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 73.795 11.905 74.115 ;
      LAYER met4 ;
        RECT 11.585 73.795 11.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 73.390 11.905 73.710 ;
      LAYER met4 ;
        RECT 11.585 73.390 11.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 72.985 11.905 73.305 ;
      LAYER met4 ;
        RECT 11.585 72.985 11.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 72.575 11.905 72.895 ;
      LAYER met4 ;
        RECT 11.585 72.575 11.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 72.165 11.905 72.485 ;
      LAYER met4 ;
        RECT 11.585 72.165 11.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 71.755 11.905 72.075 ;
      LAYER met4 ;
        RECT 11.585 71.755 11.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 71.345 11.905 71.665 ;
      LAYER met4 ;
        RECT 11.585 71.345 11.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 70.935 11.905 71.255 ;
      LAYER met4 ;
        RECT 11.585 70.935 11.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 70.525 11.905 70.845 ;
      LAYER met4 ;
        RECT 11.585 70.525 11.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 70.115 11.905 70.435 ;
      LAYER met4 ;
        RECT 11.585 70.115 11.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 69.705 11.905 70.025 ;
      LAYER met4 ;
        RECT 11.585 69.705 11.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 69.295 11.905 69.615 ;
      LAYER met4 ;
        RECT 11.585 69.295 11.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 68.885 11.905 69.205 ;
      LAYER met4 ;
        RECT 11.585 68.885 11.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 68.475 11.905 68.795 ;
      LAYER met4 ;
        RECT 11.585 68.475 11.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.585 68.065 11.905 68.385 ;
      LAYER met4 ;
        RECT 11.585 68.065 11.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 22.160 11.825 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 21.730 11.825 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 21.300 11.825 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 20.870 11.825 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 20.440 11.825 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 20.010 11.825 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 19.580 11.825 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 19.150 11.825 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 18.720 11.825 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 18.290 11.825 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.625 17.860 11.825 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 92.635 11.655 92.955 ;
      LAYER met4 ;
        RECT 11.335 92.635 11.655 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 92.225 11.655 92.545 ;
      LAYER met4 ;
        RECT 11.335 92.225 11.655 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 91.815 11.655 92.135 ;
      LAYER met4 ;
        RECT 11.335 91.815 11.655 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 91.405 11.655 91.725 ;
      LAYER met4 ;
        RECT 11.335 91.405 11.655 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 90.995 11.655 91.315 ;
      LAYER met4 ;
        RECT 11.335 90.995 11.655 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 90.585 11.655 90.905 ;
      LAYER met4 ;
        RECT 11.335 90.585 11.655 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 90.175 11.655 90.495 ;
      LAYER met4 ;
        RECT 11.335 90.175 11.655 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 89.765 11.655 90.085 ;
      LAYER met4 ;
        RECT 11.335 89.765 11.655 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 89.355 11.655 89.675 ;
      LAYER met4 ;
        RECT 11.335 89.355 11.655 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 88.945 11.655 89.265 ;
      LAYER met4 ;
        RECT 11.335 88.945 11.655 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 88.535 11.655 88.855 ;
      LAYER met4 ;
        RECT 11.335 88.535 11.655 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 88.125 11.655 88.445 ;
      LAYER met4 ;
        RECT 11.335 88.125 11.655 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 87.715 11.655 88.035 ;
      LAYER met4 ;
        RECT 11.335 87.715 11.655 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 87.305 11.655 87.625 ;
      LAYER met4 ;
        RECT 11.335 87.305 11.655 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 86.895 11.655 87.215 ;
      LAYER met4 ;
        RECT 11.335 86.895 11.655 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 86.485 11.655 86.805 ;
      LAYER met4 ;
        RECT 11.335 86.485 11.655 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 86.075 11.655 86.395 ;
      LAYER met4 ;
        RECT 11.335 86.075 11.655 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 85.665 11.655 85.985 ;
      LAYER met4 ;
        RECT 11.335 85.665 11.655 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 85.255 11.655 85.575 ;
      LAYER met4 ;
        RECT 11.335 85.255 11.655 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 84.845 11.655 85.165 ;
      LAYER met4 ;
        RECT 11.335 84.845 11.655 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 84.435 11.655 84.755 ;
      LAYER met4 ;
        RECT 11.335 84.435 11.655 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 84.025 11.655 84.345 ;
      LAYER met4 ;
        RECT 11.335 84.025 11.655 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 83.615 11.655 83.935 ;
      LAYER met4 ;
        RECT 11.335 83.615 11.655 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 83.205 11.655 83.525 ;
      LAYER met4 ;
        RECT 11.335 83.205 11.655 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.335 82.795 11.655 83.115 ;
      LAYER met4 ;
        RECT 11.335 82.795 11.655 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 82.300 11.505 82.620 ;
      LAYER met4 ;
        RECT 11.185 82.300 11.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 81.895 11.505 82.215 ;
      LAYER met4 ;
        RECT 11.185 81.895 11.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 81.490 11.505 81.810 ;
      LAYER met4 ;
        RECT 11.185 81.490 11.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 81.085 11.505 81.405 ;
      LAYER met4 ;
        RECT 11.185 81.085 11.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 80.680 11.505 81.000 ;
      LAYER met4 ;
        RECT 11.185 80.680 11.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 80.275 11.505 80.595 ;
      LAYER met4 ;
        RECT 11.185 80.275 11.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 79.870 11.505 80.190 ;
      LAYER met4 ;
        RECT 11.185 79.870 11.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 79.465 11.505 79.785 ;
      LAYER met4 ;
        RECT 11.185 79.465 11.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 79.060 11.505 79.380 ;
      LAYER met4 ;
        RECT 11.185 79.060 11.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 78.655 11.505 78.975 ;
      LAYER met4 ;
        RECT 11.185 78.655 11.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 78.250 11.505 78.570 ;
      LAYER met4 ;
        RECT 11.185 78.250 11.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 77.845 11.505 78.165 ;
      LAYER met4 ;
        RECT 11.185 77.845 11.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 77.440 11.505 77.760 ;
      LAYER met4 ;
        RECT 11.185 77.440 11.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 77.035 11.505 77.355 ;
      LAYER met4 ;
        RECT 11.185 77.035 11.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 76.630 11.505 76.950 ;
      LAYER met4 ;
        RECT 11.185 76.630 11.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 76.225 11.505 76.545 ;
      LAYER met4 ;
        RECT 11.185 76.225 11.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 75.820 11.505 76.140 ;
      LAYER met4 ;
        RECT 11.185 75.820 11.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 75.415 11.505 75.735 ;
      LAYER met4 ;
        RECT 11.185 75.415 11.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 75.010 11.505 75.330 ;
      LAYER met4 ;
        RECT 11.185 75.010 11.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 74.605 11.505 74.925 ;
      LAYER met4 ;
        RECT 11.185 74.605 11.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 74.200 11.505 74.520 ;
      LAYER met4 ;
        RECT 11.185 74.200 11.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 73.795 11.505 74.115 ;
      LAYER met4 ;
        RECT 11.185 73.795 11.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 73.390 11.505 73.710 ;
      LAYER met4 ;
        RECT 11.185 73.390 11.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 72.985 11.505 73.305 ;
      LAYER met4 ;
        RECT 11.185 72.985 11.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 72.575 11.505 72.895 ;
      LAYER met4 ;
        RECT 11.185 72.575 11.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 72.165 11.505 72.485 ;
      LAYER met4 ;
        RECT 11.185 72.165 11.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 71.755 11.505 72.075 ;
      LAYER met4 ;
        RECT 11.185 71.755 11.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 71.345 11.505 71.665 ;
      LAYER met4 ;
        RECT 11.185 71.345 11.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 70.935 11.505 71.255 ;
      LAYER met4 ;
        RECT 11.185 70.935 11.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 70.525 11.505 70.845 ;
      LAYER met4 ;
        RECT 11.185 70.525 11.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 70.115 11.505 70.435 ;
      LAYER met4 ;
        RECT 11.185 70.115 11.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 69.705 11.505 70.025 ;
      LAYER met4 ;
        RECT 11.185 69.705 11.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 69.295 11.505 69.615 ;
      LAYER met4 ;
        RECT 11.185 69.295 11.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 68.885 11.505 69.205 ;
      LAYER met4 ;
        RECT 11.185 68.885 11.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 68.475 11.505 68.795 ;
      LAYER met4 ;
        RECT 11.185 68.475 11.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 68.065 11.505 68.385 ;
      LAYER met4 ;
        RECT 11.185 68.065 11.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 22.160 11.420 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 21.730 11.420 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 21.300 11.420 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 20.870 11.420 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 20.440 11.420 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 20.010 11.420 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 19.580 11.420 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 19.150 11.420 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 18.720 11.420 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 18.290 11.420 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.220 17.860 11.420 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 92.635 11.245 92.955 ;
      LAYER met4 ;
        RECT 10.925 92.635 11.245 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 92.225 11.245 92.545 ;
      LAYER met4 ;
        RECT 10.925 92.225 11.245 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 91.815 11.245 92.135 ;
      LAYER met4 ;
        RECT 10.925 91.815 11.245 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 91.405 11.245 91.725 ;
      LAYER met4 ;
        RECT 10.925 91.405 11.245 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 90.995 11.245 91.315 ;
      LAYER met4 ;
        RECT 10.925 90.995 11.245 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 90.585 11.245 90.905 ;
      LAYER met4 ;
        RECT 10.925 90.585 11.245 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 90.175 11.245 90.495 ;
      LAYER met4 ;
        RECT 10.925 90.175 11.245 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 89.765 11.245 90.085 ;
      LAYER met4 ;
        RECT 10.925 89.765 11.245 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 89.355 11.245 89.675 ;
      LAYER met4 ;
        RECT 10.925 89.355 11.245 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 88.945 11.245 89.265 ;
      LAYER met4 ;
        RECT 10.925 88.945 11.245 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 88.535 11.245 88.855 ;
      LAYER met4 ;
        RECT 10.925 88.535 11.245 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 88.125 11.245 88.445 ;
      LAYER met4 ;
        RECT 10.925 88.125 11.245 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 87.715 11.245 88.035 ;
      LAYER met4 ;
        RECT 10.925 87.715 11.245 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 87.305 11.245 87.625 ;
      LAYER met4 ;
        RECT 10.925 87.305 11.245 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 86.895 11.245 87.215 ;
      LAYER met4 ;
        RECT 10.925 86.895 11.245 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 86.485 11.245 86.805 ;
      LAYER met4 ;
        RECT 10.925 86.485 11.245 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 86.075 11.245 86.395 ;
      LAYER met4 ;
        RECT 10.925 86.075 11.245 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 85.665 11.245 85.985 ;
      LAYER met4 ;
        RECT 10.925 85.665 11.245 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 85.255 11.245 85.575 ;
      LAYER met4 ;
        RECT 10.925 85.255 11.245 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 84.845 11.245 85.165 ;
      LAYER met4 ;
        RECT 10.925 84.845 11.245 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 84.435 11.245 84.755 ;
      LAYER met4 ;
        RECT 10.925 84.435 11.245 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 84.025 11.245 84.345 ;
      LAYER met4 ;
        RECT 10.925 84.025 11.245 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 83.615 11.245 83.935 ;
      LAYER met4 ;
        RECT 10.925 83.615 11.245 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 83.205 11.245 83.525 ;
      LAYER met4 ;
        RECT 10.925 83.205 11.245 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.925 82.795 11.245 83.115 ;
      LAYER met4 ;
        RECT 10.925 82.795 11.245 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 82.300 11.105 82.620 ;
      LAYER met4 ;
        RECT 10.785 82.300 11.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 81.895 11.105 82.215 ;
      LAYER met4 ;
        RECT 10.785 81.895 11.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 81.490 11.105 81.810 ;
      LAYER met4 ;
        RECT 10.785 81.490 11.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 81.085 11.105 81.405 ;
      LAYER met4 ;
        RECT 10.785 81.085 11.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 80.680 11.105 81.000 ;
      LAYER met4 ;
        RECT 10.785 80.680 11.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 80.275 11.105 80.595 ;
      LAYER met4 ;
        RECT 10.785 80.275 11.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 79.870 11.105 80.190 ;
      LAYER met4 ;
        RECT 10.785 79.870 11.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 79.465 11.105 79.785 ;
      LAYER met4 ;
        RECT 10.785 79.465 11.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 79.060 11.105 79.380 ;
      LAYER met4 ;
        RECT 10.785 79.060 11.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 78.655 11.105 78.975 ;
      LAYER met4 ;
        RECT 10.785 78.655 11.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 78.250 11.105 78.570 ;
      LAYER met4 ;
        RECT 10.785 78.250 11.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 77.845 11.105 78.165 ;
      LAYER met4 ;
        RECT 10.785 77.845 11.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 77.440 11.105 77.760 ;
      LAYER met4 ;
        RECT 10.785 77.440 11.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 77.035 11.105 77.355 ;
      LAYER met4 ;
        RECT 10.785 77.035 11.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 76.630 11.105 76.950 ;
      LAYER met4 ;
        RECT 10.785 76.630 11.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 76.225 11.105 76.545 ;
      LAYER met4 ;
        RECT 10.785 76.225 11.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 75.820 11.105 76.140 ;
      LAYER met4 ;
        RECT 10.785 75.820 11.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 75.415 11.105 75.735 ;
      LAYER met4 ;
        RECT 10.785 75.415 11.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 75.010 11.105 75.330 ;
      LAYER met4 ;
        RECT 10.785 75.010 11.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 74.605 11.105 74.925 ;
      LAYER met4 ;
        RECT 10.785 74.605 11.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 74.200 11.105 74.520 ;
      LAYER met4 ;
        RECT 10.785 74.200 11.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 73.795 11.105 74.115 ;
      LAYER met4 ;
        RECT 10.785 73.795 11.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 73.390 11.105 73.710 ;
      LAYER met4 ;
        RECT 10.785 73.390 11.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 72.985 11.105 73.305 ;
      LAYER met4 ;
        RECT 10.785 72.985 11.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 72.575 11.105 72.895 ;
      LAYER met4 ;
        RECT 10.785 72.575 11.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 72.165 11.105 72.485 ;
      LAYER met4 ;
        RECT 10.785 72.165 11.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 71.755 11.105 72.075 ;
      LAYER met4 ;
        RECT 10.785 71.755 11.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 71.345 11.105 71.665 ;
      LAYER met4 ;
        RECT 10.785 71.345 11.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 70.935 11.105 71.255 ;
      LAYER met4 ;
        RECT 10.785 70.935 11.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 70.525 11.105 70.845 ;
      LAYER met4 ;
        RECT 10.785 70.525 11.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 70.115 11.105 70.435 ;
      LAYER met4 ;
        RECT 10.785 70.115 11.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 69.705 11.105 70.025 ;
      LAYER met4 ;
        RECT 10.785 69.705 11.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 69.295 11.105 69.615 ;
      LAYER met4 ;
        RECT 10.785 69.295 11.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 68.885 11.105 69.205 ;
      LAYER met4 ;
        RECT 10.785 68.885 11.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 68.475 11.105 68.795 ;
      LAYER met4 ;
        RECT 10.785 68.475 11.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.785 68.065 11.105 68.385 ;
      LAYER met4 ;
        RECT 10.785 68.065 11.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 22.160 11.015 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 21.730 11.015 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 21.300 11.015 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 20.870 11.015 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 20.440 11.015 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 20.010 11.015 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 19.580 11.015 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 19.150 11.015 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 18.720 11.015 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 18.290 11.015 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.815 17.860 11.015 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 92.635 10.835 92.955 ;
      LAYER met4 ;
        RECT 10.515 92.635 10.835 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 92.225 10.835 92.545 ;
      LAYER met4 ;
        RECT 10.515 92.225 10.835 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 91.815 10.835 92.135 ;
      LAYER met4 ;
        RECT 10.515 91.815 10.835 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 91.405 10.835 91.725 ;
      LAYER met4 ;
        RECT 10.515 91.405 10.835 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 90.995 10.835 91.315 ;
      LAYER met4 ;
        RECT 10.515 90.995 10.835 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 90.585 10.835 90.905 ;
      LAYER met4 ;
        RECT 10.515 90.585 10.835 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 90.175 10.835 90.495 ;
      LAYER met4 ;
        RECT 10.515 90.175 10.835 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 89.765 10.835 90.085 ;
      LAYER met4 ;
        RECT 10.515 89.765 10.835 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 89.355 10.835 89.675 ;
      LAYER met4 ;
        RECT 10.515 89.355 10.835 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 88.945 10.835 89.265 ;
      LAYER met4 ;
        RECT 10.515 88.945 10.835 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 88.535 10.835 88.855 ;
      LAYER met4 ;
        RECT 10.515 88.535 10.835 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 88.125 10.835 88.445 ;
      LAYER met4 ;
        RECT 10.515 88.125 10.835 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 87.715 10.835 88.035 ;
      LAYER met4 ;
        RECT 10.515 87.715 10.835 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 87.305 10.835 87.625 ;
      LAYER met4 ;
        RECT 10.515 87.305 10.835 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 86.895 10.835 87.215 ;
      LAYER met4 ;
        RECT 10.515 86.895 10.835 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 86.485 10.835 86.805 ;
      LAYER met4 ;
        RECT 10.515 86.485 10.835 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 86.075 10.835 86.395 ;
      LAYER met4 ;
        RECT 10.515 86.075 10.835 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 85.665 10.835 85.985 ;
      LAYER met4 ;
        RECT 10.515 85.665 10.835 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 85.255 10.835 85.575 ;
      LAYER met4 ;
        RECT 10.515 85.255 10.835 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 84.845 10.835 85.165 ;
      LAYER met4 ;
        RECT 10.515 84.845 10.835 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 84.435 10.835 84.755 ;
      LAYER met4 ;
        RECT 10.515 84.435 10.835 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 84.025 10.835 84.345 ;
      LAYER met4 ;
        RECT 10.515 84.025 10.835 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 83.615 10.835 83.935 ;
      LAYER met4 ;
        RECT 10.515 83.615 10.835 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 83.205 10.835 83.525 ;
      LAYER met4 ;
        RECT 10.515 83.205 10.835 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.515 82.795 10.835 83.115 ;
      LAYER met4 ;
        RECT 10.515 82.795 10.835 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 82.300 10.705 82.620 ;
      LAYER met4 ;
        RECT 10.385 82.300 10.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 81.895 10.705 82.215 ;
      LAYER met4 ;
        RECT 10.385 81.895 10.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 81.490 10.705 81.810 ;
      LAYER met4 ;
        RECT 10.385 81.490 10.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 81.085 10.705 81.405 ;
      LAYER met4 ;
        RECT 10.385 81.085 10.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 80.680 10.705 81.000 ;
      LAYER met4 ;
        RECT 10.385 80.680 10.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 80.275 10.705 80.595 ;
      LAYER met4 ;
        RECT 10.385 80.275 10.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 79.870 10.705 80.190 ;
      LAYER met4 ;
        RECT 10.385 79.870 10.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 79.465 10.705 79.785 ;
      LAYER met4 ;
        RECT 10.385 79.465 10.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 79.060 10.705 79.380 ;
      LAYER met4 ;
        RECT 10.385 79.060 10.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 78.655 10.705 78.975 ;
      LAYER met4 ;
        RECT 10.385 78.655 10.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 78.250 10.705 78.570 ;
      LAYER met4 ;
        RECT 10.385 78.250 10.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 77.845 10.705 78.165 ;
      LAYER met4 ;
        RECT 10.385 77.845 10.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 77.440 10.705 77.760 ;
      LAYER met4 ;
        RECT 10.385 77.440 10.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 77.035 10.705 77.355 ;
      LAYER met4 ;
        RECT 10.385 77.035 10.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 76.630 10.705 76.950 ;
      LAYER met4 ;
        RECT 10.385 76.630 10.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 76.225 10.705 76.545 ;
      LAYER met4 ;
        RECT 10.385 76.225 10.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 75.820 10.705 76.140 ;
      LAYER met4 ;
        RECT 10.385 75.820 10.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 75.415 10.705 75.735 ;
      LAYER met4 ;
        RECT 10.385 75.415 10.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 75.010 10.705 75.330 ;
      LAYER met4 ;
        RECT 10.385 75.010 10.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 74.605 10.705 74.925 ;
      LAYER met4 ;
        RECT 10.385 74.605 10.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 74.200 10.705 74.520 ;
      LAYER met4 ;
        RECT 10.385 74.200 10.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 73.795 10.705 74.115 ;
      LAYER met4 ;
        RECT 10.385 73.795 10.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 73.390 10.705 73.710 ;
      LAYER met4 ;
        RECT 10.385 73.390 10.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 72.985 10.705 73.305 ;
      LAYER met4 ;
        RECT 10.385 72.985 10.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 72.575 10.705 72.895 ;
      LAYER met4 ;
        RECT 10.385 72.575 10.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 72.165 10.705 72.485 ;
      LAYER met4 ;
        RECT 10.385 72.165 10.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 71.755 10.705 72.075 ;
      LAYER met4 ;
        RECT 10.385 71.755 10.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 71.345 10.705 71.665 ;
      LAYER met4 ;
        RECT 10.385 71.345 10.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 70.935 10.705 71.255 ;
      LAYER met4 ;
        RECT 10.385 70.935 10.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 70.525 10.705 70.845 ;
      LAYER met4 ;
        RECT 10.385 70.525 10.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 70.115 10.705 70.435 ;
      LAYER met4 ;
        RECT 10.385 70.115 10.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 69.705 10.705 70.025 ;
      LAYER met4 ;
        RECT 10.385 69.705 10.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 69.295 10.705 69.615 ;
      LAYER met4 ;
        RECT 10.385 69.295 10.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 68.885 10.705 69.205 ;
      LAYER met4 ;
        RECT 10.385 68.885 10.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 68.475 10.705 68.795 ;
      LAYER met4 ;
        RECT 10.385 68.475 10.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.385 68.065 10.705 68.385 ;
      LAYER met4 ;
        RECT 10.385 68.065 10.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 22.160 10.610 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 21.730 10.610 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 21.300 10.610 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 20.870 10.610 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 20.440 10.610 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 20.010 10.610 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 19.580 10.610 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 19.150 10.610 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 18.720 10.610 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 18.290 10.610 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.410 17.860 10.610 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 92.635 10.425 92.955 ;
      LAYER met4 ;
        RECT 10.105 92.635 10.425 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 92.225 10.425 92.545 ;
      LAYER met4 ;
        RECT 10.105 92.225 10.425 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 91.815 10.425 92.135 ;
      LAYER met4 ;
        RECT 10.105 91.815 10.425 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 91.405 10.425 91.725 ;
      LAYER met4 ;
        RECT 10.105 91.405 10.425 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 90.995 10.425 91.315 ;
      LAYER met4 ;
        RECT 10.105 90.995 10.425 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 90.585 10.425 90.905 ;
      LAYER met4 ;
        RECT 10.105 90.585 10.425 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 90.175 10.425 90.495 ;
      LAYER met4 ;
        RECT 10.105 90.175 10.425 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 89.765 10.425 90.085 ;
      LAYER met4 ;
        RECT 10.105 89.765 10.425 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 89.355 10.425 89.675 ;
      LAYER met4 ;
        RECT 10.105 89.355 10.425 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 88.945 10.425 89.265 ;
      LAYER met4 ;
        RECT 10.105 88.945 10.425 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 88.535 10.425 88.855 ;
      LAYER met4 ;
        RECT 10.105 88.535 10.425 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 88.125 10.425 88.445 ;
      LAYER met4 ;
        RECT 10.105 88.125 10.425 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 87.715 10.425 88.035 ;
      LAYER met4 ;
        RECT 10.105 87.715 10.425 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 87.305 10.425 87.625 ;
      LAYER met4 ;
        RECT 10.105 87.305 10.425 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 86.895 10.425 87.215 ;
      LAYER met4 ;
        RECT 10.105 86.895 10.425 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 86.485 10.425 86.805 ;
      LAYER met4 ;
        RECT 10.105 86.485 10.425 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 86.075 10.425 86.395 ;
      LAYER met4 ;
        RECT 10.105 86.075 10.425 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 85.665 10.425 85.985 ;
      LAYER met4 ;
        RECT 10.105 85.665 10.425 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 85.255 10.425 85.575 ;
      LAYER met4 ;
        RECT 10.105 85.255 10.425 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 84.845 10.425 85.165 ;
      LAYER met4 ;
        RECT 10.105 84.845 10.425 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 84.435 10.425 84.755 ;
      LAYER met4 ;
        RECT 10.105 84.435 10.425 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 84.025 10.425 84.345 ;
      LAYER met4 ;
        RECT 10.105 84.025 10.425 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 83.615 10.425 83.935 ;
      LAYER met4 ;
        RECT 10.105 83.615 10.425 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 83.205 10.425 83.525 ;
      LAYER met4 ;
        RECT 10.105 83.205 10.425 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.105 82.795 10.425 83.115 ;
      LAYER met4 ;
        RECT 10.105 82.795 10.425 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 82.300 10.305 82.620 ;
      LAYER met4 ;
        RECT 9.985 82.300 10.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 81.895 10.305 82.215 ;
      LAYER met4 ;
        RECT 9.985 81.895 10.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 81.490 10.305 81.810 ;
      LAYER met4 ;
        RECT 9.985 81.490 10.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 81.085 10.305 81.405 ;
      LAYER met4 ;
        RECT 9.985 81.085 10.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 80.680 10.305 81.000 ;
      LAYER met4 ;
        RECT 9.985 80.680 10.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 80.275 10.305 80.595 ;
      LAYER met4 ;
        RECT 9.985 80.275 10.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 79.870 10.305 80.190 ;
      LAYER met4 ;
        RECT 9.985 79.870 10.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 79.465 10.305 79.785 ;
      LAYER met4 ;
        RECT 9.985 79.465 10.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 79.060 10.305 79.380 ;
      LAYER met4 ;
        RECT 9.985 79.060 10.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 78.655 10.305 78.975 ;
      LAYER met4 ;
        RECT 9.985 78.655 10.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 78.250 10.305 78.570 ;
      LAYER met4 ;
        RECT 9.985 78.250 10.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 77.845 10.305 78.165 ;
      LAYER met4 ;
        RECT 9.985 77.845 10.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 77.440 10.305 77.760 ;
      LAYER met4 ;
        RECT 9.985 77.440 10.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 77.035 10.305 77.355 ;
      LAYER met4 ;
        RECT 9.985 77.035 10.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 76.630 10.305 76.950 ;
      LAYER met4 ;
        RECT 9.985 76.630 10.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 76.225 10.305 76.545 ;
      LAYER met4 ;
        RECT 9.985 76.225 10.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 75.820 10.305 76.140 ;
      LAYER met4 ;
        RECT 9.985 75.820 10.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 75.415 10.305 75.735 ;
      LAYER met4 ;
        RECT 9.985 75.415 10.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 75.010 10.305 75.330 ;
      LAYER met4 ;
        RECT 9.985 75.010 10.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 74.605 10.305 74.925 ;
      LAYER met4 ;
        RECT 9.985 74.605 10.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 74.200 10.305 74.520 ;
      LAYER met4 ;
        RECT 9.985 74.200 10.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 73.795 10.305 74.115 ;
      LAYER met4 ;
        RECT 9.985 73.795 10.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 73.390 10.305 73.710 ;
      LAYER met4 ;
        RECT 9.985 73.390 10.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 72.985 10.305 73.305 ;
      LAYER met4 ;
        RECT 9.985 72.985 10.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 72.575 10.305 72.895 ;
      LAYER met4 ;
        RECT 9.985 72.575 10.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 72.165 10.305 72.485 ;
      LAYER met4 ;
        RECT 9.985 72.165 10.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 71.755 10.305 72.075 ;
      LAYER met4 ;
        RECT 9.985 71.755 10.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 71.345 10.305 71.665 ;
      LAYER met4 ;
        RECT 9.985 71.345 10.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 70.935 10.305 71.255 ;
      LAYER met4 ;
        RECT 9.985 70.935 10.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 70.525 10.305 70.845 ;
      LAYER met4 ;
        RECT 9.985 70.525 10.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 70.115 10.305 70.435 ;
      LAYER met4 ;
        RECT 9.985 70.115 10.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 69.705 10.305 70.025 ;
      LAYER met4 ;
        RECT 9.985 69.705 10.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 69.295 10.305 69.615 ;
      LAYER met4 ;
        RECT 9.985 69.295 10.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 68.885 10.305 69.205 ;
      LAYER met4 ;
        RECT 9.985 68.885 10.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 68.475 10.305 68.795 ;
      LAYER met4 ;
        RECT 9.985 68.475 10.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.985 68.065 10.305 68.385 ;
      LAYER met4 ;
        RECT 9.985 68.065 10.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 22.160 10.205 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 21.730 10.205 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 21.300 10.205 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 20.870 10.205 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 20.440 10.205 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 20.010 10.205 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 19.580 10.205 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 19.150 10.205 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 18.720 10.205 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 18.290 10.205 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.005 17.860 10.205 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 92.635 10.015 92.955 ;
      LAYER met4 ;
        RECT 9.695 92.635 10.015 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 92.225 10.015 92.545 ;
      LAYER met4 ;
        RECT 9.695 92.225 10.015 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 91.815 10.015 92.135 ;
      LAYER met4 ;
        RECT 9.695 91.815 10.015 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 91.405 10.015 91.725 ;
      LAYER met4 ;
        RECT 9.695 91.405 10.015 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 90.995 10.015 91.315 ;
      LAYER met4 ;
        RECT 9.695 90.995 10.015 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 90.585 10.015 90.905 ;
      LAYER met4 ;
        RECT 9.695 90.585 10.015 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 90.175 10.015 90.495 ;
      LAYER met4 ;
        RECT 9.695 90.175 10.015 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 89.765 10.015 90.085 ;
      LAYER met4 ;
        RECT 9.695 89.765 10.015 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 89.355 10.015 89.675 ;
      LAYER met4 ;
        RECT 9.695 89.355 10.015 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 88.945 10.015 89.265 ;
      LAYER met4 ;
        RECT 9.695 88.945 10.015 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 88.535 10.015 88.855 ;
      LAYER met4 ;
        RECT 9.695 88.535 10.015 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 88.125 10.015 88.445 ;
      LAYER met4 ;
        RECT 9.695 88.125 10.015 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 87.715 10.015 88.035 ;
      LAYER met4 ;
        RECT 9.695 87.715 10.015 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 87.305 10.015 87.625 ;
      LAYER met4 ;
        RECT 9.695 87.305 10.015 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 86.895 10.015 87.215 ;
      LAYER met4 ;
        RECT 9.695 86.895 10.015 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 86.485 10.015 86.805 ;
      LAYER met4 ;
        RECT 9.695 86.485 10.015 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 86.075 10.015 86.395 ;
      LAYER met4 ;
        RECT 9.695 86.075 10.015 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 85.665 10.015 85.985 ;
      LAYER met4 ;
        RECT 9.695 85.665 10.015 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 85.255 10.015 85.575 ;
      LAYER met4 ;
        RECT 9.695 85.255 10.015 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 84.845 10.015 85.165 ;
      LAYER met4 ;
        RECT 9.695 84.845 10.015 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 84.435 10.015 84.755 ;
      LAYER met4 ;
        RECT 9.695 84.435 10.015 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 84.025 10.015 84.345 ;
      LAYER met4 ;
        RECT 9.695 84.025 10.015 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 83.615 10.015 83.935 ;
      LAYER met4 ;
        RECT 9.695 83.615 10.015 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 83.205 10.015 83.525 ;
      LAYER met4 ;
        RECT 9.695 83.205 10.015 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.695 82.795 10.015 83.115 ;
      LAYER met4 ;
        RECT 9.695 82.795 10.015 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 82.300 9.905 82.620 ;
      LAYER met4 ;
        RECT 9.585 82.300 9.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 81.895 9.905 82.215 ;
      LAYER met4 ;
        RECT 9.585 81.895 9.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 81.490 9.905 81.810 ;
      LAYER met4 ;
        RECT 9.585 81.490 9.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 81.085 9.905 81.405 ;
      LAYER met4 ;
        RECT 9.585 81.085 9.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 80.680 9.905 81.000 ;
      LAYER met4 ;
        RECT 9.585 80.680 9.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 80.275 9.905 80.595 ;
      LAYER met4 ;
        RECT 9.585 80.275 9.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 79.870 9.905 80.190 ;
      LAYER met4 ;
        RECT 9.585 79.870 9.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 79.465 9.905 79.785 ;
      LAYER met4 ;
        RECT 9.585 79.465 9.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 79.060 9.905 79.380 ;
      LAYER met4 ;
        RECT 9.585 79.060 9.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 78.655 9.905 78.975 ;
      LAYER met4 ;
        RECT 9.585 78.655 9.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 78.250 9.905 78.570 ;
      LAYER met4 ;
        RECT 9.585 78.250 9.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 77.845 9.905 78.165 ;
      LAYER met4 ;
        RECT 9.585 77.845 9.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 77.440 9.905 77.760 ;
      LAYER met4 ;
        RECT 9.585 77.440 9.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 77.035 9.905 77.355 ;
      LAYER met4 ;
        RECT 9.585 77.035 9.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 76.630 9.905 76.950 ;
      LAYER met4 ;
        RECT 9.585 76.630 9.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 76.225 9.905 76.545 ;
      LAYER met4 ;
        RECT 9.585 76.225 9.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 75.820 9.905 76.140 ;
      LAYER met4 ;
        RECT 9.585 75.820 9.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 75.415 9.905 75.735 ;
      LAYER met4 ;
        RECT 9.585 75.415 9.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 75.010 9.905 75.330 ;
      LAYER met4 ;
        RECT 9.585 75.010 9.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 74.605 9.905 74.925 ;
      LAYER met4 ;
        RECT 9.585 74.605 9.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 74.200 9.905 74.520 ;
      LAYER met4 ;
        RECT 9.585 74.200 9.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 73.795 9.905 74.115 ;
      LAYER met4 ;
        RECT 9.585 73.795 9.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 73.390 9.905 73.710 ;
      LAYER met4 ;
        RECT 9.585 73.390 9.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 72.985 9.905 73.305 ;
      LAYER met4 ;
        RECT 9.585 72.985 9.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 72.575 9.905 72.895 ;
      LAYER met4 ;
        RECT 9.585 72.575 9.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 72.165 9.905 72.485 ;
      LAYER met4 ;
        RECT 9.585 72.165 9.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 71.755 9.905 72.075 ;
      LAYER met4 ;
        RECT 9.585 71.755 9.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 71.345 9.905 71.665 ;
      LAYER met4 ;
        RECT 9.585 71.345 9.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 70.935 9.905 71.255 ;
      LAYER met4 ;
        RECT 9.585 70.935 9.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 70.525 9.905 70.845 ;
      LAYER met4 ;
        RECT 9.585 70.525 9.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 70.115 9.905 70.435 ;
      LAYER met4 ;
        RECT 9.585 70.115 9.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 69.705 9.905 70.025 ;
      LAYER met4 ;
        RECT 9.585 69.705 9.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 69.295 9.905 69.615 ;
      LAYER met4 ;
        RECT 9.585 69.295 9.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 68.885 9.905 69.205 ;
      LAYER met4 ;
        RECT 9.585 68.885 9.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 68.475 9.905 68.795 ;
      LAYER met4 ;
        RECT 9.585 68.475 9.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.585 68.065 9.905 68.385 ;
      LAYER met4 ;
        RECT 9.585 68.065 9.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 22.160 9.800 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 21.730 9.800 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 21.300 9.800 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 20.870 9.800 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 20.440 9.800 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 20.010 9.800 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 19.580 9.800 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 19.150 9.800 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 18.720 9.800 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 18.290 9.800 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.600 17.860 9.800 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 92.635 9.605 92.955 ;
      LAYER met4 ;
        RECT 9.285 92.635 9.605 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 92.225 9.605 92.545 ;
      LAYER met4 ;
        RECT 9.285 92.225 9.605 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 91.815 9.605 92.135 ;
      LAYER met4 ;
        RECT 9.285 91.815 9.605 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 91.405 9.605 91.725 ;
      LAYER met4 ;
        RECT 9.285 91.405 9.605 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 90.995 9.605 91.315 ;
      LAYER met4 ;
        RECT 9.285 90.995 9.605 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 90.585 9.605 90.905 ;
      LAYER met4 ;
        RECT 9.285 90.585 9.605 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 90.175 9.605 90.495 ;
      LAYER met4 ;
        RECT 9.285 90.175 9.605 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 89.765 9.605 90.085 ;
      LAYER met4 ;
        RECT 9.285 89.765 9.605 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 89.355 9.605 89.675 ;
      LAYER met4 ;
        RECT 9.285 89.355 9.605 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 88.945 9.605 89.265 ;
      LAYER met4 ;
        RECT 9.285 88.945 9.605 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 88.535 9.605 88.855 ;
      LAYER met4 ;
        RECT 9.285 88.535 9.605 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 88.125 9.605 88.445 ;
      LAYER met4 ;
        RECT 9.285 88.125 9.605 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 87.715 9.605 88.035 ;
      LAYER met4 ;
        RECT 9.285 87.715 9.605 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 87.305 9.605 87.625 ;
      LAYER met4 ;
        RECT 9.285 87.305 9.605 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 86.895 9.605 87.215 ;
      LAYER met4 ;
        RECT 9.285 86.895 9.605 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 86.485 9.605 86.805 ;
      LAYER met4 ;
        RECT 9.285 86.485 9.605 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 86.075 9.605 86.395 ;
      LAYER met4 ;
        RECT 9.285 86.075 9.605 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 85.665 9.605 85.985 ;
      LAYER met4 ;
        RECT 9.285 85.665 9.605 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 85.255 9.605 85.575 ;
      LAYER met4 ;
        RECT 9.285 85.255 9.605 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 84.845 9.605 85.165 ;
      LAYER met4 ;
        RECT 9.285 84.845 9.605 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 84.435 9.605 84.755 ;
      LAYER met4 ;
        RECT 9.285 84.435 9.605 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 84.025 9.605 84.345 ;
      LAYER met4 ;
        RECT 9.285 84.025 9.605 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 83.615 9.605 83.935 ;
      LAYER met4 ;
        RECT 9.285 83.615 9.605 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 83.205 9.605 83.525 ;
      LAYER met4 ;
        RECT 9.285 83.205 9.605 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.285 82.795 9.605 83.115 ;
      LAYER met4 ;
        RECT 9.285 82.795 9.605 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 82.300 9.505 82.620 ;
      LAYER met4 ;
        RECT 9.185 82.300 9.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 81.895 9.505 82.215 ;
      LAYER met4 ;
        RECT 9.185 81.895 9.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 81.490 9.505 81.810 ;
      LAYER met4 ;
        RECT 9.185 81.490 9.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 81.085 9.505 81.405 ;
      LAYER met4 ;
        RECT 9.185 81.085 9.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 80.680 9.505 81.000 ;
      LAYER met4 ;
        RECT 9.185 80.680 9.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 80.275 9.505 80.595 ;
      LAYER met4 ;
        RECT 9.185 80.275 9.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 79.870 9.505 80.190 ;
      LAYER met4 ;
        RECT 9.185 79.870 9.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 79.465 9.505 79.785 ;
      LAYER met4 ;
        RECT 9.185 79.465 9.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 79.060 9.505 79.380 ;
      LAYER met4 ;
        RECT 9.185 79.060 9.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 78.655 9.505 78.975 ;
      LAYER met4 ;
        RECT 9.185 78.655 9.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 78.250 9.505 78.570 ;
      LAYER met4 ;
        RECT 9.185 78.250 9.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 77.845 9.505 78.165 ;
      LAYER met4 ;
        RECT 9.185 77.845 9.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 77.440 9.505 77.760 ;
      LAYER met4 ;
        RECT 9.185 77.440 9.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 77.035 9.505 77.355 ;
      LAYER met4 ;
        RECT 9.185 77.035 9.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 76.630 9.505 76.950 ;
      LAYER met4 ;
        RECT 9.185 76.630 9.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 76.225 9.505 76.545 ;
      LAYER met4 ;
        RECT 9.185 76.225 9.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 75.820 9.505 76.140 ;
      LAYER met4 ;
        RECT 9.185 75.820 9.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 75.415 9.505 75.735 ;
      LAYER met4 ;
        RECT 9.185 75.415 9.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 75.010 9.505 75.330 ;
      LAYER met4 ;
        RECT 9.185 75.010 9.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 74.605 9.505 74.925 ;
      LAYER met4 ;
        RECT 9.185 74.605 9.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 74.200 9.505 74.520 ;
      LAYER met4 ;
        RECT 9.185 74.200 9.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 73.795 9.505 74.115 ;
      LAYER met4 ;
        RECT 9.185 73.795 9.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 73.390 9.505 73.710 ;
      LAYER met4 ;
        RECT 9.185 73.390 9.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 72.985 9.505 73.305 ;
      LAYER met4 ;
        RECT 9.185 72.985 9.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 72.575 9.505 72.895 ;
      LAYER met4 ;
        RECT 9.185 72.575 9.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 72.165 9.505 72.485 ;
      LAYER met4 ;
        RECT 9.185 72.165 9.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 71.755 9.505 72.075 ;
      LAYER met4 ;
        RECT 9.185 71.755 9.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 71.345 9.505 71.665 ;
      LAYER met4 ;
        RECT 9.185 71.345 9.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 70.935 9.505 71.255 ;
      LAYER met4 ;
        RECT 9.185 70.935 9.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 70.525 9.505 70.845 ;
      LAYER met4 ;
        RECT 9.185 70.525 9.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 70.115 9.505 70.435 ;
      LAYER met4 ;
        RECT 9.185 70.115 9.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 69.705 9.505 70.025 ;
      LAYER met4 ;
        RECT 9.185 69.705 9.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 69.295 9.505 69.615 ;
      LAYER met4 ;
        RECT 9.185 69.295 9.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 68.885 9.505 69.205 ;
      LAYER met4 ;
        RECT 9.185 68.885 9.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 68.475 9.505 68.795 ;
      LAYER met4 ;
        RECT 9.185 68.475 9.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.185 68.065 9.505 68.385 ;
      LAYER met4 ;
        RECT 9.185 68.065 9.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 22.160 9.395 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 21.730 9.395 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 21.300 9.395 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 20.870 9.395 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 20.440 9.395 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 20.010 9.395 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 19.580 9.395 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 19.150 9.395 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 18.720 9.395 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 18.290 9.395 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.195 17.860 9.395 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 92.635 9.195 92.955 ;
      LAYER met4 ;
        RECT 8.875 92.635 9.195 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 92.225 9.195 92.545 ;
      LAYER met4 ;
        RECT 8.875 92.225 9.195 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 91.815 9.195 92.135 ;
      LAYER met4 ;
        RECT 8.875 91.815 9.195 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 91.405 9.195 91.725 ;
      LAYER met4 ;
        RECT 8.875 91.405 9.195 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 90.995 9.195 91.315 ;
      LAYER met4 ;
        RECT 8.875 90.995 9.195 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 90.585 9.195 90.905 ;
      LAYER met4 ;
        RECT 8.875 90.585 9.195 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 90.175 9.195 90.495 ;
      LAYER met4 ;
        RECT 8.875 90.175 9.195 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 89.765 9.195 90.085 ;
      LAYER met4 ;
        RECT 8.875 89.765 9.195 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 89.355 9.195 89.675 ;
      LAYER met4 ;
        RECT 8.875 89.355 9.195 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 88.945 9.195 89.265 ;
      LAYER met4 ;
        RECT 8.875 88.945 9.195 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 88.535 9.195 88.855 ;
      LAYER met4 ;
        RECT 8.875 88.535 9.195 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 88.125 9.195 88.445 ;
      LAYER met4 ;
        RECT 8.875 88.125 9.195 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 87.715 9.195 88.035 ;
      LAYER met4 ;
        RECT 8.875 87.715 9.195 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 87.305 9.195 87.625 ;
      LAYER met4 ;
        RECT 8.875 87.305 9.195 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 86.895 9.195 87.215 ;
      LAYER met4 ;
        RECT 8.875 86.895 9.195 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 86.485 9.195 86.805 ;
      LAYER met4 ;
        RECT 8.875 86.485 9.195 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 86.075 9.195 86.395 ;
      LAYER met4 ;
        RECT 8.875 86.075 9.195 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 85.665 9.195 85.985 ;
      LAYER met4 ;
        RECT 8.875 85.665 9.195 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 85.255 9.195 85.575 ;
      LAYER met4 ;
        RECT 8.875 85.255 9.195 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 84.845 9.195 85.165 ;
      LAYER met4 ;
        RECT 8.875 84.845 9.195 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 84.435 9.195 84.755 ;
      LAYER met4 ;
        RECT 8.875 84.435 9.195 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 84.025 9.195 84.345 ;
      LAYER met4 ;
        RECT 8.875 84.025 9.195 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 83.615 9.195 83.935 ;
      LAYER met4 ;
        RECT 8.875 83.615 9.195 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 83.205 9.195 83.525 ;
      LAYER met4 ;
        RECT 8.875 83.205 9.195 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.875 82.795 9.195 83.115 ;
      LAYER met4 ;
        RECT 8.875 82.795 9.195 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 82.300 9.105 82.620 ;
      LAYER met4 ;
        RECT 8.785 82.300 9.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 81.895 9.105 82.215 ;
      LAYER met4 ;
        RECT 8.785 81.895 9.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 81.490 9.105 81.810 ;
      LAYER met4 ;
        RECT 8.785 81.490 9.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 81.085 9.105 81.405 ;
      LAYER met4 ;
        RECT 8.785 81.085 9.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 80.680 9.105 81.000 ;
      LAYER met4 ;
        RECT 8.785 80.680 9.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 80.275 9.105 80.595 ;
      LAYER met4 ;
        RECT 8.785 80.275 9.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 79.870 9.105 80.190 ;
      LAYER met4 ;
        RECT 8.785 79.870 9.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 79.465 9.105 79.785 ;
      LAYER met4 ;
        RECT 8.785 79.465 9.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 79.060 9.105 79.380 ;
      LAYER met4 ;
        RECT 8.785 79.060 9.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 78.655 9.105 78.975 ;
      LAYER met4 ;
        RECT 8.785 78.655 9.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 78.250 9.105 78.570 ;
      LAYER met4 ;
        RECT 8.785 78.250 9.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 77.845 9.105 78.165 ;
      LAYER met4 ;
        RECT 8.785 77.845 9.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 77.440 9.105 77.760 ;
      LAYER met4 ;
        RECT 8.785 77.440 9.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 77.035 9.105 77.355 ;
      LAYER met4 ;
        RECT 8.785 77.035 9.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 76.630 9.105 76.950 ;
      LAYER met4 ;
        RECT 8.785 76.630 9.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 76.225 9.105 76.545 ;
      LAYER met4 ;
        RECT 8.785 76.225 9.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 75.820 9.105 76.140 ;
      LAYER met4 ;
        RECT 8.785 75.820 9.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 75.415 9.105 75.735 ;
      LAYER met4 ;
        RECT 8.785 75.415 9.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 75.010 9.105 75.330 ;
      LAYER met4 ;
        RECT 8.785 75.010 9.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 74.605 9.105 74.925 ;
      LAYER met4 ;
        RECT 8.785 74.605 9.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 74.200 9.105 74.520 ;
      LAYER met4 ;
        RECT 8.785 74.200 9.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 73.795 9.105 74.115 ;
      LAYER met4 ;
        RECT 8.785 73.795 9.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 73.390 9.105 73.710 ;
      LAYER met4 ;
        RECT 8.785 73.390 9.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 72.985 9.105 73.305 ;
      LAYER met4 ;
        RECT 8.785 72.985 9.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 72.575 9.105 72.895 ;
      LAYER met4 ;
        RECT 8.785 72.575 9.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 72.165 9.105 72.485 ;
      LAYER met4 ;
        RECT 8.785 72.165 9.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 71.755 9.105 72.075 ;
      LAYER met4 ;
        RECT 8.785 71.755 9.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 71.345 9.105 71.665 ;
      LAYER met4 ;
        RECT 8.785 71.345 9.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 70.935 9.105 71.255 ;
      LAYER met4 ;
        RECT 8.785 70.935 9.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 70.525 9.105 70.845 ;
      LAYER met4 ;
        RECT 8.785 70.525 9.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 70.115 9.105 70.435 ;
      LAYER met4 ;
        RECT 8.785 70.115 9.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 69.705 9.105 70.025 ;
      LAYER met4 ;
        RECT 8.785 69.705 9.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 69.295 9.105 69.615 ;
      LAYER met4 ;
        RECT 8.785 69.295 9.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 68.885 9.105 69.205 ;
      LAYER met4 ;
        RECT 8.785 68.885 9.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 68.475 9.105 68.795 ;
      LAYER met4 ;
        RECT 8.785 68.475 9.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.785 68.065 9.105 68.385 ;
      LAYER met4 ;
        RECT 8.785 68.065 9.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 22.160 8.990 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 21.730 8.990 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 21.300 8.990 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 20.870 8.990 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 20.440 8.990 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 20.010 8.990 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 19.580 8.990 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 19.150 8.990 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 18.720 8.990 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 18.290 8.990 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.790 17.860 8.990 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 92.635 8.785 92.955 ;
      LAYER met4 ;
        RECT 8.465 92.635 8.785 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 92.225 8.785 92.545 ;
      LAYER met4 ;
        RECT 8.465 92.225 8.785 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 91.815 8.785 92.135 ;
      LAYER met4 ;
        RECT 8.465 91.815 8.785 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 91.405 8.785 91.725 ;
      LAYER met4 ;
        RECT 8.465 91.405 8.785 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 90.995 8.785 91.315 ;
      LAYER met4 ;
        RECT 8.465 90.995 8.785 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 90.585 8.785 90.905 ;
      LAYER met4 ;
        RECT 8.465 90.585 8.785 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 90.175 8.785 90.495 ;
      LAYER met4 ;
        RECT 8.465 90.175 8.785 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 89.765 8.785 90.085 ;
      LAYER met4 ;
        RECT 8.465 89.765 8.785 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 89.355 8.785 89.675 ;
      LAYER met4 ;
        RECT 8.465 89.355 8.785 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 88.945 8.785 89.265 ;
      LAYER met4 ;
        RECT 8.465 88.945 8.785 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 88.535 8.785 88.855 ;
      LAYER met4 ;
        RECT 8.465 88.535 8.785 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 88.125 8.785 88.445 ;
      LAYER met4 ;
        RECT 8.465 88.125 8.785 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 87.715 8.785 88.035 ;
      LAYER met4 ;
        RECT 8.465 87.715 8.785 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 87.305 8.785 87.625 ;
      LAYER met4 ;
        RECT 8.465 87.305 8.785 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 86.895 8.785 87.215 ;
      LAYER met4 ;
        RECT 8.465 86.895 8.785 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 86.485 8.785 86.805 ;
      LAYER met4 ;
        RECT 8.465 86.485 8.785 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 86.075 8.785 86.395 ;
      LAYER met4 ;
        RECT 8.465 86.075 8.785 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 85.665 8.785 85.985 ;
      LAYER met4 ;
        RECT 8.465 85.665 8.785 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 85.255 8.785 85.575 ;
      LAYER met4 ;
        RECT 8.465 85.255 8.785 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 84.845 8.785 85.165 ;
      LAYER met4 ;
        RECT 8.465 84.845 8.785 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 84.435 8.785 84.755 ;
      LAYER met4 ;
        RECT 8.465 84.435 8.785 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 84.025 8.785 84.345 ;
      LAYER met4 ;
        RECT 8.465 84.025 8.785 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 83.615 8.785 83.935 ;
      LAYER met4 ;
        RECT 8.465 83.615 8.785 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 83.205 8.785 83.525 ;
      LAYER met4 ;
        RECT 8.465 83.205 8.785 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.465 82.795 8.785 83.115 ;
      LAYER met4 ;
        RECT 8.465 82.795 8.785 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 82.300 8.705 82.620 ;
      LAYER met4 ;
        RECT 8.385 82.300 8.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 81.895 8.705 82.215 ;
      LAYER met4 ;
        RECT 8.385 81.895 8.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 81.490 8.705 81.810 ;
      LAYER met4 ;
        RECT 8.385 81.490 8.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 81.085 8.705 81.405 ;
      LAYER met4 ;
        RECT 8.385 81.085 8.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 80.680 8.705 81.000 ;
      LAYER met4 ;
        RECT 8.385 80.680 8.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 80.275 8.705 80.595 ;
      LAYER met4 ;
        RECT 8.385 80.275 8.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 79.870 8.705 80.190 ;
      LAYER met4 ;
        RECT 8.385 79.870 8.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 79.465 8.705 79.785 ;
      LAYER met4 ;
        RECT 8.385 79.465 8.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 79.060 8.705 79.380 ;
      LAYER met4 ;
        RECT 8.385 79.060 8.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 78.655 8.705 78.975 ;
      LAYER met4 ;
        RECT 8.385 78.655 8.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 78.250 8.705 78.570 ;
      LAYER met4 ;
        RECT 8.385 78.250 8.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 77.845 8.705 78.165 ;
      LAYER met4 ;
        RECT 8.385 77.845 8.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 77.440 8.705 77.760 ;
      LAYER met4 ;
        RECT 8.385 77.440 8.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 77.035 8.705 77.355 ;
      LAYER met4 ;
        RECT 8.385 77.035 8.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 76.630 8.705 76.950 ;
      LAYER met4 ;
        RECT 8.385 76.630 8.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 76.225 8.705 76.545 ;
      LAYER met4 ;
        RECT 8.385 76.225 8.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 75.820 8.705 76.140 ;
      LAYER met4 ;
        RECT 8.385 75.820 8.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 75.415 8.705 75.735 ;
      LAYER met4 ;
        RECT 8.385 75.415 8.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 75.010 8.705 75.330 ;
      LAYER met4 ;
        RECT 8.385 75.010 8.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 74.605 8.705 74.925 ;
      LAYER met4 ;
        RECT 8.385 74.605 8.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 74.200 8.705 74.520 ;
      LAYER met4 ;
        RECT 8.385 74.200 8.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 73.795 8.705 74.115 ;
      LAYER met4 ;
        RECT 8.385 73.795 8.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 73.390 8.705 73.710 ;
      LAYER met4 ;
        RECT 8.385 73.390 8.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 72.985 8.705 73.305 ;
      LAYER met4 ;
        RECT 8.385 72.985 8.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 72.575 8.705 72.895 ;
      LAYER met4 ;
        RECT 8.385 72.575 8.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 72.165 8.705 72.485 ;
      LAYER met4 ;
        RECT 8.385 72.165 8.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 71.755 8.705 72.075 ;
      LAYER met4 ;
        RECT 8.385 71.755 8.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 71.345 8.705 71.665 ;
      LAYER met4 ;
        RECT 8.385 71.345 8.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 70.935 8.705 71.255 ;
      LAYER met4 ;
        RECT 8.385 70.935 8.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 70.525 8.705 70.845 ;
      LAYER met4 ;
        RECT 8.385 70.525 8.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 70.115 8.705 70.435 ;
      LAYER met4 ;
        RECT 8.385 70.115 8.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 69.705 8.705 70.025 ;
      LAYER met4 ;
        RECT 8.385 69.705 8.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 69.295 8.705 69.615 ;
      LAYER met4 ;
        RECT 8.385 69.295 8.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 68.885 8.705 69.205 ;
      LAYER met4 ;
        RECT 8.385 68.885 8.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 68.475 8.705 68.795 ;
      LAYER met4 ;
        RECT 8.385 68.475 8.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 68.065 8.705 68.385 ;
      LAYER met4 ;
        RECT 8.385 68.065 8.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 22.160 8.585 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 21.730 8.585 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 21.300 8.585 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 20.870 8.585 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 20.440 8.585 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 20.010 8.585 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 19.580 8.585 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 19.150 8.585 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 18.720 8.585 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 18.290 8.585 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.385 17.860 8.585 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 92.635 8.375 92.955 ;
      LAYER met4 ;
        RECT 8.055 92.635 8.375 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 92.225 8.375 92.545 ;
      LAYER met4 ;
        RECT 8.055 92.225 8.375 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 91.815 8.375 92.135 ;
      LAYER met4 ;
        RECT 8.055 91.815 8.375 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 91.405 8.375 91.725 ;
      LAYER met4 ;
        RECT 8.055 91.405 8.375 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 90.995 8.375 91.315 ;
      LAYER met4 ;
        RECT 8.055 90.995 8.375 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 90.585 8.375 90.905 ;
      LAYER met4 ;
        RECT 8.055 90.585 8.375 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 90.175 8.375 90.495 ;
      LAYER met4 ;
        RECT 8.055 90.175 8.375 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 89.765 8.375 90.085 ;
      LAYER met4 ;
        RECT 8.055 89.765 8.375 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 89.355 8.375 89.675 ;
      LAYER met4 ;
        RECT 8.055 89.355 8.375 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 88.945 8.375 89.265 ;
      LAYER met4 ;
        RECT 8.055 88.945 8.375 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 88.535 8.375 88.855 ;
      LAYER met4 ;
        RECT 8.055 88.535 8.375 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 88.125 8.375 88.445 ;
      LAYER met4 ;
        RECT 8.055 88.125 8.375 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 87.715 8.375 88.035 ;
      LAYER met4 ;
        RECT 8.055 87.715 8.375 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 87.305 8.375 87.625 ;
      LAYER met4 ;
        RECT 8.055 87.305 8.375 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 86.895 8.375 87.215 ;
      LAYER met4 ;
        RECT 8.055 86.895 8.375 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 86.485 8.375 86.805 ;
      LAYER met4 ;
        RECT 8.055 86.485 8.375 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 86.075 8.375 86.395 ;
      LAYER met4 ;
        RECT 8.055 86.075 8.375 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 85.665 8.375 85.985 ;
      LAYER met4 ;
        RECT 8.055 85.665 8.375 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 85.255 8.375 85.575 ;
      LAYER met4 ;
        RECT 8.055 85.255 8.375 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 84.845 8.375 85.165 ;
      LAYER met4 ;
        RECT 8.055 84.845 8.375 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 84.435 8.375 84.755 ;
      LAYER met4 ;
        RECT 8.055 84.435 8.375 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 84.025 8.375 84.345 ;
      LAYER met4 ;
        RECT 8.055 84.025 8.375 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 83.615 8.375 83.935 ;
      LAYER met4 ;
        RECT 8.055 83.615 8.375 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 83.205 8.375 83.525 ;
      LAYER met4 ;
        RECT 8.055 83.205 8.375 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.055 82.795 8.375 83.115 ;
      LAYER met4 ;
        RECT 8.055 82.795 8.375 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 82.300 8.305 82.620 ;
      LAYER met4 ;
        RECT 7.985 82.300 8.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 81.895 8.305 82.215 ;
      LAYER met4 ;
        RECT 7.985 81.895 8.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 81.490 8.305 81.810 ;
      LAYER met4 ;
        RECT 7.985 81.490 8.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 81.085 8.305 81.405 ;
      LAYER met4 ;
        RECT 7.985 81.085 8.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 80.680 8.305 81.000 ;
      LAYER met4 ;
        RECT 7.985 80.680 8.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 80.275 8.305 80.595 ;
      LAYER met4 ;
        RECT 7.985 80.275 8.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 79.870 8.305 80.190 ;
      LAYER met4 ;
        RECT 7.985 79.870 8.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 79.465 8.305 79.785 ;
      LAYER met4 ;
        RECT 7.985 79.465 8.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 79.060 8.305 79.380 ;
      LAYER met4 ;
        RECT 7.985 79.060 8.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 78.655 8.305 78.975 ;
      LAYER met4 ;
        RECT 7.985 78.655 8.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 78.250 8.305 78.570 ;
      LAYER met4 ;
        RECT 7.985 78.250 8.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 77.845 8.305 78.165 ;
      LAYER met4 ;
        RECT 7.985 77.845 8.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 77.440 8.305 77.760 ;
      LAYER met4 ;
        RECT 7.985 77.440 8.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 77.035 8.305 77.355 ;
      LAYER met4 ;
        RECT 7.985 77.035 8.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 76.630 8.305 76.950 ;
      LAYER met4 ;
        RECT 7.985 76.630 8.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 76.225 8.305 76.545 ;
      LAYER met4 ;
        RECT 7.985 76.225 8.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 75.820 8.305 76.140 ;
      LAYER met4 ;
        RECT 7.985 75.820 8.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 75.415 8.305 75.735 ;
      LAYER met4 ;
        RECT 7.985 75.415 8.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 75.010 8.305 75.330 ;
      LAYER met4 ;
        RECT 7.985 75.010 8.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 74.605 8.305 74.925 ;
      LAYER met4 ;
        RECT 7.985 74.605 8.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 74.200 8.305 74.520 ;
      LAYER met4 ;
        RECT 7.985 74.200 8.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 73.795 8.305 74.115 ;
      LAYER met4 ;
        RECT 7.985 73.795 8.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 73.390 8.305 73.710 ;
      LAYER met4 ;
        RECT 7.985 73.390 8.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 72.985 8.305 73.305 ;
      LAYER met4 ;
        RECT 7.985 72.985 8.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 72.575 8.305 72.895 ;
      LAYER met4 ;
        RECT 7.985 72.575 8.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 72.165 8.305 72.485 ;
      LAYER met4 ;
        RECT 7.985 72.165 8.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 71.755 8.305 72.075 ;
      LAYER met4 ;
        RECT 7.985 71.755 8.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 71.345 8.305 71.665 ;
      LAYER met4 ;
        RECT 7.985 71.345 8.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 70.935 8.305 71.255 ;
      LAYER met4 ;
        RECT 7.985 70.935 8.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 70.525 8.305 70.845 ;
      LAYER met4 ;
        RECT 7.985 70.525 8.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 70.115 8.305 70.435 ;
      LAYER met4 ;
        RECT 7.985 70.115 8.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 69.705 8.305 70.025 ;
      LAYER met4 ;
        RECT 7.985 69.705 8.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 69.295 8.305 69.615 ;
      LAYER met4 ;
        RECT 7.985 69.295 8.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 68.885 8.305 69.205 ;
      LAYER met4 ;
        RECT 7.985 68.885 8.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 68.475 8.305 68.795 ;
      LAYER met4 ;
        RECT 7.985 68.475 8.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.985 68.065 8.305 68.385 ;
      LAYER met4 ;
        RECT 7.985 68.065 8.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 22.160 8.180 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 21.730 8.180 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 21.300 8.180 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 20.870 8.180 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 20.440 8.180 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 20.010 8.180 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 19.580 8.180 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 19.150 8.180 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 18.720 8.180 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 18.290 8.180 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.980 17.860 8.180 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 92.635 7.965 92.955 ;
      LAYER met4 ;
        RECT 7.645 92.635 7.965 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 92.225 7.965 92.545 ;
      LAYER met4 ;
        RECT 7.645 92.225 7.965 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 91.815 7.965 92.135 ;
      LAYER met4 ;
        RECT 7.645 91.815 7.965 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 91.405 7.965 91.725 ;
      LAYER met4 ;
        RECT 7.645 91.405 7.965 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 90.995 7.965 91.315 ;
      LAYER met4 ;
        RECT 7.645 90.995 7.965 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 90.585 7.965 90.905 ;
      LAYER met4 ;
        RECT 7.645 90.585 7.965 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 90.175 7.965 90.495 ;
      LAYER met4 ;
        RECT 7.645 90.175 7.965 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 89.765 7.965 90.085 ;
      LAYER met4 ;
        RECT 7.645 89.765 7.965 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 89.355 7.965 89.675 ;
      LAYER met4 ;
        RECT 7.645 89.355 7.965 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 88.945 7.965 89.265 ;
      LAYER met4 ;
        RECT 7.645 88.945 7.965 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 88.535 7.965 88.855 ;
      LAYER met4 ;
        RECT 7.645 88.535 7.965 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 88.125 7.965 88.445 ;
      LAYER met4 ;
        RECT 7.645 88.125 7.965 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 87.715 7.965 88.035 ;
      LAYER met4 ;
        RECT 7.645 87.715 7.965 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 87.305 7.965 87.625 ;
      LAYER met4 ;
        RECT 7.645 87.305 7.965 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 86.895 7.965 87.215 ;
      LAYER met4 ;
        RECT 7.645 86.895 7.965 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 86.485 7.965 86.805 ;
      LAYER met4 ;
        RECT 7.645 86.485 7.965 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 86.075 7.965 86.395 ;
      LAYER met4 ;
        RECT 7.645 86.075 7.965 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 85.665 7.965 85.985 ;
      LAYER met4 ;
        RECT 7.645 85.665 7.965 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 85.255 7.965 85.575 ;
      LAYER met4 ;
        RECT 7.645 85.255 7.965 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 84.845 7.965 85.165 ;
      LAYER met4 ;
        RECT 7.645 84.845 7.965 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 84.435 7.965 84.755 ;
      LAYER met4 ;
        RECT 7.645 84.435 7.965 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 84.025 7.965 84.345 ;
      LAYER met4 ;
        RECT 7.645 84.025 7.965 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 83.615 7.965 83.935 ;
      LAYER met4 ;
        RECT 7.645 83.615 7.965 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 83.205 7.965 83.525 ;
      LAYER met4 ;
        RECT 7.645 83.205 7.965 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.645 82.795 7.965 83.115 ;
      LAYER met4 ;
        RECT 7.645 82.795 7.965 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 82.300 7.905 82.620 ;
      LAYER met4 ;
        RECT 7.585 82.300 7.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 81.895 7.905 82.215 ;
      LAYER met4 ;
        RECT 7.585 81.895 7.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 81.490 7.905 81.810 ;
      LAYER met4 ;
        RECT 7.585 81.490 7.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 81.085 7.905 81.405 ;
      LAYER met4 ;
        RECT 7.585 81.085 7.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 80.680 7.905 81.000 ;
      LAYER met4 ;
        RECT 7.585 80.680 7.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 80.275 7.905 80.595 ;
      LAYER met4 ;
        RECT 7.585 80.275 7.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 79.870 7.905 80.190 ;
      LAYER met4 ;
        RECT 7.585 79.870 7.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 79.465 7.905 79.785 ;
      LAYER met4 ;
        RECT 7.585 79.465 7.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 79.060 7.905 79.380 ;
      LAYER met4 ;
        RECT 7.585 79.060 7.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 78.655 7.905 78.975 ;
      LAYER met4 ;
        RECT 7.585 78.655 7.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 78.250 7.905 78.570 ;
      LAYER met4 ;
        RECT 7.585 78.250 7.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 77.845 7.905 78.165 ;
      LAYER met4 ;
        RECT 7.585 77.845 7.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 77.440 7.905 77.760 ;
      LAYER met4 ;
        RECT 7.585 77.440 7.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 77.035 7.905 77.355 ;
      LAYER met4 ;
        RECT 7.585 77.035 7.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 76.630 7.905 76.950 ;
      LAYER met4 ;
        RECT 7.585 76.630 7.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 76.225 7.905 76.545 ;
      LAYER met4 ;
        RECT 7.585 76.225 7.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 75.820 7.905 76.140 ;
      LAYER met4 ;
        RECT 7.585 75.820 7.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 75.415 7.905 75.735 ;
      LAYER met4 ;
        RECT 7.585 75.415 7.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 75.010 7.905 75.330 ;
      LAYER met4 ;
        RECT 7.585 75.010 7.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 74.605 7.905 74.925 ;
      LAYER met4 ;
        RECT 7.585 74.605 7.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 74.200 7.905 74.520 ;
      LAYER met4 ;
        RECT 7.585 74.200 7.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 73.795 7.905 74.115 ;
      LAYER met4 ;
        RECT 7.585 73.795 7.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 73.390 7.905 73.710 ;
      LAYER met4 ;
        RECT 7.585 73.390 7.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 72.985 7.905 73.305 ;
      LAYER met4 ;
        RECT 7.585 72.985 7.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 72.575 7.905 72.895 ;
      LAYER met4 ;
        RECT 7.585 72.575 7.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 72.165 7.905 72.485 ;
      LAYER met4 ;
        RECT 7.585 72.165 7.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 71.755 7.905 72.075 ;
      LAYER met4 ;
        RECT 7.585 71.755 7.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 71.345 7.905 71.665 ;
      LAYER met4 ;
        RECT 7.585 71.345 7.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 70.935 7.905 71.255 ;
      LAYER met4 ;
        RECT 7.585 70.935 7.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 70.525 7.905 70.845 ;
      LAYER met4 ;
        RECT 7.585 70.525 7.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 70.115 7.905 70.435 ;
      LAYER met4 ;
        RECT 7.585 70.115 7.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 69.705 7.905 70.025 ;
      LAYER met4 ;
        RECT 7.585 69.705 7.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 69.295 7.905 69.615 ;
      LAYER met4 ;
        RECT 7.585 69.295 7.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 68.885 7.905 69.205 ;
      LAYER met4 ;
        RECT 7.585 68.885 7.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 68.475 7.905 68.795 ;
      LAYER met4 ;
        RECT 7.585 68.475 7.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.585 68.065 7.905 68.385 ;
      LAYER met4 ;
        RECT 7.585 68.065 7.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 22.160 7.775 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 21.730 7.775 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 21.300 7.775 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 20.870 7.775 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 20.440 7.775 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 20.010 7.775 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 19.580 7.775 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 19.150 7.775 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 18.720 7.775 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 18.290 7.775 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.575 17.860 7.775 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 92.635 7.555 92.955 ;
      LAYER met4 ;
        RECT 7.235 92.635 7.555 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 92.225 7.555 92.545 ;
      LAYER met4 ;
        RECT 7.235 92.225 7.555 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 91.815 7.555 92.135 ;
      LAYER met4 ;
        RECT 7.235 91.815 7.555 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 91.405 7.555 91.725 ;
      LAYER met4 ;
        RECT 7.235 91.405 7.555 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 90.995 7.555 91.315 ;
      LAYER met4 ;
        RECT 7.235 90.995 7.555 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 90.585 7.555 90.905 ;
      LAYER met4 ;
        RECT 7.235 90.585 7.555 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 90.175 7.555 90.495 ;
      LAYER met4 ;
        RECT 7.235 90.175 7.555 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 89.765 7.555 90.085 ;
      LAYER met4 ;
        RECT 7.235 89.765 7.555 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 89.355 7.555 89.675 ;
      LAYER met4 ;
        RECT 7.235 89.355 7.555 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 88.945 7.555 89.265 ;
      LAYER met4 ;
        RECT 7.235 88.945 7.555 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 88.535 7.555 88.855 ;
      LAYER met4 ;
        RECT 7.235 88.535 7.555 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 88.125 7.555 88.445 ;
      LAYER met4 ;
        RECT 7.235 88.125 7.555 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 87.715 7.555 88.035 ;
      LAYER met4 ;
        RECT 7.235 87.715 7.555 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 87.305 7.555 87.625 ;
      LAYER met4 ;
        RECT 7.235 87.305 7.555 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 86.895 7.555 87.215 ;
      LAYER met4 ;
        RECT 7.235 86.895 7.555 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 86.485 7.555 86.805 ;
      LAYER met4 ;
        RECT 7.235 86.485 7.555 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 86.075 7.555 86.395 ;
      LAYER met4 ;
        RECT 7.235 86.075 7.555 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 85.665 7.555 85.985 ;
      LAYER met4 ;
        RECT 7.235 85.665 7.555 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 85.255 7.555 85.575 ;
      LAYER met4 ;
        RECT 7.235 85.255 7.555 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 84.845 7.555 85.165 ;
      LAYER met4 ;
        RECT 7.235 84.845 7.555 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 84.435 7.555 84.755 ;
      LAYER met4 ;
        RECT 7.235 84.435 7.555 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 84.025 7.555 84.345 ;
      LAYER met4 ;
        RECT 7.235 84.025 7.555 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 83.615 7.555 83.935 ;
      LAYER met4 ;
        RECT 7.235 83.615 7.555 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 83.205 7.555 83.525 ;
      LAYER met4 ;
        RECT 7.235 83.205 7.555 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.235 82.795 7.555 83.115 ;
      LAYER met4 ;
        RECT 7.235 82.795 7.555 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 82.300 7.505 82.620 ;
      LAYER met4 ;
        RECT 7.185 82.300 7.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 81.895 7.505 82.215 ;
      LAYER met4 ;
        RECT 7.185 81.895 7.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 81.490 7.505 81.810 ;
      LAYER met4 ;
        RECT 7.185 81.490 7.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 81.085 7.505 81.405 ;
      LAYER met4 ;
        RECT 7.185 81.085 7.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 80.680 7.505 81.000 ;
      LAYER met4 ;
        RECT 7.185 80.680 7.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 80.275 7.505 80.595 ;
      LAYER met4 ;
        RECT 7.185 80.275 7.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 79.870 7.505 80.190 ;
      LAYER met4 ;
        RECT 7.185 79.870 7.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 79.465 7.505 79.785 ;
      LAYER met4 ;
        RECT 7.185 79.465 7.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 79.060 7.505 79.380 ;
      LAYER met4 ;
        RECT 7.185 79.060 7.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 78.655 7.505 78.975 ;
      LAYER met4 ;
        RECT 7.185 78.655 7.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 78.250 7.505 78.570 ;
      LAYER met4 ;
        RECT 7.185 78.250 7.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 77.845 7.505 78.165 ;
      LAYER met4 ;
        RECT 7.185 77.845 7.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 77.440 7.505 77.760 ;
      LAYER met4 ;
        RECT 7.185 77.440 7.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 77.035 7.505 77.355 ;
      LAYER met4 ;
        RECT 7.185 77.035 7.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 76.630 7.505 76.950 ;
      LAYER met4 ;
        RECT 7.185 76.630 7.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 76.225 7.505 76.545 ;
      LAYER met4 ;
        RECT 7.185 76.225 7.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 75.820 7.505 76.140 ;
      LAYER met4 ;
        RECT 7.185 75.820 7.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 75.415 7.505 75.735 ;
      LAYER met4 ;
        RECT 7.185 75.415 7.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 75.010 7.505 75.330 ;
      LAYER met4 ;
        RECT 7.185 75.010 7.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 74.605 7.505 74.925 ;
      LAYER met4 ;
        RECT 7.185 74.605 7.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 74.200 7.505 74.520 ;
      LAYER met4 ;
        RECT 7.185 74.200 7.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 73.795 7.505 74.115 ;
      LAYER met4 ;
        RECT 7.185 73.795 7.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 73.390 7.505 73.710 ;
      LAYER met4 ;
        RECT 7.185 73.390 7.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 72.985 7.505 73.305 ;
      LAYER met4 ;
        RECT 7.185 72.985 7.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 72.575 7.505 72.895 ;
      LAYER met4 ;
        RECT 7.185 72.575 7.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 72.165 7.505 72.485 ;
      LAYER met4 ;
        RECT 7.185 72.165 7.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 71.755 7.505 72.075 ;
      LAYER met4 ;
        RECT 7.185 71.755 7.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 71.345 7.505 71.665 ;
      LAYER met4 ;
        RECT 7.185 71.345 7.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 70.935 7.505 71.255 ;
      LAYER met4 ;
        RECT 7.185 70.935 7.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 70.525 7.505 70.845 ;
      LAYER met4 ;
        RECT 7.185 70.525 7.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 70.115 7.505 70.435 ;
      LAYER met4 ;
        RECT 7.185 70.115 7.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 69.705 7.505 70.025 ;
      LAYER met4 ;
        RECT 7.185 69.705 7.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 69.295 7.505 69.615 ;
      LAYER met4 ;
        RECT 7.185 69.295 7.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 68.885 7.505 69.205 ;
      LAYER met4 ;
        RECT 7.185 68.885 7.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 68.475 7.505 68.795 ;
      LAYER met4 ;
        RECT 7.185 68.475 7.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.185 68.065 7.505 68.385 ;
      LAYER met4 ;
        RECT 7.185 68.065 7.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 22.160 7.370 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 21.730 7.370 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 21.300 7.370 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 20.870 7.370 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 20.440 7.370 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 20.010 7.370 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 19.580 7.370 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 19.150 7.370 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 18.720 7.370 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 18.290 7.370 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.170 17.860 7.370 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 92.635 7.145 92.955 ;
      LAYER met4 ;
        RECT 6.825 92.635 7.145 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 92.225 7.145 92.545 ;
      LAYER met4 ;
        RECT 6.825 92.225 7.145 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 91.815 7.145 92.135 ;
      LAYER met4 ;
        RECT 6.825 91.815 7.145 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 91.405 7.145 91.725 ;
      LAYER met4 ;
        RECT 6.825 91.405 7.145 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 90.995 7.145 91.315 ;
      LAYER met4 ;
        RECT 6.825 90.995 7.145 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 90.585 7.145 90.905 ;
      LAYER met4 ;
        RECT 6.825 90.585 7.145 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 90.175 7.145 90.495 ;
      LAYER met4 ;
        RECT 6.825 90.175 7.145 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 89.765 7.145 90.085 ;
      LAYER met4 ;
        RECT 6.825 89.765 7.145 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 89.355 7.145 89.675 ;
      LAYER met4 ;
        RECT 6.825 89.355 7.145 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 88.945 7.145 89.265 ;
      LAYER met4 ;
        RECT 6.825 88.945 7.145 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 88.535 7.145 88.855 ;
      LAYER met4 ;
        RECT 6.825 88.535 7.145 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 88.125 7.145 88.445 ;
      LAYER met4 ;
        RECT 6.825 88.125 7.145 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 87.715 7.145 88.035 ;
      LAYER met4 ;
        RECT 6.825 87.715 7.145 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 87.305 7.145 87.625 ;
      LAYER met4 ;
        RECT 6.825 87.305 7.145 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 86.895 7.145 87.215 ;
      LAYER met4 ;
        RECT 6.825 86.895 7.145 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 86.485 7.145 86.805 ;
      LAYER met4 ;
        RECT 6.825 86.485 7.145 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 86.075 7.145 86.395 ;
      LAYER met4 ;
        RECT 6.825 86.075 7.145 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 85.665 7.145 85.985 ;
      LAYER met4 ;
        RECT 6.825 85.665 7.145 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 85.255 7.145 85.575 ;
      LAYER met4 ;
        RECT 6.825 85.255 7.145 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 84.845 7.145 85.165 ;
      LAYER met4 ;
        RECT 6.825 84.845 7.145 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 84.435 7.145 84.755 ;
      LAYER met4 ;
        RECT 6.825 84.435 7.145 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 84.025 7.145 84.345 ;
      LAYER met4 ;
        RECT 6.825 84.025 7.145 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 83.615 7.145 83.935 ;
      LAYER met4 ;
        RECT 6.825 83.615 7.145 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 83.205 7.145 83.525 ;
      LAYER met4 ;
        RECT 6.825 83.205 7.145 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.825 82.795 7.145 83.115 ;
      LAYER met4 ;
        RECT 6.825 82.795 7.145 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 82.300 7.105 82.620 ;
      LAYER met4 ;
        RECT 6.785 82.300 7.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 81.895 7.105 82.215 ;
      LAYER met4 ;
        RECT 6.785 81.895 7.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 81.490 7.105 81.810 ;
      LAYER met4 ;
        RECT 6.785 81.490 7.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 81.085 7.105 81.405 ;
      LAYER met4 ;
        RECT 6.785 81.085 7.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 80.680 7.105 81.000 ;
      LAYER met4 ;
        RECT 6.785 80.680 7.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 80.275 7.105 80.595 ;
      LAYER met4 ;
        RECT 6.785 80.275 7.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 79.870 7.105 80.190 ;
      LAYER met4 ;
        RECT 6.785 79.870 7.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 79.465 7.105 79.785 ;
      LAYER met4 ;
        RECT 6.785 79.465 7.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 79.060 7.105 79.380 ;
      LAYER met4 ;
        RECT 6.785 79.060 7.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 78.655 7.105 78.975 ;
      LAYER met4 ;
        RECT 6.785 78.655 7.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 78.250 7.105 78.570 ;
      LAYER met4 ;
        RECT 6.785 78.250 7.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 77.845 7.105 78.165 ;
      LAYER met4 ;
        RECT 6.785 77.845 7.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 77.440 7.105 77.760 ;
      LAYER met4 ;
        RECT 6.785 77.440 7.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 77.035 7.105 77.355 ;
      LAYER met4 ;
        RECT 6.785 77.035 7.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 76.630 7.105 76.950 ;
      LAYER met4 ;
        RECT 6.785 76.630 7.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 76.225 7.105 76.545 ;
      LAYER met4 ;
        RECT 6.785 76.225 7.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 75.820 7.105 76.140 ;
      LAYER met4 ;
        RECT 6.785 75.820 7.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 75.415 7.105 75.735 ;
      LAYER met4 ;
        RECT 6.785 75.415 7.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 75.010 7.105 75.330 ;
      LAYER met4 ;
        RECT 6.785 75.010 7.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 74.605 7.105 74.925 ;
      LAYER met4 ;
        RECT 6.785 74.605 7.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 74.200 7.105 74.520 ;
      LAYER met4 ;
        RECT 6.785 74.200 7.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 73.795 7.105 74.115 ;
      LAYER met4 ;
        RECT 6.785 73.795 7.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 73.390 7.105 73.710 ;
      LAYER met4 ;
        RECT 6.785 73.390 7.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 72.985 7.105 73.305 ;
      LAYER met4 ;
        RECT 6.785 72.985 7.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 72.575 7.105 72.895 ;
      LAYER met4 ;
        RECT 6.785 72.575 7.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 72.165 7.105 72.485 ;
      LAYER met4 ;
        RECT 6.785 72.165 7.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 71.755 7.105 72.075 ;
      LAYER met4 ;
        RECT 6.785 71.755 7.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 71.345 7.105 71.665 ;
      LAYER met4 ;
        RECT 6.785 71.345 7.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 70.935 7.105 71.255 ;
      LAYER met4 ;
        RECT 6.785 70.935 7.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 70.525 7.105 70.845 ;
      LAYER met4 ;
        RECT 6.785 70.525 7.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 70.115 7.105 70.435 ;
      LAYER met4 ;
        RECT 6.785 70.115 7.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 69.705 7.105 70.025 ;
      LAYER met4 ;
        RECT 6.785 69.705 7.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 69.295 7.105 69.615 ;
      LAYER met4 ;
        RECT 6.785 69.295 7.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 68.885 7.105 69.205 ;
      LAYER met4 ;
        RECT 6.785 68.885 7.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 68.475 7.105 68.795 ;
      LAYER met4 ;
        RECT 6.785 68.475 7.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.785 68.065 7.105 68.385 ;
      LAYER met4 ;
        RECT 6.785 68.065 7.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 22.160 6.965 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 21.730 6.965 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 21.300 6.965 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 20.870 6.965 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 20.440 6.965 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 20.010 6.965 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 19.580 6.965 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 19.150 6.965 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 18.720 6.965 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 18.290 6.965 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.765 17.860 6.965 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 92.635 6.735 92.955 ;
      LAYER met4 ;
        RECT 6.415 92.635 6.735 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 92.225 6.735 92.545 ;
      LAYER met4 ;
        RECT 6.415 92.225 6.735 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 91.815 6.735 92.135 ;
      LAYER met4 ;
        RECT 6.415 91.815 6.735 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 91.405 6.735 91.725 ;
      LAYER met4 ;
        RECT 6.415 91.405 6.735 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 90.995 6.735 91.315 ;
      LAYER met4 ;
        RECT 6.415 90.995 6.735 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 90.585 6.735 90.905 ;
      LAYER met4 ;
        RECT 6.415 90.585 6.735 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 90.175 6.735 90.495 ;
      LAYER met4 ;
        RECT 6.415 90.175 6.735 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 89.765 6.735 90.085 ;
      LAYER met4 ;
        RECT 6.415 89.765 6.735 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 89.355 6.735 89.675 ;
      LAYER met4 ;
        RECT 6.415 89.355 6.735 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 88.945 6.735 89.265 ;
      LAYER met4 ;
        RECT 6.415 88.945 6.735 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 88.535 6.735 88.855 ;
      LAYER met4 ;
        RECT 6.415 88.535 6.735 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 88.125 6.735 88.445 ;
      LAYER met4 ;
        RECT 6.415 88.125 6.735 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 87.715 6.735 88.035 ;
      LAYER met4 ;
        RECT 6.415 87.715 6.735 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 87.305 6.735 87.625 ;
      LAYER met4 ;
        RECT 6.415 87.305 6.735 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 86.895 6.735 87.215 ;
      LAYER met4 ;
        RECT 6.415 86.895 6.735 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 86.485 6.735 86.805 ;
      LAYER met4 ;
        RECT 6.415 86.485 6.735 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 86.075 6.735 86.395 ;
      LAYER met4 ;
        RECT 6.415 86.075 6.735 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 85.665 6.735 85.985 ;
      LAYER met4 ;
        RECT 6.415 85.665 6.735 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 85.255 6.735 85.575 ;
      LAYER met4 ;
        RECT 6.415 85.255 6.735 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 84.845 6.735 85.165 ;
      LAYER met4 ;
        RECT 6.415 84.845 6.735 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 84.435 6.735 84.755 ;
      LAYER met4 ;
        RECT 6.415 84.435 6.735 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 84.025 6.735 84.345 ;
      LAYER met4 ;
        RECT 6.415 84.025 6.735 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 83.615 6.735 83.935 ;
      LAYER met4 ;
        RECT 6.415 83.615 6.735 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 83.205 6.735 83.525 ;
      LAYER met4 ;
        RECT 6.415 83.205 6.735 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.415 82.795 6.735 83.115 ;
      LAYER met4 ;
        RECT 6.415 82.795 6.735 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 82.300 6.705 82.620 ;
      LAYER met4 ;
        RECT 6.385 82.300 6.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 81.895 6.705 82.215 ;
      LAYER met4 ;
        RECT 6.385 81.895 6.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 81.490 6.705 81.810 ;
      LAYER met4 ;
        RECT 6.385 81.490 6.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 81.085 6.705 81.405 ;
      LAYER met4 ;
        RECT 6.385 81.085 6.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 80.680 6.705 81.000 ;
      LAYER met4 ;
        RECT 6.385 80.680 6.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 80.275 6.705 80.595 ;
      LAYER met4 ;
        RECT 6.385 80.275 6.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 79.870 6.705 80.190 ;
      LAYER met4 ;
        RECT 6.385 79.870 6.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 79.465 6.705 79.785 ;
      LAYER met4 ;
        RECT 6.385 79.465 6.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 79.060 6.705 79.380 ;
      LAYER met4 ;
        RECT 6.385 79.060 6.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 78.655 6.705 78.975 ;
      LAYER met4 ;
        RECT 6.385 78.655 6.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 78.250 6.705 78.570 ;
      LAYER met4 ;
        RECT 6.385 78.250 6.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 77.845 6.705 78.165 ;
      LAYER met4 ;
        RECT 6.385 77.845 6.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 77.440 6.705 77.760 ;
      LAYER met4 ;
        RECT 6.385 77.440 6.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 77.035 6.705 77.355 ;
      LAYER met4 ;
        RECT 6.385 77.035 6.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 76.630 6.705 76.950 ;
      LAYER met4 ;
        RECT 6.385 76.630 6.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 76.225 6.705 76.545 ;
      LAYER met4 ;
        RECT 6.385 76.225 6.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 75.820 6.705 76.140 ;
      LAYER met4 ;
        RECT 6.385 75.820 6.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 75.415 6.705 75.735 ;
      LAYER met4 ;
        RECT 6.385 75.415 6.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 75.010 6.705 75.330 ;
      LAYER met4 ;
        RECT 6.385 75.010 6.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 74.605 6.705 74.925 ;
      LAYER met4 ;
        RECT 6.385 74.605 6.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 74.200 6.705 74.520 ;
      LAYER met4 ;
        RECT 6.385 74.200 6.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 73.795 6.705 74.115 ;
      LAYER met4 ;
        RECT 6.385 73.795 6.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 73.390 6.705 73.710 ;
      LAYER met4 ;
        RECT 6.385 73.390 6.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 72.985 6.705 73.305 ;
      LAYER met4 ;
        RECT 6.385 72.985 6.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 72.575 6.705 72.895 ;
      LAYER met4 ;
        RECT 6.385 72.575 6.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 72.165 6.705 72.485 ;
      LAYER met4 ;
        RECT 6.385 72.165 6.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 71.755 6.705 72.075 ;
      LAYER met4 ;
        RECT 6.385 71.755 6.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 71.345 6.705 71.665 ;
      LAYER met4 ;
        RECT 6.385 71.345 6.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 70.935 6.705 71.255 ;
      LAYER met4 ;
        RECT 6.385 70.935 6.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 70.525 6.705 70.845 ;
      LAYER met4 ;
        RECT 6.385 70.525 6.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 70.115 6.705 70.435 ;
      LAYER met4 ;
        RECT 6.385 70.115 6.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 69.705 6.705 70.025 ;
      LAYER met4 ;
        RECT 6.385 69.705 6.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 69.295 6.705 69.615 ;
      LAYER met4 ;
        RECT 6.385 69.295 6.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 68.885 6.705 69.205 ;
      LAYER met4 ;
        RECT 6.385 68.885 6.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 68.475 6.705 68.795 ;
      LAYER met4 ;
        RECT 6.385 68.475 6.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.385 68.065 6.705 68.385 ;
      LAYER met4 ;
        RECT 6.385 68.065 6.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 22.160 6.560 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 21.730 6.560 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 21.300 6.560 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 20.870 6.560 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 20.440 6.560 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 20.010 6.560 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 19.580 6.560 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 19.150 6.560 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 18.720 6.560 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 18.290 6.560 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.360 17.860 6.560 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 92.635 6.325 92.955 ;
      LAYER met4 ;
        RECT 6.005 92.635 6.325 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 92.225 6.325 92.545 ;
      LAYER met4 ;
        RECT 6.005 92.225 6.325 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 91.815 6.325 92.135 ;
      LAYER met4 ;
        RECT 6.005 91.815 6.325 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 91.405 6.325 91.725 ;
      LAYER met4 ;
        RECT 6.005 91.405 6.325 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 90.995 6.325 91.315 ;
      LAYER met4 ;
        RECT 6.005 90.995 6.325 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 90.585 6.325 90.905 ;
      LAYER met4 ;
        RECT 6.005 90.585 6.325 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 90.175 6.325 90.495 ;
      LAYER met4 ;
        RECT 6.005 90.175 6.325 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 89.765 6.325 90.085 ;
      LAYER met4 ;
        RECT 6.005 89.765 6.325 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 89.355 6.325 89.675 ;
      LAYER met4 ;
        RECT 6.005 89.355 6.325 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 88.945 6.325 89.265 ;
      LAYER met4 ;
        RECT 6.005 88.945 6.325 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 88.535 6.325 88.855 ;
      LAYER met4 ;
        RECT 6.005 88.535 6.325 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 88.125 6.325 88.445 ;
      LAYER met4 ;
        RECT 6.005 88.125 6.325 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 87.715 6.325 88.035 ;
      LAYER met4 ;
        RECT 6.005 87.715 6.325 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 87.305 6.325 87.625 ;
      LAYER met4 ;
        RECT 6.005 87.305 6.325 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 86.895 6.325 87.215 ;
      LAYER met4 ;
        RECT 6.005 86.895 6.325 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 86.485 6.325 86.805 ;
      LAYER met4 ;
        RECT 6.005 86.485 6.325 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 86.075 6.325 86.395 ;
      LAYER met4 ;
        RECT 6.005 86.075 6.325 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 85.665 6.325 85.985 ;
      LAYER met4 ;
        RECT 6.005 85.665 6.325 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 85.255 6.325 85.575 ;
      LAYER met4 ;
        RECT 6.005 85.255 6.325 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 84.845 6.325 85.165 ;
      LAYER met4 ;
        RECT 6.005 84.845 6.325 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 84.435 6.325 84.755 ;
      LAYER met4 ;
        RECT 6.005 84.435 6.325 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 84.025 6.325 84.345 ;
      LAYER met4 ;
        RECT 6.005 84.025 6.325 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 83.615 6.325 83.935 ;
      LAYER met4 ;
        RECT 6.005 83.615 6.325 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 83.205 6.325 83.525 ;
      LAYER met4 ;
        RECT 6.005 83.205 6.325 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.005 82.795 6.325 83.115 ;
      LAYER met4 ;
        RECT 6.005 82.795 6.325 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 82.300 6.305 82.620 ;
      LAYER met4 ;
        RECT 5.985 82.300 6.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 81.895 6.305 82.215 ;
      LAYER met4 ;
        RECT 5.985 81.895 6.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 81.490 6.305 81.810 ;
      LAYER met4 ;
        RECT 5.985 81.490 6.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 81.085 6.305 81.405 ;
      LAYER met4 ;
        RECT 5.985 81.085 6.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 80.680 6.305 81.000 ;
      LAYER met4 ;
        RECT 5.985 80.680 6.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 80.275 6.305 80.595 ;
      LAYER met4 ;
        RECT 5.985 80.275 6.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 79.870 6.305 80.190 ;
      LAYER met4 ;
        RECT 5.985 79.870 6.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 79.465 6.305 79.785 ;
      LAYER met4 ;
        RECT 5.985 79.465 6.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 79.060 6.305 79.380 ;
      LAYER met4 ;
        RECT 5.985 79.060 6.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 78.655 6.305 78.975 ;
      LAYER met4 ;
        RECT 5.985 78.655 6.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 78.250 6.305 78.570 ;
      LAYER met4 ;
        RECT 5.985 78.250 6.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 77.845 6.305 78.165 ;
      LAYER met4 ;
        RECT 5.985 77.845 6.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 77.440 6.305 77.760 ;
      LAYER met4 ;
        RECT 5.985 77.440 6.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 77.035 6.305 77.355 ;
      LAYER met4 ;
        RECT 5.985 77.035 6.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 76.630 6.305 76.950 ;
      LAYER met4 ;
        RECT 5.985 76.630 6.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 76.225 6.305 76.545 ;
      LAYER met4 ;
        RECT 5.985 76.225 6.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 75.820 6.305 76.140 ;
      LAYER met4 ;
        RECT 5.985 75.820 6.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 75.415 6.305 75.735 ;
      LAYER met4 ;
        RECT 5.985 75.415 6.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 75.010 6.305 75.330 ;
      LAYER met4 ;
        RECT 5.985 75.010 6.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 74.605 6.305 74.925 ;
      LAYER met4 ;
        RECT 5.985 74.605 6.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 74.200 6.305 74.520 ;
      LAYER met4 ;
        RECT 5.985 74.200 6.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 73.795 6.305 74.115 ;
      LAYER met4 ;
        RECT 5.985 73.795 6.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 73.390 6.305 73.710 ;
      LAYER met4 ;
        RECT 5.985 73.390 6.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 72.985 6.305 73.305 ;
      LAYER met4 ;
        RECT 5.985 72.985 6.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 72.575 6.305 72.895 ;
      LAYER met4 ;
        RECT 5.985 72.575 6.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 72.165 6.305 72.485 ;
      LAYER met4 ;
        RECT 5.985 72.165 6.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 71.755 6.305 72.075 ;
      LAYER met4 ;
        RECT 5.985 71.755 6.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 71.345 6.305 71.665 ;
      LAYER met4 ;
        RECT 5.985 71.345 6.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 70.935 6.305 71.255 ;
      LAYER met4 ;
        RECT 5.985 70.935 6.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 70.525 6.305 70.845 ;
      LAYER met4 ;
        RECT 5.985 70.525 6.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 70.115 6.305 70.435 ;
      LAYER met4 ;
        RECT 5.985 70.115 6.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 69.705 6.305 70.025 ;
      LAYER met4 ;
        RECT 5.985 69.705 6.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 69.295 6.305 69.615 ;
      LAYER met4 ;
        RECT 5.985 69.295 6.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 68.885 6.305 69.205 ;
      LAYER met4 ;
        RECT 5.985 68.885 6.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 68.475 6.305 68.795 ;
      LAYER met4 ;
        RECT 5.985 68.475 6.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.985 68.065 6.305 68.385 ;
      LAYER met4 ;
        RECT 5.985 68.065 6.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 22.160 6.155 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 21.730 6.155 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 21.300 6.155 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 20.870 6.155 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 20.440 6.155 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 20.010 6.155 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 19.580 6.155 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 19.150 6.155 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 18.720 6.155 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 18.290 6.155 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 17.860 6.155 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 92.635 5.915 92.955 ;
      LAYER met4 ;
        RECT 5.595 92.635 5.915 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 92.225 5.915 92.545 ;
      LAYER met4 ;
        RECT 5.595 92.225 5.915 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 91.815 5.915 92.135 ;
      LAYER met4 ;
        RECT 5.595 91.815 5.915 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 91.405 5.915 91.725 ;
      LAYER met4 ;
        RECT 5.595 91.405 5.915 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 90.995 5.915 91.315 ;
      LAYER met4 ;
        RECT 5.595 90.995 5.915 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 90.585 5.915 90.905 ;
      LAYER met4 ;
        RECT 5.595 90.585 5.915 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 90.175 5.915 90.495 ;
      LAYER met4 ;
        RECT 5.595 90.175 5.915 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 89.765 5.915 90.085 ;
      LAYER met4 ;
        RECT 5.595 89.765 5.915 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 89.355 5.915 89.675 ;
      LAYER met4 ;
        RECT 5.595 89.355 5.915 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 88.945 5.915 89.265 ;
      LAYER met4 ;
        RECT 5.595 88.945 5.915 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 88.535 5.915 88.855 ;
      LAYER met4 ;
        RECT 5.595 88.535 5.915 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 88.125 5.915 88.445 ;
      LAYER met4 ;
        RECT 5.595 88.125 5.915 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 87.715 5.915 88.035 ;
      LAYER met4 ;
        RECT 5.595 87.715 5.915 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 87.305 5.915 87.625 ;
      LAYER met4 ;
        RECT 5.595 87.305 5.915 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 86.895 5.915 87.215 ;
      LAYER met4 ;
        RECT 5.595 86.895 5.915 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 86.485 5.915 86.805 ;
      LAYER met4 ;
        RECT 5.595 86.485 5.915 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 86.075 5.915 86.395 ;
      LAYER met4 ;
        RECT 5.595 86.075 5.915 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 85.665 5.915 85.985 ;
      LAYER met4 ;
        RECT 5.595 85.665 5.915 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 85.255 5.915 85.575 ;
      LAYER met4 ;
        RECT 5.595 85.255 5.915 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 84.845 5.915 85.165 ;
      LAYER met4 ;
        RECT 5.595 84.845 5.915 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 84.435 5.915 84.755 ;
      LAYER met4 ;
        RECT 5.595 84.435 5.915 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 84.025 5.915 84.345 ;
      LAYER met4 ;
        RECT 5.595 84.025 5.915 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 83.615 5.915 83.935 ;
      LAYER met4 ;
        RECT 5.595 83.615 5.915 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 83.205 5.915 83.525 ;
      LAYER met4 ;
        RECT 5.595 83.205 5.915 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.595 82.795 5.915 83.115 ;
      LAYER met4 ;
        RECT 5.595 82.795 5.915 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 82.300 5.905 82.620 ;
      LAYER met4 ;
        RECT 5.585 82.300 5.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 81.895 5.905 82.215 ;
      LAYER met4 ;
        RECT 5.585 81.895 5.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 81.490 5.905 81.810 ;
      LAYER met4 ;
        RECT 5.585 81.490 5.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 81.085 5.905 81.405 ;
      LAYER met4 ;
        RECT 5.585 81.085 5.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 80.680 5.905 81.000 ;
      LAYER met4 ;
        RECT 5.585 80.680 5.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 80.275 5.905 80.595 ;
      LAYER met4 ;
        RECT 5.585 80.275 5.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 79.870 5.905 80.190 ;
      LAYER met4 ;
        RECT 5.585 79.870 5.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 79.465 5.905 79.785 ;
      LAYER met4 ;
        RECT 5.585 79.465 5.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 79.060 5.905 79.380 ;
      LAYER met4 ;
        RECT 5.585 79.060 5.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 78.655 5.905 78.975 ;
      LAYER met4 ;
        RECT 5.585 78.655 5.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 78.250 5.905 78.570 ;
      LAYER met4 ;
        RECT 5.585 78.250 5.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 77.845 5.905 78.165 ;
      LAYER met4 ;
        RECT 5.585 77.845 5.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 77.440 5.905 77.760 ;
      LAYER met4 ;
        RECT 5.585 77.440 5.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 77.035 5.905 77.355 ;
      LAYER met4 ;
        RECT 5.585 77.035 5.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 76.630 5.905 76.950 ;
      LAYER met4 ;
        RECT 5.585 76.630 5.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 76.225 5.905 76.545 ;
      LAYER met4 ;
        RECT 5.585 76.225 5.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 75.820 5.905 76.140 ;
      LAYER met4 ;
        RECT 5.585 75.820 5.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 75.415 5.905 75.735 ;
      LAYER met4 ;
        RECT 5.585 75.415 5.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 75.010 5.905 75.330 ;
      LAYER met4 ;
        RECT 5.585 75.010 5.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 74.605 5.905 74.925 ;
      LAYER met4 ;
        RECT 5.585 74.605 5.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 74.200 5.905 74.520 ;
      LAYER met4 ;
        RECT 5.585 74.200 5.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 73.795 5.905 74.115 ;
      LAYER met4 ;
        RECT 5.585 73.795 5.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 73.390 5.905 73.710 ;
      LAYER met4 ;
        RECT 5.585 73.390 5.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 72.985 5.905 73.305 ;
      LAYER met4 ;
        RECT 5.585 72.985 5.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 72.575 5.905 72.895 ;
      LAYER met4 ;
        RECT 5.585 72.575 5.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 72.165 5.905 72.485 ;
      LAYER met4 ;
        RECT 5.585 72.165 5.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 71.755 5.905 72.075 ;
      LAYER met4 ;
        RECT 5.585 71.755 5.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 71.345 5.905 71.665 ;
      LAYER met4 ;
        RECT 5.585 71.345 5.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 70.935 5.905 71.255 ;
      LAYER met4 ;
        RECT 5.585 70.935 5.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 70.525 5.905 70.845 ;
      LAYER met4 ;
        RECT 5.585 70.525 5.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 70.115 5.905 70.435 ;
      LAYER met4 ;
        RECT 5.585 70.115 5.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 69.705 5.905 70.025 ;
      LAYER met4 ;
        RECT 5.585 69.705 5.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 69.295 5.905 69.615 ;
      LAYER met4 ;
        RECT 5.585 69.295 5.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 68.885 5.905 69.205 ;
      LAYER met4 ;
        RECT 5.585 68.885 5.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 68.475 5.905 68.795 ;
      LAYER met4 ;
        RECT 5.585 68.475 5.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.585 68.065 5.905 68.385 ;
      LAYER met4 ;
        RECT 5.585 68.065 5.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 22.160 5.750 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 21.730 5.750 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 21.300 5.750 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 20.870 5.750 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 20.440 5.750 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 20.010 5.750 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 19.580 5.750 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 19.150 5.750 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 18.720 5.750 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 18.290 5.750 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.550 17.860 5.750 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 92.635 5.505 92.955 ;
      LAYER met4 ;
        RECT 5.185 92.635 5.505 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 92.225 5.505 92.545 ;
      LAYER met4 ;
        RECT 5.185 92.225 5.505 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 91.815 5.505 92.135 ;
      LAYER met4 ;
        RECT 5.185 91.815 5.505 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 91.405 5.505 91.725 ;
      LAYER met4 ;
        RECT 5.185 91.405 5.505 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 90.995 5.505 91.315 ;
      LAYER met4 ;
        RECT 5.185 90.995 5.505 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 90.585 5.505 90.905 ;
      LAYER met4 ;
        RECT 5.185 90.585 5.505 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 90.175 5.505 90.495 ;
      LAYER met4 ;
        RECT 5.185 90.175 5.505 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 89.765 5.505 90.085 ;
      LAYER met4 ;
        RECT 5.185 89.765 5.505 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 89.355 5.505 89.675 ;
      LAYER met4 ;
        RECT 5.185 89.355 5.505 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 88.945 5.505 89.265 ;
      LAYER met4 ;
        RECT 5.185 88.945 5.505 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 88.535 5.505 88.855 ;
      LAYER met4 ;
        RECT 5.185 88.535 5.505 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 88.125 5.505 88.445 ;
      LAYER met4 ;
        RECT 5.185 88.125 5.505 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 87.715 5.505 88.035 ;
      LAYER met4 ;
        RECT 5.185 87.715 5.505 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 87.305 5.505 87.625 ;
      LAYER met4 ;
        RECT 5.185 87.305 5.505 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 86.895 5.505 87.215 ;
      LAYER met4 ;
        RECT 5.185 86.895 5.505 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 86.485 5.505 86.805 ;
      LAYER met4 ;
        RECT 5.185 86.485 5.505 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 86.075 5.505 86.395 ;
      LAYER met4 ;
        RECT 5.185 86.075 5.505 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 85.665 5.505 85.985 ;
      LAYER met4 ;
        RECT 5.185 85.665 5.505 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 85.255 5.505 85.575 ;
      LAYER met4 ;
        RECT 5.185 85.255 5.505 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 84.845 5.505 85.165 ;
      LAYER met4 ;
        RECT 5.185 84.845 5.505 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 84.435 5.505 84.755 ;
      LAYER met4 ;
        RECT 5.185 84.435 5.505 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 84.025 5.505 84.345 ;
      LAYER met4 ;
        RECT 5.185 84.025 5.505 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 83.615 5.505 83.935 ;
      LAYER met4 ;
        RECT 5.185 83.615 5.505 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 83.205 5.505 83.525 ;
      LAYER met4 ;
        RECT 5.185 83.205 5.505 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 82.795 5.505 83.115 ;
      LAYER met4 ;
        RECT 5.185 82.795 5.505 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 82.300 5.505 82.620 ;
      LAYER met4 ;
        RECT 5.185 82.300 5.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 81.895 5.505 82.215 ;
      LAYER met4 ;
        RECT 5.185 81.895 5.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 81.490 5.505 81.810 ;
      LAYER met4 ;
        RECT 5.185 81.490 5.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 81.085 5.505 81.405 ;
      LAYER met4 ;
        RECT 5.185 81.085 5.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 80.680 5.505 81.000 ;
      LAYER met4 ;
        RECT 5.185 80.680 5.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 80.275 5.505 80.595 ;
      LAYER met4 ;
        RECT 5.185 80.275 5.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 79.870 5.505 80.190 ;
      LAYER met4 ;
        RECT 5.185 79.870 5.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 79.465 5.505 79.785 ;
      LAYER met4 ;
        RECT 5.185 79.465 5.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 79.060 5.505 79.380 ;
      LAYER met4 ;
        RECT 5.185 79.060 5.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 78.655 5.505 78.975 ;
      LAYER met4 ;
        RECT 5.185 78.655 5.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 78.250 5.505 78.570 ;
      LAYER met4 ;
        RECT 5.185 78.250 5.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 77.845 5.505 78.165 ;
      LAYER met4 ;
        RECT 5.185 77.845 5.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 77.440 5.505 77.760 ;
      LAYER met4 ;
        RECT 5.185 77.440 5.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 77.035 5.505 77.355 ;
      LAYER met4 ;
        RECT 5.185 77.035 5.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 76.630 5.505 76.950 ;
      LAYER met4 ;
        RECT 5.185 76.630 5.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 76.225 5.505 76.545 ;
      LAYER met4 ;
        RECT 5.185 76.225 5.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 75.820 5.505 76.140 ;
      LAYER met4 ;
        RECT 5.185 75.820 5.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 75.415 5.505 75.735 ;
      LAYER met4 ;
        RECT 5.185 75.415 5.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 75.010 5.505 75.330 ;
      LAYER met4 ;
        RECT 5.185 75.010 5.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 74.605 5.505 74.925 ;
      LAYER met4 ;
        RECT 5.185 74.605 5.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 74.200 5.505 74.520 ;
      LAYER met4 ;
        RECT 5.185 74.200 5.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 73.795 5.505 74.115 ;
      LAYER met4 ;
        RECT 5.185 73.795 5.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 73.390 5.505 73.710 ;
      LAYER met4 ;
        RECT 5.185 73.390 5.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 72.985 5.505 73.305 ;
      LAYER met4 ;
        RECT 5.185 72.985 5.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 72.575 5.505 72.895 ;
      LAYER met4 ;
        RECT 5.185 72.575 5.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 72.165 5.505 72.485 ;
      LAYER met4 ;
        RECT 5.185 72.165 5.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 71.755 5.505 72.075 ;
      LAYER met4 ;
        RECT 5.185 71.755 5.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 71.345 5.505 71.665 ;
      LAYER met4 ;
        RECT 5.185 71.345 5.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 70.935 5.505 71.255 ;
      LAYER met4 ;
        RECT 5.185 70.935 5.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 70.525 5.505 70.845 ;
      LAYER met4 ;
        RECT 5.185 70.525 5.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 70.115 5.505 70.435 ;
      LAYER met4 ;
        RECT 5.185 70.115 5.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 69.705 5.505 70.025 ;
      LAYER met4 ;
        RECT 5.185 69.705 5.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 69.295 5.505 69.615 ;
      LAYER met4 ;
        RECT 5.185 69.295 5.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 68.885 5.505 69.205 ;
      LAYER met4 ;
        RECT 5.185 68.885 5.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 68.475 5.505 68.795 ;
      LAYER met4 ;
        RECT 5.185 68.475 5.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.185 68.065 5.505 68.385 ;
      LAYER met4 ;
        RECT 5.185 68.065 5.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 22.160 5.345 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 21.730 5.345 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 21.300 5.345 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 20.870 5.345 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 20.440 5.345 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 20.010 5.345 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 19.580 5.345 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 19.150 5.345 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 18.720 5.345 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 18.290 5.345 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.145 17.860 5.345 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 82.300 5.105 82.620 ;
      LAYER met4 ;
        RECT 4.785 82.300 5.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 81.895 5.105 82.215 ;
      LAYER met4 ;
        RECT 4.785 81.895 5.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 81.490 5.105 81.810 ;
      LAYER met4 ;
        RECT 4.785 81.490 5.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 81.085 5.105 81.405 ;
      LAYER met4 ;
        RECT 4.785 81.085 5.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 80.680 5.105 81.000 ;
      LAYER met4 ;
        RECT 4.785 80.680 5.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 80.275 5.105 80.595 ;
      LAYER met4 ;
        RECT 4.785 80.275 5.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 79.870 5.105 80.190 ;
      LAYER met4 ;
        RECT 4.785 79.870 5.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 79.465 5.105 79.785 ;
      LAYER met4 ;
        RECT 4.785 79.465 5.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 79.060 5.105 79.380 ;
      LAYER met4 ;
        RECT 4.785 79.060 5.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 78.655 5.105 78.975 ;
      LAYER met4 ;
        RECT 4.785 78.655 5.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 78.250 5.105 78.570 ;
      LAYER met4 ;
        RECT 4.785 78.250 5.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 77.845 5.105 78.165 ;
      LAYER met4 ;
        RECT 4.785 77.845 5.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 77.440 5.105 77.760 ;
      LAYER met4 ;
        RECT 4.785 77.440 5.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 77.035 5.105 77.355 ;
      LAYER met4 ;
        RECT 4.785 77.035 5.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 76.630 5.105 76.950 ;
      LAYER met4 ;
        RECT 4.785 76.630 5.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 76.225 5.105 76.545 ;
      LAYER met4 ;
        RECT 4.785 76.225 5.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 75.820 5.105 76.140 ;
      LAYER met4 ;
        RECT 4.785 75.820 5.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 75.415 5.105 75.735 ;
      LAYER met4 ;
        RECT 4.785 75.415 5.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 75.010 5.105 75.330 ;
      LAYER met4 ;
        RECT 4.785 75.010 5.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 74.605 5.105 74.925 ;
      LAYER met4 ;
        RECT 4.785 74.605 5.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 74.200 5.105 74.520 ;
      LAYER met4 ;
        RECT 4.785 74.200 5.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 73.795 5.105 74.115 ;
      LAYER met4 ;
        RECT 4.785 73.795 5.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 73.390 5.105 73.710 ;
      LAYER met4 ;
        RECT 4.785 73.390 5.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 72.985 5.105 73.305 ;
      LAYER met4 ;
        RECT 4.785 72.985 5.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 72.575 5.105 72.895 ;
      LAYER met4 ;
        RECT 4.785 72.575 5.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 72.165 5.105 72.485 ;
      LAYER met4 ;
        RECT 4.785 72.165 5.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 71.755 5.105 72.075 ;
      LAYER met4 ;
        RECT 4.785 71.755 5.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 71.345 5.105 71.665 ;
      LAYER met4 ;
        RECT 4.785 71.345 5.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 70.935 5.105 71.255 ;
      LAYER met4 ;
        RECT 4.785 70.935 5.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 70.525 5.105 70.845 ;
      LAYER met4 ;
        RECT 4.785 70.525 5.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 70.115 5.105 70.435 ;
      LAYER met4 ;
        RECT 4.785 70.115 5.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 69.705 5.105 70.025 ;
      LAYER met4 ;
        RECT 4.785 69.705 5.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 69.295 5.105 69.615 ;
      LAYER met4 ;
        RECT 4.785 69.295 5.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 68.885 5.105 69.205 ;
      LAYER met4 ;
        RECT 4.785 68.885 5.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 68.475 5.105 68.795 ;
      LAYER met4 ;
        RECT 4.785 68.475 5.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.785 68.065 5.105 68.385 ;
      LAYER met4 ;
        RECT 4.785 68.065 5.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 92.635 5.095 92.955 ;
      LAYER met4 ;
        RECT 4.775 92.635 5.095 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 92.225 5.095 92.545 ;
      LAYER met4 ;
        RECT 4.775 92.225 5.095 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 91.815 5.095 92.135 ;
      LAYER met4 ;
        RECT 4.775 91.815 5.095 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 91.405 5.095 91.725 ;
      LAYER met4 ;
        RECT 4.775 91.405 5.095 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 90.995 5.095 91.315 ;
      LAYER met4 ;
        RECT 4.775 90.995 5.095 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 90.585 5.095 90.905 ;
      LAYER met4 ;
        RECT 4.775 90.585 5.095 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 90.175 5.095 90.495 ;
      LAYER met4 ;
        RECT 4.775 90.175 5.095 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 89.765 5.095 90.085 ;
      LAYER met4 ;
        RECT 4.775 89.765 5.095 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 89.355 5.095 89.675 ;
      LAYER met4 ;
        RECT 4.775 89.355 5.095 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 88.945 5.095 89.265 ;
      LAYER met4 ;
        RECT 4.775 88.945 5.095 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 88.535 5.095 88.855 ;
      LAYER met4 ;
        RECT 4.775 88.535 5.095 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 88.125 5.095 88.445 ;
      LAYER met4 ;
        RECT 4.775 88.125 5.095 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 87.715 5.095 88.035 ;
      LAYER met4 ;
        RECT 4.775 87.715 5.095 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 87.305 5.095 87.625 ;
      LAYER met4 ;
        RECT 4.775 87.305 5.095 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 86.895 5.095 87.215 ;
      LAYER met4 ;
        RECT 4.775 86.895 5.095 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 86.485 5.095 86.805 ;
      LAYER met4 ;
        RECT 4.775 86.485 5.095 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 86.075 5.095 86.395 ;
      LAYER met4 ;
        RECT 4.775 86.075 5.095 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 85.665 5.095 85.985 ;
      LAYER met4 ;
        RECT 4.775 85.665 5.095 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 85.255 5.095 85.575 ;
      LAYER met4 ;
        RECT 4.775 85.255 5.095 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 84.845 5.095 85.165 ;
      LAYER met4 ;
        RECT 4.775 84.845 5.095 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 84.435 5.095 84.755 ;
      LAYER met4 ;
        RECT 4.775 84.435 5.095 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 84.025 5.095 84.345 ;
      LAYER met4 ;
        RECT 4.775 84.025 5.095 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 83.615 5.095 83.935 ;
      LAYER met4 ;
        RECT 4.775 83.615 5.095 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 83.205 5.095 83.525 ;
      LAYER met4 ;
        RECT 4.775 83.205 5.095 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.775 82.795 5.095 83.115 ;
      LAYER met4 ;
        RECT 4.775 82.795 5.095 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 22.160 4.940 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 21.730 4.940 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 21.300 4.940 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 20.870 4.940 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 20.440 4.940 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 20.010 4.940 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 19.580 4.940 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 19.150 4.940 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 18.720 4.940 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 18.290 4.940 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.740 17.860 4.940 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 82.300 4.705 82.620 ;
      LAYER met4 ;
        RECT 4.385 82.300 4.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 81.895 4.705 82.215 ;
      LAYER met4 ;
        RECT 4.385 81.895 4.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 81.490 4.705 81.810 ;
      LAYER met4 ;
        RECT 4.385 81.490 4.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 81.085 4.705 81.405 ;
      LAYER met4 ;
        RECT 4.385 81.085 4.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 80.680 4.705 81.000 ;
      LAYER met4 ;
        RECT 4.385 80.680 4.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 80.275 4.705 80.595 ;
      LAYER met4 ;
        RECT 4.385 80.275 4.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 79.870 4.705 80.190 ;
      LAYER met4 ;
        RECT 4.385 79.870 4.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 79.465 4.705 79.785 ;
      LAYER met4 ;
        RECT 4.385 79.465 4.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 79.060 4.705 79.380 ;
      LAYER met4 ;
        RECT 4.385 79.060 4.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 78.655 4.705 78.975 ;
      LAYER met4 ;
        RECT 4.385 78.655 4.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 78.250 4.705 78.570 ;
      LAYER met4 ;
        RECT 4.385 78.250 4.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 77.845 4.705 78.165 ;
      LAYER met4 ;
        RECT 4.385 77.845 4.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 77.440 4.705 77.760 ;
      LAYER met4 ;
        RECT 4.385 77.440 4.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 77.035 4.705 77.355 ;
      LAYER met4 ;
        RECT 4.385 77.035 4.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 76.630 4.705 76.950 ;
      LAYER met4 ;
        RECT 4.385 76.630 4.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 76.225 4.705 76.545 ;
      LAYER met4 ;
        RECT 4.385 76.225 4.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 75.820 4.705 76.140 ;
      LAYER met4 ;
        RECT 4.385 75.820 4.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 75.415 4.705 75.735 ;
      LAYER met4 ;
        RECT 4.385 75.415 4.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 75.010 4.705 75.330 ;
      LAYER met4 ;
        RECT 4.385 75.010 4.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 74.605 4.705 74.925 ;
      LAYER met4 ;
        RECT 4.385 74.605 4.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 74.200 4.705 74.520 ;
      LAYER met4 ;
        RECT 4.385 74.200 4.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 73.795 4.705 74.115 ;
      LAYER met4 ;
        RECT 4.385 73.795 4.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 73.390 4.705 73.710 ;
      LAYER met4 ;
        RECT 4.385 73.390 4.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 72.985 4.705 73.305 ;
      LAYER met4 ;
        RECT 4.385 72.985 4.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 72.575 4.705 72.895 ;
      LAYER met4 ;
        RECT 4.385 72.575 4.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 72.165 4.705 72.485 ;
      LAYER met4 ;
        RECT 4.385 72.165 4.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 71.755 4.705 72.075 ;
      LAYER met4 ;
        RECT 4.385 71.755 4.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 71.345 4.705 71.665 ;
      LAYER met4 ;
        RECT 4.385 71.345 4.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 70.935 4.705 71.255 ;
      LAYER met4 ;
        RECT 4.385 70.935 4.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 70.525 4.705 70.845 ;
      LAYER met4 ;
        RECT 4.385 70.525 4.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 70.115 4.705 70.435 ;
      LAYER met4 ;
        RECT 4.385 70.115 4.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 69.705 4.705 70.025 ;
      LAYER met4 ;
        RECT 4.385 69.705 4.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 69.295 4.705 69.615 ;
      LAYER met4 ;
        RECT 4.385 69.295 4.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 68.885 4.705 69.205 ;
      LAYER met4 ;
        RECT 4.385 68.885 4.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 68.475 4.705 68.795 ;
      LAYER met4 ;
        RECT 4.385 68.475 4.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.385 68.065 4.705 68.385 ;
      LAYER met4 ;
        RECT 4.385 68.065 4.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 92.635 4.685 92.955 ;
      LAYER met4 ;
        RECT 4.365 92.635 4.685 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 92.225 4.685 92.545 ;
      LAYER met4 ;
        RECT 4.365 92.225 4.685 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 91.815 4.685 92.135 ;
      LAYER met4 ;
        RECT 4.365 91.815 4.685 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 91.405 4.685 91.725 ;
      LAYER met4 ;
        RECT 4.365 91.405 4.685 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 90.995 4.685 91.315 ;
      LAYER met4 ;
        RECT 4.365 90.995 4.685 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 90.585 4.685 90.905 ;
      LAYER met4 ;
        RECT 4.365 90.585 4.685 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 90.175 4.685 90.495 ;
      LAYER met4 ;
        RECT 4.365 90.175 4.685 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 89.765 4.685 90.085 ;
      LAYER met4 ;
        RECT 4.365 89.765 4.685 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 89.355 4.685 89.675 ;
      LAYER met4 ;
        RECT 4.365 89.355 4.685 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 88.945 4.685 89.265 ;
      LAYER met4 ;
        RECT 4.365 88.945 4.685 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 88.535 4.685 88.855 ;
      LAYER met4 ;
        RECT 4.365 88.535 4.685 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 88.125 4.685 88.445 ;
      LAYER met4 ;
        RECT 4.365 88.125 4.685 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 87.715 4.685 88.035 ;
      LAYER met4 ;
        RECT 4.365 87.715 4.685 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 87.305 4.685 87.625 ;
      LAYER met4 ;
        RECT 4.365 87.305 4.685 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 86.895 4.685 87.215 ;
      LAYER met4 ;
        RECT 4.365 86.895 4.685 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 86.485 4.685 86.805 ;
      LAYER met4 ;
        RECT 4.365 86.485 4.685 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 86.075 4.685 86.395 ;
      LAYER met4 ;
        RECT 4.365 86.075 4.685 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 85.665 4.685 85.985 ;
      LAYER met4 ;
        RECT 4.365 85.665 4.685 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 85.255 4.685 85.575 ;
      LAYER met4 ;
        RECT 4.365 85.255 4.685 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 84.845 4.685 85.165 ;
      LAYER met4 ;
        RECT 4.365 84.845 4.685 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 84.435 4.685 84.755 ;
      LAYER met4 ;
        RECT 4.365 84.435 4.685 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 84.025 4.685 84.345 ;
      LAYER met4 ;
        RECT 4.365 84.025 4.685 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 83.615 4.685 83.935 ;
      LAYER met4 ;
        RECT 4.365 83.615 4.685 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 83.205 4.685 83.525 ;
      LAYER met4 ;
        RECT 4.365 83.205 4.685 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.365 82.795 4.685 83.115 ;
      LAYER met4 ;
        RECT 4.365 82.795 4.685 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 22.160 4.535 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 21.730 4.535 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 21.300 4.535 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 20.870 4.535 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 20.440 4.535 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 20.010 4.535 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 19.580 4.535 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 19.150 4.535 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 18.720 4.535 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 18.290 4.535 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.335 17.860 4.535 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 82.300 4.305 82.620 ;
      LAYER met4 ;
        RECT 3.985 82.300 4.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 81.895 4.305 82.215 ;
      LAYER met4 ;
        RECT 3.985 81.895 4.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 81.490 4.305 81.810 ;
      LAYER met4 ;
        RECT 3.985 81.490 4.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 81.085 4.305 81.405 ;
      LAYER met4 ;
        RECT 3.985 81.085 4.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 80.680 4.305 81.000 ;
      LAYER met4 ;
        RECT 3.985 80.680 4.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 80.275 4.305 80.595 ;
      LAYER met4 ;
        RECT 3.985 80.275 4.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 79.870 4.305 80.190 ;
      LAYER met4 ;
        RECT 3.985 79.870 4.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 79.465 4.305 79.785 ;
      LAYER met4 ;
        RECT 3.985 79.465 4.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 79.060 4.305 79.380 ;
      LAYER met4 ;
        RECT 3.985 79.060 4.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 78.655 4.305 78.975 ;
      LAYER met4 ;
        RECT 3.985 78.655 4.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 78.250 4.305 78.570 ;
      LAYER met4 ;
        RECT 3.985 78.250 4.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 77.845 4.305 78.165 ;
      LAYER met4 ;
        RECT 3.985 77.845 4.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 77.440 4.305 77.760 ;
      LAYER met4 ;
        RECT 3.985 77.440 4.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 77.035 4.305 77.355 ;
      LAYER met4 ;
        RECT 3.985 77.035 4.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 76.630 4.305 76.950 ;
      LAYER met4 ;
        RECT 3.985 76.630 4.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 76.225 4.305 76.545 ;
      LAYER met4 ;
        RECT 3.985 76.225 4.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 75.820 4.305 76.140 ;
      LAYER met4 ;
        RECT 3.985 75.820 4.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 75.415 4.305 75.735 ;
      LAYER met4 ;
        RECT 3.985 75.415 4.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 75.010 4.305 75.330 ;
      LAYER met4 ;
        RECT 3.985 75.010 4.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 74.605 4.305 74.925 ;
      LAYER met4 ;
        RECT 3.985 74.605 4.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 74.200 4.305 74.520 ;
      LAYER met4 ;
        RECT 3.985 74.200 4.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 73.795 4.305 74.115 ;
      LAYER met4 ;
        RECT 3.985 73.795 4.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 73.390 4.305 73.710 ;
      LAYER met4 ;
        RECT 3.985 73.390 4.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 72.985 4.305 73.305 ;
      LAYER met4 ;
        RECT 3.985 72.985 4.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 72.575 4.305 72.895 ;
      LAYER met4 ;
        RECT 3.985 72.575 4.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 72.165 4.305 72.485 ;
      LAYER met4 ;
        RECT 3.985 72.165 4.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 71.755 4.305 72.075 ;
      LAYER met4 ;
        RECT 3.985 71.755 4.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 71.345 4.305 71.665 ;
      LAYER met4 ;
        RECT 3.985 71.345 4.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 70.935 4.305 71.255 ;
      LAYER met4 ;
        RECT 3.985 70.935 4.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 70.525 4.305 70.845 ;
      LAYER met4 ;
        RECT 3.985 70.525 4.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 70.115 4.305 70.435 ;
      LAYER met4 ;
        RECT 3.985 70.115 4.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 69.705 4.305 70.025 ;
      LAYER met4 ;
        RECT 3.985 69.705 4.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 69.295 4.305 69.615 ;
      LAYER met4 ;
        RECT 3.985 69.295 4.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 68.885 4.305 69.205 ;
      LAYER met4 ;
        RECT 3.985 68.885 4.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 68.475 4.305 68.795 ;
      LAYER met4 ;
        RECT 3.985 68.475 4.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.985 68.065 4.305 68.385 ;
      LAYER met4 ;
        RECT 3.985 68.065 4.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 92.635 4.275 92.955 ;
      LAYER met4 ;
        RECT 3.955 92.635 4.275 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 92.225 4.275 92.545 ;
      LAYER met4 ;
        RECT 3.955 92.225 4.275 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 91.815 4.275 92.135 ;
      LAYER met4 ;
        RECT 3.955 91.815 4.275 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 91.405 4.275 91.725 ;
      LAYER met4 ;
        RECT 3.955 91.405 4.275 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 90.995 4.275 91.315 ;
      LAYER met4 ;
        RECT 3.955 90.995 4.275 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 90.585 4.275 90.905 ;
      LAYER met4 ;
        RECT 3.955 90.585 4.275 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 90.175 4.275 90.495 ;
      LAYER met4 ;
        RECT 3.955 90.175 4.275 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 89.765 4.275 90.085 ;
      LAYER met4 ;
        RECT 3.955 89.765 4.275 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 89.355 4.275 89.675 ;
      LAYER met4 ;
        RECT 3.955 89.355 4.275 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 88.945 4.275 89.265 ;
      LAYER met4 ;
        RECT 3.955 88.945 4.275 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 88.535 4.275 88.855 ;
      LAYER met4 ;
        RECT 3.955 88.535 4.275 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 88.125 4.275 88.445 ;
      LAYER met4 ;
        RECT 3.955 88.125 4.275 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 87.715 4.275 88.035 ;
      LAYER met4 ;
        RECT 3.955 87.715 4.275 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 87.305 4.275 87.625 ;
      LAYER met4 ;
        RECT 3.955 87.305 4.275 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 86.895 4.275 87.215 ;
      LAYER met4 ;
        RECT 3.955 86.895 4.275 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 86.485 4.275 86.805 ;
      LAYER met4 ;
        RECT 3.955 86.485 4.275 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 86.075 4.275 86.395 ;
      LAYER met4 ;
        RECT 3.955 86.075 4.275 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 85.665 4.275 85.985 ;
      LAYER met4 ;
        RECT 3.955 85.665 4.275 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 85.255 4.275 85.575 ;
      LAYER met4 ;
        RECT 3.955 85.255 4.275 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 84.845 4.275 85.165 ;
      LAYER met4 ;
        RECT 3.955 84.845 4.275 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 84.435 4.275 84.755 ;
      LAYER met4 ;
        RECT 3.955 84.435 4.275 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 84.025 4.275 84.345 ;
      LAYER met4 ;
        RECT 3.955 84.025 4.275 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 83.615 4.275 83.935 ;
      LAYER met4 ;
        RECT 3.955 83.615 4.275 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 83.205 4.275 83.525 ;
      LAYER met4 ;
        RECT 3.955 83.205 4.275 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.955 82.795 4.275 83.115 ;
      LAYER met4 ;
        RECT 3.955 82.795 4.275 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 22.160 4.130 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 21.730 4.130 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 21.300 4.130 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 20.870 4.130 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 20.440 4.130 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 20.010 4.130 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 19.580 4.130 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 19.150 4.130 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 18.720 4.130 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 18.290 4.130 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.930 17.860 4.130 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 82.300 3.905 82.620 ;
      LAYER met4 ;
        RECT 3.585 82.300 3.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 81.895 3.905 82.215 ;
      LAYER met4 ;
        RECT 3.585 81.895 3.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 81.490 3.905 81.810 ;
      LAYER met4 ;
        RECT 3.585 81.490 3.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 81.085 3.905 81.405 ;
      LAYER met4 ;
        RECT 3.585 81.085 3.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 80.680 3.905 81.000 ;
      LAYER met4 ;
        RECT 3.585 80.680 3.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 80.275 3.905 80.595 ;
      LAYER met4 ;
        RECT 3.585 80.275 3.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 79.870 3.905 80.190 ;
      LAYER met4 ;
        RECT 3.585 79.870 3.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 79.465 3.905 79.785 ;
      LAYER met4 ;
        RECT 3.585 79.465 3.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 79.060 3.905 79.380 ;
      LAYER met4 ;
        RECT 3.585 79.060 3.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 78.655 3.905 78.975 ;
      LAYER met4 ;
        RECT 3.585 78.655 3.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 78.250 3.905 78.570 ;
      LAYER met4 ;
        RECT 3.585 78.250 3.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 77.845 3.905 78.165 ;
      LAYER met4 ;
        RECT 3.585 77.845 3.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 77.440 3.905 77.760 ;
      LAYER met4 ;
        RECT 3.585 77.440 3.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 77.035 3.905 77.355 ;
      LAYER met4 ;
        RECT 3.585 77.035 3.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 76.630 3.905 76.950 ;
      LAYER met4 ;
        RECT 3.585 76.630 3.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 76.225 3.905 76.545 ;
      LAYER met4 ;
        RECT 3.585 76.225 3.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 75.820 3.905 76.140 ;
      LAYER met4 ;
        RECT 3.585 75.820 3.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 75.415 3.905 75.735 ;
      LAYER met4 ;
        RECT 3.585 75.415 3.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 75.010 3.905 75.330 ;
      LAYER met4 ;
        RECT 3.585 75.010 3.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 74.605 3.905 74.925 ;
      LAYER met4 ;
        RECT 3.585 74.605 3.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 74.200 3.905 74.520 ;
      LAYER met4 ;
        RECT 3.585 74.200 3.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 73.795 3.905 74.115 ;
      LAYER met4 ;
        RECT 3.585 73.795 3.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 73.390 3.905 73.710 ;
      LAYER met4 ;
        RECT 3.585 73.390 3.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 72.985 3.905 73.305 ;
      LAYER met4 ;
        RECT 3.585 72.985 3.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 72.575 3.905 72.895 ;
      LAYER met4 ;
        RECT 3.585 72.575 3.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 72.165 3.905 72.485 ;
      LAYER met4 ;
        RECT 3.585 72.165 3.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 71.755 3.905 72.075 ;
      LAYER met4 ;
        RECT 3.585 71.755 3.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 71.345 3.905 71.665 ;
      LAYER met4 ;
        RECT 3.585 71.345 3.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 70.935 3.905 71.255 ;
      LAYER met4 ;
        RECT 3.585 70.935 3.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 70.525 3.905 70.845 ;
      LAYER met4 ;
        RECT 3.585 70.525 3.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 70.115 3.905 70.435 ;
      LAYER met4 ;
        RECT 3.585 70.115 3.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 69.705 3.905 70.025 ;
      LAYER met4 ;
        RECT 3.585 69.705 3.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 69.295 3.905 69.615 ;
      LAYER met4 ;
        RECT 3.585 69.295 3.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 68.885 3.905 69.205 ;
      LAYER met4 ;
        RECT 3.585 68.885 3.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 68.475 3.905 68.795 ;
      LAYER met4 ;
        RECT 3.585 68.475 3.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.585 68.065 3.905 68.385 ;
      LAYER met4 ;
        RECT 3.585 68.065 3.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 92.635 3.865 92.955 ;
      LAYER met4 ;
        RECT 3.545 92.635 3.865 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 92.225 3.865 92.545 ;
      LAYER met4 ;
        RECT 3.545 92.225 3.865 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 91.815 3.865 92.135 ;
      LAYER met4 ;
        RECT 3.545 91.815 3.865 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 91.405 3.865 91.725 ;
      LAYER met4 ;
        RECT 3.545 91.405 3.865 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 90.995 3.865 91.315 ;
      LAYER met4 ;
        RECT 3.545 90.995 3.865 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 90.585 3.865 90.905 ;
      LAYER met4 ;
        RECT 3.545 90.585 3.865 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 90.175 3.865 90.495 ;
      LAYER met4 ;
        RECT 3.545 90.175 3.865 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 89.765 3.865 90.085 ;
      LAYER met4 ;
        RECT 3.545 89.765 3.865 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 89.355 3.865 89.675 ;
      LAYER met4 ;
        RECT 3.545 89.355 3.865 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 88.945 3.865 89.265 ;
      LAYER met4 ;
        RECT 3.545 88.945 3.865 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 88.535 3.865 88.855 ;
      LAYER met4 ;
        RECT 3.545 88.535 3.865 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 88.125 3.865 88.445 ;
      LAYER met4 ;
        RECT 3.545 88.125 3.865 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 87.715 3.865 88.035 ;
      LAYER met4 ;
        RECT 3.545 87.715 3.865 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 87.305 3.865 87.625 ;
      LAYER met4 ;
        RECT 3.545 87.305 3.865 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 86.895 3.865 87.215 ;
      LAYER met4 ;
        RECT 3.545 86.895 3.865 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 86.485 3.865 86.805 ;
      LAYER met4 ;
        RECT 3.545 86.485 3.865 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 86.075 3.865 86.395 ;
      LAYER met4 ;
        RECT 3.545 86.075 3.865 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 85.665 3.865 85.985 ;
      LAYER met4 ;
        RECT 3.545 85.665 3.865 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 85.255 3.865 85.575 ;
      LAYER met4 ;
        RECT 3.545 85.255 3.865 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 84.845 3.865 85.165 ;
      LAYER met4 ;
        RECT 3.545 84.845 3.865 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 84.435 3.865 84.755 ;
      LAYER met4 ;
        RECT 3.545 84.435 3.865 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 84.025 3.865 84.345 ;
      LAYER met4 ;
        RECT 3.545 84.025 3.865 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 83.615 3.865 83.935 ;
      LAYER met4 ;
        RECT 3.545 83.615 3.865 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 83.205 3.865 83.525 ;
      LAYER met4 ;
        RECT 3.545 83.205 3.865 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.545 82.795 3.865 83.115 ;
      LAYER met4 ;
        RECT 3.545 82.795 3.865 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 22.160 3.725 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 21.730 3.725 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 21.300 3.725 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 20.870 3.725 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 20.440 3.725 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 20.010 3.725 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 19.580 3.725 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 19.150 3.725 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 18.720 3.725 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 18.290 3.725 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.525 17.860 3.725 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 82.300 3.505 82.620 ;
      LAYER met4 ;
        RECT 3.185 82.300 3.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 81.895 3.505 82.215 ;
      LAYER met4 ;
        RECT 3.185 81.895 3.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 81.490 3.505 81.810 ;
      LAYER met4 ;
        RECT 3.185 81.490 3.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 81.085 3.505 81.405 ;
      LAYER met4 ;
        RECT 3.185 81.085 3.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 80.680 3.505 81.000 ;
      LAYER met4 ;
        RECT 3.185 80.680 3.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 80.275 3.505 80.595 ;
      LAYER met4 ;
        RECT 3.185 80.275 3.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 79.870 3.505 80.190 ;
      LAYER met4 ;
        RECT 3.185 79.870 3.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 79.465 3.505 79.785 ;
      LAYER met4 ;
        RECT 3.185 79.465 3.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 79.060 3.505 79.380 ;
      LAYER met4 ;
        RECT 3.185 79.060 3.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 78.655 3.505 78.975 ;
      LAYER met4 ;
        RECT 3.185 78.655 3.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 78.250 3.505 78.570 ;
      LAYER met4 ;
        RECT 3.185 78.250 3.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 77.845 3.505 78.165 ;
      LAYER met4 ;
        RECT 3.185 77.845 3.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 77.440 3.505 77.760 ;
      LAYER met4 ;
        RECT 3.185 77.440 3.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 77.035 3.505 77.355 ;
      LAYER met4 ;
        RECT 3.185 77.035 3.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 76.630 3.505 76.950 ;
      LAYER met4 ;
        RECT 3.185 76.630 3.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 76.225 3.505 76.545 ;
      LAYER met4 ;
        RECT 3.185 76.225 3.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 75.820 3.505 76.140 ;
      LAYER met4 ;
        RECT 3.185 75.820 3.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 75.415 3.505 75.735 ;
      LAYER met4 ;
        RECT 3.185 75.415 3.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 75.010 3.505 75.330 ;
      LAYER met4 ;
        RECT 3.185 75.010 3.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 74.605 3.505 74.925 ;
      LAYER met4 ;
        RECT 3.185 74.605 3.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 74.200 3.505 74.520 ;
      LAYER met4 ;
        RECT 3.185 74.200 3.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 73.795 3.505 74.115 ;
      LAYER met4 ;
        RECT 3.185 73.795 3.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 73.390 3.505 73.710 ;
      LAYER met4 ;
        RECT 3.185 73.390 3.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 72.985 3.505 73.305 ;
      LAYER met4 ;
        RECT 3.185 72.985 3.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 72.575 3.505 72.895 ;
      LAYER met4 ;
        RECT 3.185 72.575 3.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 72.165 3.505 72.485 ;
      LAYER met4 ;
        RECT 3.185 72.165 3.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 71.755 3.505 72.075 ;
      LAYER met4 ;
        RECT 3.185 71.755 3.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 71.345 3.505 71.665 ;
      LAYER met4 ;
        RECT 3.185 71.345 3.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 70.935 3.505 71.255 ;
      LAYER met4 ;
        RECT 3.185 70.935 3.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 70.525 3.505 70.845 ;
      LAYER met4 ;
        RECT 3.185 70.525 3.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 70.115 3.505 70.435 ;
      LAYER met4 ;
        RECT 3.185 70.115 3.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 69.705 3.505 70.025 ;
      LAYER met4 ;
        RECT 3.185 69.705 3.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 69.295 3.505 69.615 ;
      LAYER met4 ;
        RECT 3.185 69.295 3.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 68.885 3.505 69.205 ;
      LAYER met4 ;
        RECT 3.185 68.885 3.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 68.475 3.505 68.795 ;
      LAYER met4 ;
        RECT 3.185 68.475 3.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.185 68.065 3.505 68.385 ;
      LAYER met4 ;
        RECT 3.185 68.065 3.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 92.635 3.455 92.955 ;
      LAYER met4 ;
        RECT 3.135 92.635 3.455 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 92.225 3.455 92.545 ;
      LAYER met4 ;
        RECT 3.135 92.225 3.455 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 91.815 3.455 92.135 ;
      LAYER met4 ;
        RECT 3.135 91.815 3.455 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 91.405 3.455 91.725 ;
      LAYER met4 ;
        RECT 3.135 91.405 3.455 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 90.995 3.455 91.315 ;
      LAYER met4 ;
        RECT 3.135 90.995 3.455 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 90.585 3.455 90.905 ;
      LAYER met4 ;
        RECT 3.135 90.585 3.455 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 90.175 3.455 90.495 ;
      LAYER met4 ;
        RECT 3.135 90.175 3.455 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 89.765 3.455 90.085 ;
      LAYER met4 ;
        RECT 3.135 89.765 3.455 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 89.355 3.455 89.675 ;
      LAYER met4 ;
        RECT 3.135 89.355 3.455 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 88.945 3.455 89.265 ;
      LAYER met4 ;
        RECT 3.135 88.945 3.455 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 88.535 3.455 88.855 ;
      LAYER met4 ;
        RECT 3.135 88.535 3.455 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 88.125 3.455 88.445 ;
      LAYER met4 ;
        RECT 3.135 88.125 3.455 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 87.715 3.455 88.035 ;
      LAYER met4 ;
        RECT 3.135 87.715 3.455 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 87.305 3.455 87.625 ;
      LAYER met4 ;
        RECT 3.135 87.305 3.455 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 86.895 3.455 87.215 ;
      LAYER met4 ;
        RECT 3.135 86.895 3.455 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 86.485 3.455 86.805 ;
      LAYER met4 ;
        RECT 3.135 86.485 3.455 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 86.075 3.455 86.395 ;
      LAYER met4 ;
        RECT 3.135 86.075 3.455 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 85.665 3.455 85.985 ;
      LAYER met4 ;
        RECT 3.135 85.665 3.455 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 85.255 3.455 85.575 ;
      LAYER met4 ;
        RECT 3.135 85.255 3.455 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 84.845 3.455 85.165 ;
      LAYER met4 ;
        RECT 3.135 84.845 3.455 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 84.435 3.455 84.755 ;
      LAYER met4 ;
        RECT 3.135 84.435 3.455 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 84.025 3.455 84.345 ;
      LAYER met4 ;
        RECT 3.135 84.025 3.455 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 83.615 3.455 83.935 ;
      LAYER met4 ;
        RECT 3.135 83.615 3.455 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 83.205 3.455 83.525 ;
      LAYER met4 ;
        RECT 3.135 83.205 3.455 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.135 82.795 3.455 83.115 ;
      LAYER met4 ;
        RECT 3.135 82.795 3.455 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 22.160 3.320 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 21.730 3.320 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 21.300 3.320 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 20.870 3.320 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 20.440 3.320 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 20.010 3.320 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 19.580 3.320 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 19.150 3.320 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 18.720 3.320 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 18.290 3.320 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.120 17.860 3.320 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 82.300 3.105 82.620 ;
      LAYER met4 ;
        RECT 2.785 82.300 3.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 81.895 3.105 82.215 ;
      LAYER met4 ;
        RECT 2.785 81.895 3.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 81.490 3.105 81.810 ;
      LAYER met4 ;
        RECT 2.785 81.490 3.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 81.085 3.105 81.405 ;
      LAYER met4 ;
        RECT 2.785 81.085 3.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 80.680 3.105 81.000 ;
      LAYER met4 ;
        RECT 2.785 80.680 3.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 80.275 3.105 80.595 ;
      LAYER met4 ;
        RECT 2.785 80.275 3.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 79.870 3.105 80.190 ;
      LAYER met4 ;
        RECT 2.785 79.870 3.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 79.465 3.105 79.785 ;
      LAYER met4 ;
        RECT 2.785 79.465 3.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 79.060 3.105 79.380 ;
      LAYER met4 ;
        RECT 2.785 79.060 3.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 78.655 3.105 78.975 ;
      LAYER met4 ;
        RECT 2.785 78.655 3.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 78.250 3.105 78.570 ;
      LAYER met4 ;
        RECT 2.785 78.250 3.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 77.845 3.105 78.165 ;
      LAYER met4 ;
        RECT 2.785 77.845 3.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 77.440 3.105 77.760 ;
      LAYER met4 ;
        RECT 2.785 77.440 3.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 77.035 3.105 77.355 ;
      LAYER met4 ;
        RECT 2.785 77.035 3.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 76.630 3.105 76.950 ;
      LAYER met4 ;
        RECT 2.785 76.630 3.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 76.225 3.105 76.545 ;
      LAYER met4 ;
        RECT 2.785 76.225 3.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 75.820 3.105 76.140 ;
      LAYER met4 ;
        RECT 2.785 75.820 3.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 75.415 3.105 75.735 ;
      LAYER met4 ;
        RECT 2.785 75.415 3.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 75.010 3.105 75.330 ;
      LAYER met4 ;
        RECT 2.785 75.010 3.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 74.605 3.105 74.925 ;
      LAYER met4 ;
        RECT 2.785 74.605 3.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 74.200 3.105 74.520 ;
      LAYER met4 ;
        RECT 2.785 74.200 3.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 73.795 3.105 74.115 ;
      LAYER met4 ;
        RECT 2.785 73.795 3.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 73.390 3.105 73.710 ;
      LAYER met4 ;
        RECT 2.785 73.390 3.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 72.985 3.105 73.305 ;
      LAYER met4 ;
        RECT 2.785 72.985 3.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 72.575 3.105 72.895 ;
      LAYER met4 ;
        RECT 2.785 72.575 3.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 72.165 3.105 72.485 ;
      LAYER met4 ;
        RECT 2.785 72.165 3.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 71.755 3.105 72.075 ;
      LAYER met4 ;
        RECT 2.785 71.755 3.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 71.345 3.105 71.665 ;
      LAYER met4 ;
        RECT 2.785 71.345 3.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 70.935 3.105 71.255 ;
      LAYER met4 ;
        RECT 2.785 70.935 3.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 70.525 3.105 70.845 ;
      LAYER met4 ;
        RECT 2.785 70.525 3.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 70.115 3.105 70.435 ;
      LAYER met4 ;
        RECT 2.785 70.115 3.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 69.705 3.105 70.025 ;
      LAYER met4 ;
        RECT 2.785 69.705 3.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 69.295 3.105 69.615 ;
      LAYER met4 ;
        RECT 2.785 69.295 3.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 68.885 3.105 69.205 ;
      LAYER met4 ;
        RECT 2.785 68.885 3.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 68.475 3.105 68.795 ;
      LAYER met4 ;
        RECT 2.785 68.475 3.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.785 68.065 3.105 68.385 ;
      LAYER met4 ;
        RECT 2.785 68.065 3.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 92.635 3.045 92.955 ;
      LAYER met4 ;
        RECT 2.725 92.635 3.045 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 92.225 3.045 92.545 ;
      LAYER met4 ;
        RECT 2.725 92.225 3.045 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 91.815 3.045 92.135 ;
      LAYER met4 ;
        RECT 2.725 91.815 3.045 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 91.405 3.045 91.725 ;
      LAYER met4 ;
        RECT 2.725 91.405 3.045 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 90.995 3.045 91.315 ;
      LAYER met4 ;
        RECT 2.725 90.995 3.045 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 90.585 3.045 90.905 ;
      LAYER met4 ;
        RECT 2.725 90.585 3.045 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 90.175 3.045 90.495 ;
      LAYER met4 ;
        RECT 2.725 90.175 3.045 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 89.765 3.045 90.085 ;
      LAYER met4 ;
        RECT 2.725 89.765 3.045 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 89.355 3.045 89.675 ;
      LAYER met4 ;
        RECT 2.725 89.355 3.045 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 88.945 3.045 89.265 ;
      LAYER met4 ;
        RECT 2.725 88.945 3.045 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 88.535 3.045 88.855 ;
      LAYER met4 ;
        RECT 2.725 88.535 3.045 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 88.125 3.045 88.445 ;
      LAYER met4 ;
        RECT 2.725 88.125 3.045 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 87.715 3.045 88.035 ;
      LAYER met4 ;
        RECT 2.725 87.715 3.045 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 87.305 3.045 87.625 ;
      LAYER met4 ;
        RECT 2.725 87.305 3.045 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 86.895 3.045 87.215 ;
      LAYER met4 ;
        RECT 2.725 86.895 3.045 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 86.485 3.045 86.805 ;
      LAYER met4 ;
        RECT 2.725 86.485 3.045 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 86.075 3.045 86.395 ;
      LAYER met4 ;
        RECT 2.725 86.075 3.045 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 85.665 3.045 85.985 ;
      LAYER met4 ;
        RECT 2.725 85.665 3.045 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 85.255 3.045 85.575 ;
      LAYER met4 ;
        RECT 2.725 85.255 3.045 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 84.845 3.045 85.165 ;
      LAYER met4 ;
        RECT 2.725 84.845 3.045 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 84.435 3.045 84.755 ;
      LAYER met4 ;
        RECT 2.725 84.435 3.045 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 84.025 3.045 84.345 ;
      LAYER met4 ;
        RECT 2.725 84.025 3.045 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 83.615 3.045 83.935 ;
      LAYER met4 ;
        RECT 2.725 83.615 3.045 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 83.205 3.045 83.525 ;
      LAYER met4 ;
        RECT 2.725 83.205 3.045 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.725 82.795 3.045 83.115 ;
      LAYER met4 ;
        RECT 2.725 82.795 3.045 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 22.160 2.915 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 21.730 2.915 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 21.300 2.915 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 20.870 2.915 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 20.440 2.915 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 20.010 2.915 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 19.580 2.915 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 19.150 2.915 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 18.720 2.915 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 18.290 2.915 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.715 17.860 2.915 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 82.300 2.705 82.620 ;
      LAYER met4 ;
        RECT 2.385 82.300 2.705 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 81.895 2.705 82.215 ;
      LAYER met4 ;
        RECT 2.385 81.895 2.705 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 81.490 2.705 81.810 ;
      LAYER met4 ;
        RECT 2.385 81.490 2.705 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 81.085 2.705 81.405 ;
      LAYER met4 ;
        RECT 2.385 81.085 2.705 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 80.680 2.705 81.000 ;
      LAYER met4 ;
        RECT 2.385 80.680 2.705 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 80.275 2.705 80.595 ;
      LAYER met4 ;
        RECT 2.385 80.275 2.705 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 79.870 2.705 80.190 ;
      LAYER met4 ;
        RECT 2.385 79.870 2.705 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 79.465 2.705 79.785 ;
      LAYER met4 ;
        RECT 2.385 79.465 2.705 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 79.060 2.705 79.380 ;
      LAYER met4 ;
        RECT 2.385 79.060 2.705 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 78.655 2.705 78.975 ;
      LAYER met4 ;
        RECT 2.385 78.655 2.705 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 78.250 2.705 78.570 ;
      LAYER met4 ;
        RECT 2.385 78.250 2.705 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 77.845 2.705 78.165 ;
      LAYER met4 ;
        RECT 2.385 77.845 2.705 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 77.440 2.705 77.760 ;
      LAYER met4 ;
        RECT 2.385 77.440 2.705 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 77.035 2.705 77.355 ;
      LAYER met4 ;
        RECT 2.385 77.035 2.705 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 76.630 2.705 76.950 ;
      LAYER met4 ;
        RECT 2.385 76.630 2.705 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 76.225 2.705 76.545 ;
      LAYER met4 ;
        RECT 2.385 76.225 2.705 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 75.820 2.705 76.140 ;
      LAYER met4 ;
        RECT 2.385 75.820 2.705 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 75.415 2.705 75.735 ;
      LAYER met4 ;
        RECT 2.385 75.415 2.705 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 75.010 2.705 75.330 ;
      LAYER met4 ;
        RECT 2.385 75.010 2.705 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 74.605 2.705 74.925 ;
      LAYER met4 ;
        RECT 2.385 74.605 2.705 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 74.200 2.705 74.520 ;
      LAYER met4 ;
        RECT 2.385 74.200 2.705 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 73.795 2.705 74.115 ;
      LAYER met4 ;
        RECT 2.385 73.795 2.705 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 73.390 2.705 73.710 ;
      LAYER met4 ;
        RECT 2.385 73.390 2.705 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 72.985 2.705 73.305 ;
      LAYER met4 ;
        RECT 2.385 72.985 2.705 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 72.575 2.705 72.895 ;
      LAYER met4 ;
        RECT 2.385 72.575 2.705 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 72.165 2.705 72.485 ;
      LAYER met4 ;
        RECT 2.385 72.165 2.705 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 71.755 2.705 72.075 ;
      LAYER met4 ;
        RECT 2.385 71.755 2.705 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 71.345 2.705 71.665 ;
      LAYER met4 ;
        RECT 2.385 71.345 2.705 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 70.935 2.705 71.255 ;
      LAYER met4 ;
        RECT 2.385 70.935 2.705 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 70.525 2.705 70.845 ;
      LAYER met4 ;
        RECT 2.385 70.525 2.705 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 70.115 2.705 70.435 ;
      LAYER met4 ;
        RECT 2.385 70.115 2.705 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 69.705 2.705 70.025 ;
      LAYER met4 ;
        RECT 2.385 69.705 2.705 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 69.295 2.705 69.615 ;
      LAYER met4 ;
        RECT 2.385 69.295 2.705 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 68.885 2.705 69.205 ;
      LAYER met4 ;
        RECT 2.385 68.885 2.705 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 68.475 2.705 68.795 ;
      LAYER met4 ;
        RECT 2.385 68.475 2.705 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.385 68.065 2.705 68.385 ;
      LAYER met4 ;
        RECT 2.385 68.065 2.705 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 92.635 2.635 92.955 ;
      LAYER met4 ;
        RECT 2.315 92.635 2.635 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 92.225 2.635 92.545 ;
      LAYER met4 ;
        RECT 2.315 92.225 2.635 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 91.815 2.635 92.135 ;
      LAYER met4 ;
        RECT 2.315 91.815 2.635 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 91.405 2.635 91.725 ;
      LAYER met4 ;
        RECT 2.315 91.405 2.635 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 90.995 2.635 91.315 ;
      LAYER met4 ;
        RECT 2.315 90.995 2.635 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 90.585 2.635 90.905 ;
      LAYER met4 ;
        RECT 2.315 90.585 2.635 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 90.175 2.635 90.495 ;
      LAYER met4 ;
        RECT 2.315 90.175 2.635 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 89.765 2.635 90.085 ;
      LAYER met4 ;
        RECT 2.315 89.765 2.635 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 89.355 2.635 89.675 ;
      LAYER met4 ;
        RECT 2.315 89.355 2.635 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 88.945 2.635 89.265 ;
      LAYER met4 ;
        RECT 2.315 88.945 2.635 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 88.535 2.635 88.855 ;
      LAYER met4 ;
        RECT 2.315 88.535 2.635 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 88.125 2.635 88.445 ;
      LAYER met4 ;
        RECT 2.315 88.125 2.635 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 87.715 2.635 88.035 ;
      LAYER met4 ;
        RECT 2.315 87.715 2.635 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 87.305 2.635 87.625 ;
      LAYER met4 ;
        RECT 2.315 87.305 2.635 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 86.895 2.635 87.215 ;
      LAYER met4 ;
        RECT 2.315 86.895 2.635 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 86.485 2.635 86.805 ;
      LAYER met4 ;
        RECT 2.315 86.485 2.635 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 86.075 2.635 86.395 ;
      LAYER met4 ;
        RECT 2.315 86.075 2.635 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 85.665 2.635 85.985 ;
      LAYER met4 ;
        RECT 2.315 85.665 2.635 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 85.255 2.635 85.575 ;
      LAYER met4 ;
        RECT 2.315 85.255 2.635 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 84.845 2.635 85.165 ;
      LAYER met4 ;
        RECT 2.315 84.845 2.635 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 84.435 2.635 84.755 ;
      LAYER met4 ;
        RECT 2.315 84.435 2.635 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 84.025 2.635 84.345 ;
      LAYER met4 ;
        RECT 2.315 84.025 2.635 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 83.615 2.635 83.935 ;
      LAYER met4 ;
        RECT 2.315 83.615 2.635 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 83.205 2.635 83.525 ;
      LAYER met4 ;
        RECT 2.315 83.205 2.635 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.315 82.795 2.635 83.115 ;
      LAYER met4 ;
        RECT 2.315 82.795 2.635 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 22.160 2.510 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 21.730 2.510 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 21.300 2.510 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 20.870 2.510 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 20.440 2.510 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 20.010 2.510 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 19.580 2.510 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 19.150 2.510 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 18.720 2.510 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 18.290 2.510 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.310 17.860 2.510 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 82.300 2.305 82.620 ;
      LAYER met4 ;
        RECT 1.985 82.300 2.305 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 81.895 2.305 82.215 ;
      LAYER met4 ;
        RECT 1.985 81.895 2.305 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 81.490 2.305 81.810 ;
      LAYER met4 ;
        RECT 1.985 81.490 2.305 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 81.085 2.305 81.405 ;
      LAYER met4 ;
        RECT 1.985 81.085 2.305 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 80.680 2.305 81.000 ;
      LAYER met4 ;
        RECT 1.985 80.680 2.305 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 80.275 2.305 80.595 ;
      LAYER met4 ;
        RECT 1.985 80.275 2.305 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 79.870 2.305 80.190 ;
      LAYER met4 ;
        RECT 1.985 79.870 2.305 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 79.465 2.305 79.785 ;
      LAYER met4 ;
        RECT 1.985 79.465 2.305 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 79.060 2.305 79.380 ;
      LAYER met4 ;
        RECT 1.985 79.060 2.305 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 78.655 2.305 78.975 ;
      LAYER met4 ;
        RECT 1.985 78.655 2.305 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 78.250 2.305 78.570 ;
      LAYER met4 ;
        RECT 1.985 78.250 2.305 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 77.845 2.305 78.165 ;
      LAYER met4 ;
        RECT 1.985 77.845 2.305 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 77.440 2.305 77.760 ;
      LAYER met4 ;
        RECT 1.985 77.440 2.305 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 77.035 2.305 77.355 ;
      LAYER met4 ;
        RECT 1.985 77.035 2.305 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 76.630 2.305 76.950 ;
      LAYER met4 ;
        RECT 1.985 76.630 2.305 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 76.225 2.305 76.545 ;
      LAYER met4 ;
        RECT 1.985 76.225 2.305 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 75.820 2.305 76.140 ;
      LAYER met4 ;
        RECT 1.985 75.820 2.305 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 75.415 2.305 75.735 ;
      LAYER met4 ;
        RECT 1.985 75.415 2.305 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 75.010 2.305 75.330 ;
      LAYER met4 ;
        RECT 1.985 75.010 2.305 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 74.605 2.305 74.925 ;
      LAYER met4 ;
        RECT 1.985 74.605 2.305 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 74.200 2.305 74.520 ;
      LAYER met4 ;
        RECT 1.985 74.200 2.305 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 73.795 2.305 74.115 ;
      LAYER met4 ;
        RECT 1.985 73.795 2.305 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 73.390 2.305 73.710 ;
      LAYER met4 ;
        RECT 1.985 73.390 2.305 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 72.985 2.305 73.305 ;
      LAYER met4 ;
        RECT 1.985 72.985 2.305 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 72.575 2.305 72.895 ;
      LAYER met4 ;
        RECT 1.985 72.575 2.305 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 72.165 2.305 72.485 ;
      LAYER met4 ;
        RECT 1.985 72.165 2.305 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 71.755 2.305 72.075 ;
      LAYER met4 ;
        RECT 1.985 71.755 2.305 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 71.345 2.305 71.665 ;
      LAYER met4 ;
        RECT 1.985 71.345 2.305 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 70.935 2.305 71.255 ;
      LAYER met4 ;
        RECT 1.985 70.935 2.305 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 70.525 2.305 70.845 ;
      LAYER met4 ;
        RECT 1.985 70.525 2.305 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 70.115 2.305 70.435 ;
      LAYER met4 ;
        RECT 1.985 70.115 2.305 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 69.705 2.305 70.025 ;
      LAYER met4 ;
        RECT 1.985 69.705 2.305 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 69.295 2.305 69.615 ;
      LAYER met4 ;
        RECT 1.985 69.295 2.305 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 68.885 2.305 69.205 ;
      LAYER met4 ;
        RECT 1.985 68.885 2.305 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 68.475 2.305 68.795 ;
      LAYER met4 ;
        RECT 1.985 68.475 2.305 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.985 68.065 2.305 68.385 ;
      LAYER met4 ;
        RECT 1.985 68.065 2.305 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 92.635 2.225 92.955 ;
      LAYER met4 ;
        RECT 1.905 92.635 2.225 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 92.225 2.225 92.545 ;
      LAYER met4 ;
        RECT 1.905 92.225 2.225 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 91.815 2.225 92.135 ;
      LAYER met4 ;
        RECT 1.905 91.815 2.225 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 91.405 2.225 91.725 ;
      LAYER met4 ;
        RECT 1.905 91.405 2.225 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 90.995 2.225 91.315 ;
      LAYER met4 ;
        RECT 1.905 90.995 2.225 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 90.585 2.225 90.905 ;
      LAYER met4 ;
        RECT 1.905 90.585 2.225 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 90.175 2.225 90.495 ;
      LAYER met4 ;
        RECT 1.905 90.175 2.225 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 89.765 2.225 90.085 ;
      LAYER met4 ;
        RECT 1.905 89.765 2.225 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 89.355 2.225 89.675 ;
      LAYER met4 ;
        RECT 1.905 89.355 2.225 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 88.945 2.225 89.265 ;
      LAYER met4 ;
        RECT 1.905 88.945 2.225 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 88.535 2.225 88.855 ;
      LAYER met4 ;
        RECT 1.905 88.535 2.225 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 88.125 2.225 88.445 ;
      LAYER met4 ;
        RECT 1.905 88.125 2.225 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 87.715 2.225 88.035 ;
      LAYER met4 ;
        RECT 1.905 87.715 2.225 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 87.305 2.225 87.625 ;
      LAYER met4 ;
        RECT 1.905 87.305 2.225 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 86.895 2.225 87.215 ;
      LAYER met4 ;
        RECT 1.905 86.895 2.225 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 86.485 2.225 86.805 ;
      LAYER met4 ;
        RECT 1.905 86.485 2.225 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 86.075 2.225 86.395 ;
      LAYER met4 ;
        RECT 1.905 86.075 2.225 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 85.665 2.225 85.985 ;
      LAYER met4 ;
        RECT 1.905 85.665 2.225 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 85.255 2.225 85.575 ;
      LAYER met4 ;
        RECT 1.905 85.255 2.225 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 84.845 2.225 85.165 ;
      LAYER met4 ;
        RECT 1.905 84.845 2.225 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 84.435 2.225 84.755 ;
      LAYER met4 ;
        RECT 1.905 84.435 2.225 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 84.025 2.225 84.345 ;
      LAYER met4 ;
        RECT 1.905 84.025 2.225 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 83.615 2.225 83.935 ;
      LAYER met4 ;
        RECT 1.905 83.615 2.225 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 83.205 2.225 83.525 ;
      LAYER met4 ;
        RECT 1.905 83.205 2.225 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 82.795 2.225 83.115 ;
      LAYER met4 ;
        RECT 1.905 82.795 2.225 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 22.160 2.105 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 21.730 2.105 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 21.300 2.105 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 20.870 2.105 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 20.440 2.105 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 20.010 2.105 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 19.580 2.105 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 19.150 2.105 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 18.720 2.105 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 18.290 2.105 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.905 17.860 2.105 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 82.300 1.905 82.620 ;
      LAYER met4 ;
        RECT 1.585 82.300 1.905 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 81.895 1.905 82.215 ;
      LAYER met4 ;
        RECT 1.585 81.895 1.905 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 81.490 1.905 81.810 ;
      LAYER met4 ;
        RECT 1.585 81.490 1.905 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 81.085 1.905 81.405 ;
      LAYER met4 ;
        RECT 1.585 81.085 1.905 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 80.680 1.905 81.000 ;
      LAYER met4 ;
        RECT 1.585 80.680 1.905 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 80.275 1.905 80.595 ;
      LAYER met4 ;
        RECT 1.585 80.275 1.905 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 79.870 1.905 80.190 ;
      LAYER met4 ;
        RECT 1.585 79.870 1.905 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 79.465 1.905 79.785 ;
      LAYER met4 ;
        RECT 1.585 79.465 1.905 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 79.060 1.905 79.380 ;
      LAYER met4 ;
        RECT 1.585 79.060 1.905 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 78.655 1.905 78.975 ;
      LAYER met4 ;
        RECT 1.585 78.655 1.905 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 78.250 1.905 78.570 ;
      LAYER met4 ;
        RECT 1.585 78.250 1.905 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 77.845 1.905 78.165 ;
      LAYER met4 ;
        RECT 1.585 77.845 1.905 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 77.440 1.905 77.760 ;
      LAYER met4 ;
        RECT 1.585 77.440 1.905 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 77.035 1.905 77.355 ;
      LAYER met4 ;
        RECT 1.585 77.035 1.905 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 76.630 1.905 76.950 ;
      LAYER met4 ;
        RECT 1.585 76.630 1.905 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 76.225 1.905 76.545 ;
      LAYER met4 ;
        RECT 1.585 76.225 1.905 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 75.820 1.905 76.140 ;
      LAYER met4 ;
        RECT 1.585 75.820 1.905 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 75.415 1.905 75.735 ;
      LAYER met4 ;
        RECT 1.585 75.415 1.905 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 75.010 1.905 75.330 ;
      LAYER met4 ;
        RECT 1.585 75.010 1.905 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 74.605 1.905 74.925 ;
      LAYER met4 ;
        RECT 1.585 74.605 1.905 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 74.200 1.905 74.520 ;
      LAYER met4 ;
        RECT 1.585 74.200 1.905 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 73.795 1.905 74.115 ;
      LAYER met4 ;
        RECT 1.585 73.795 1.905 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 73.390 1.905 73.710 ;
      LAYER met4 ;
        RECT 1.585 73.390 1.905 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 72.985 1.905 73.305 ;
      LAYER met4 ;
        RECT 1.585 72.985 1.905 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 72.575 1.905 72.895 ;
      LAYER met4 ;
        RECT 1.585 72.575 1.905 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 72.165 1.905 72.485 ;
      LAYER met4 ;
        RECT 1.585 72.165 1.905 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 71.755 1.905 72.075 ;
      LAYER met4 ;
        RECT 1.585 71.755 1.905 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 71.345 1.905 71.665 ;
      LAYER met4 ;
        RECT 1.585 71.345 1.905 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 70.935 1.905 71.255 ;
      LAYER met4 ;
        RECT 1.585 70.935 1.905 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 70.525 1.905 70.845 ;
      LAYER met4 ;
        RECT 1.585 70.525 1.905 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 70.115 1.905 70.435 ;
      LAYER met4 ;
        RECT 1.585 70.115 1.905 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 69.705 1.905 70.025 ;
      LAYER met4 ;
        RECT 1.585 69.705 1.905 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 69.295 1.905 69.615 ;
      LAYER met4 ;
        RECT 1.585 69.295 1.905 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 68.885 1.905 69.205 ;
      LAYER met4 ;
        RECT 1.585 68.885 1.905 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 68.475 1.905 68.795 ;
      LAYER met4 ;
        RECT 1.585 68.475 1.905 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.585 68.065 1.905 68.385 ;
      LAYER met4 ;
        RECT 1.585 68.065 1.905 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 92.635 1.815 92.955 ;
      LAYER met4 ;
        RECT 1.495 92.635 1.815 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 92.225 1.815 92.545 ;
      LAYER met4 ;
        RECT 1.495 92.225 1.815 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 91.815 1.815 92.135 ;
      LAYER met4 ;
        RECT 1.495 91.815 1.815 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 91.405 1.815 91.725 ;
      LAYER met4 ;
        RECT 1.495 91.405 1.815 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 90.995 1.815 91.315 ;
      LAYER met4 ;
        RECT 1.495 90.995 1.815 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 90.585 1.815 90.905 ;
      LAYER met4 ;
        RECT 1.495 90.585 1.815 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 90.175 1.815 90.495 ;
      LAYER met4 ;
        RECT 1.495 90.175 1.815 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 89.765 1.815 90.085 ;
      LAYER met4 ;
        RECT 1.495 89.765 1.815 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 89.355 1.815 89.675 ;
      LAYER met4 ;
        RECT 1.495 89.355 1.815 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 88.945 1.815 89.265 ;
      LAYER met4 ;
        RECT 1.495 88.945 1.815 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 88.535 1.815 88.855 ;
      LAYER met4 ;
        RECT 1.495 88.535 1.815 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 88.125 1.815 88.445 ;
      LAYER met4 ;
        RECT 1.495 88.125 1.815 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 87.715 1.815 88.035 ;
      LAYER met4 ;
        RECT 1.495 87.715 1.815 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 87.305 1.815 87.625 ;
      LAYER met4 ;
        RECT 1.495 87.305 1.815 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 86.895 1.815 87.215 ;
      LAYER met4 ;
        RECT 1.495 86.895 1.815 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 86.485 1.815 86.805 ;
      LAYER met4 ;
        RECT 1.495 86.485 1.815 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 86.075 1.815 86.395 ;
      LAYER met4 ;
        RECT 1.495 86.075 1.815 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 85.665 1.815 85.985 ;
      LAYER met4 ;
        RECT 1.495 85.665 1.815 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 85.255 1.815 85.575 ;
      LAYER met4 ;
        RECT 1.495 85.255 1.815 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 84.845 1.815 85.165 ;
      LAYER met4 ;
        RECT 1.495 84.845 1.815 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 84.435 1.815 84.755 ;
      LAYER met4 ;
        RECT 1.495 84.435 1.815 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 84.025 1.815 84.345 ;
      LAYER met4 ;
        RECT 1.495 84.025 1.815 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 83.615 1.815 83.935 ;
      LAYER met4 ;
        RECT 1.495 83.615 1.815 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 83.205 1.815 83.525 ;
      LAYER met4 ;
        RECT 1.495 83.205 1.815 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.495 82.795 1.815 83.115 ;
      LAYER met4 ;
        RECT 1.495 82.795 1.815 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 22.160 1.700 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 21.730 1.700 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 21.300 1.700 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 20.870 1.700 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 20.440 1.700 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 20.010 1.700 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 19.580 1.700 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 19.150 1.700 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 18.720 1.700 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 18.290 1.700 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.500 17.860 1.700 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 82.300 1.505 82.620 ;
      LAYER met4 ;
        RECT 1.270 82.300 1.505 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 81.895 1.505 82.215 ;
      LAYER met4 ;
        RECT 1.270 81.895 1.505 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 81.490 1.505 81.810 ;
      LAYER met4 ;
        RECT 1.270 81.490 1.505 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 81.085 1.505 81.405 ;
      LAYER met4 ;
        RECT 1.270 81.085 1.505 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 80.680 1.505 81.000 ;
      LAYER met4 ;
        RECT 1.270 80.680 1.505 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 80.275 1.505 80.595 ;
      LAYER met4 ;
        RECT 1.270 80.275 1.505 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 79.870 1.505 80.190 ;
      LAYER met4 ;
        RECT 1.270 79.870 1.505 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 79.465 1.505 79.785 ;
      LAYER met4 ;
        RECT 1.270 79.465 1.505 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 79.060 1.505 79.380 ;
      LAYER met4 ;
        RECT 1.270 79.060 1.505 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 78.655 1.505 78.975 ;
      LAYER met4 ;
        RECT 1.270 78.655 1.505 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 78.250 1.505 78.570 ;
      LAYER met4 ;
        RECT 1.270 78.250 1.505 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 77.845 1.505 78.165 ;
      LAYER met4 ;
        RECT 1.270 77.845 1.505 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 77.440 1.505 77.760 ;
      LAYER met4 ;
        RECT 1.270 77.440 1.505 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 77.035 1.505 77.355 ;
      LAYER met4 ;
        RECT 1.270 77.035 1.505 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 76.630 1.505 76.950 ;
      LAYER met4 ;
        RECT 1.270 76.630 1.505 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 76.225 1.505 76.545 ;
      LAYER met4 ;
        RECT 1.270 76.225 1.505 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 75.820 1.505 76.140 ;
      LAYER met4 ;
        RECT 1.270 75.820 1.505 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 75.415 1.505 75.735 ;
      LAYER met4 ;
        RECT 1.270 75.415 1.505 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 75.010 1.505 75.330 ;
      LAYER met4 ;
        RECT 1.270 75.010 1.505 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 74.605 1.505 74.925 ;
      LAYER met4 ;
        RECT 1.270 74.605 1.505 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 74.200 1.505 74.520 ;
      LAYER met4 ;
        RECT 1.270 74.200 1.505 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 73.795 1.505 74.115 ;
      LAYER met4 ;
        RECT 1.270 73.795 1.505 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 73.390 1.505 73.710 ;
      LAYER met4 ;
        RECT 1.270 73.390 1.505 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 72.985 1.505 73.305 ;
      LAYER met4 ;
        RECT 1.270 72.985 1.505 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 72.575 1.505 72.895 ;
      LAYER met4 ;
        RECT 1.270 72.575 1.505 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 72.165 1.505 72.485 ;
      LAYER met4 ;
        RECT 1.270 72.165 1.505 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 71.755 1.505 72.075 ;
      LAYER met4 ;
        RECT 1.270 71.755 1.505 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 71.345 1.505 71.665 ;
      LAYER met4 ;
        RECT 1.270 71.345 1.505 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 70.935 1.505 71.255 ;
      LAYER met4 ;
        RECT 1.270 70.935 1.505 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 70.525 1.505 70.845 ;
      LAYER met4 ;
        RECT 1.270 70.525 1.505 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 70.115 1.505 70.435 ;
      LAYER met4 ;
        RECT 1.270 70.115 1.505 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 69.705 1.505 70.025 ;
      LAYER met4 ;
        RECT 1.270 69.705 1.505 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 69.295 1.505 69.615 ;
      LAYER met4 ;
        RECT 1.270 69.295 1.505 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 68.885 1.505 69.205 ;
      LAYER met4 ;
        RECT 1.270 68.885 1.505 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 68.475 1.505 68.795 ;
      LAYER met4 ;
        RECT 1.270 68.475 1.505 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.185 68.065 1.505 68.385 ;
      LAYER met4 ;
        RECT 1.270 68.065 1.505 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 92.635 1.405 92.955 ;
      LAYER met4 ;
        RECT 1.270 92.635 1.405 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 92.225 1.405 92.545 ;
      LAYER met4 ;
        RECT 1.270 92.225 1.405 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 91.815 1.405 92.135 ;
      LAYER met4 ;
        RECT 1.270 91.815 1.405 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 91.405 1.405 91.725 ;
      LAYER met4 ;
        RECT 1.270 91.405 1.405 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 90.995 1.405 91.315 ;
      LAYER met4 ;
        RECT 1.270 90.995 1.405 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 90.585 1.405 90.905 ;
      LAYER met4 ;
        RECT 1.270 90.585 1.405 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 90.175 1.405 90.495 ;
      LAYER met4 ;
        RECT 1.270 90.175 1.405 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 89.765 1.405 90.085 ;
      LAYER met4 ;
        RECT 1.270 89.765 1.405 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 89.355 1.405 89.675 ;
      LAYER met4 ;
        RECT 1.270 89.355 1.405 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 88.945 1.405 89.265 ;
      LAYER met4 ;
        RECT 1.270 88.945 1.405 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 88.535 1.405 88.855 ;
      LAYER met4 ;
        RECT 1.270 88.535 1.405 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 88.125 1.405 88.445 ;
      LAYER met4 ;
        RECT 1.270 88.125 1.405 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 87.715 1.405 88.035 ;
      LAYER met4 ;
        RECT 1.270 87.715 1.405 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 87.305 1.405 87.625 ;
      LAYER met4 ;
        RECT 1.270 87.305 1.405 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 86.895 1.405 87.215 ;
      LAYER met4 ;
        RECT 1.270 86.895 1.405 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 86.485 1.405 86.805 ;
      LAYER met4 ;
        RECT 1.270 86.485 1.405 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 86.075 1.405 86.395 ;
      LAYER met4 ;
        RECT 1.270 86.075 1.405 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 85.665 1.405 85.985 ;
      LAYER met4 ;
        RECT 1.270 85.665 1.405 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 85.255 1.405 85.575 ;
      LAYER met4 ;
        RECT 1.270 85.255 1.405 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 84.845 1.405 85.165 ;
      LAYER met4 ;
        RECT 1.270 84.845 1.405 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 84.435 1.405 84.755 ;
      LAYER met4 ;
        RECT 1.270 84.435 1.405 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 84.025 1.405 84.345 ;
      LAYER met4 ;
        RECT 1.270 84.025 1.405 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 83.615 1.405 83.935 ;
      LAYER met4 ;
        RECT 1.270 83.615 1.405 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 83.205 1.405 83.525 ;
      LAYER met4 ;
        RECT 1.270 83.205 1.405 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.085 82.795 1.405 83.115 ;
      LAYER met4 ;
        RECT 1.270 82.795 1.405 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 22.160 1.295 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 21.730 1.295 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 21.300 1.295 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 20.870 1.295 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 20.440 1.295 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 20.010 1.295 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 19.580 1.295 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 19.150 1.295 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 18.720 1.295 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 18.290 1.295 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.095 17.860 1.295 18.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 82.300 1.105 82.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 81.895 1.105 82.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 81.490 1.105 81.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 81.085 1.105 81.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 80.680 1.105 81.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 80.275 1.105 80.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 79.870 1.105 80.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 79.465 1.105 79.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 79.060 1.105 79.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 78.655 1.105 78.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 78.250 1.105 78.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 77.845 1.105 78.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 77.440 1.105 77.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 77.035 1.105 77.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 76.630 1.105 76.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 76.225 1.105 76.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 75.820 1.105 76.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 75.415 1.105 75.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 75.010 1.105 75.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 74.605 1.105 74.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 74.200 1.105 74.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 73.795 1.105 74.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 73.390 1.105 73.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 72.985 1.105 73.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 72.575 1.105 72.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 72.165 1.105 72.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 71.755 1.105 72.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 71.345 1.105 71.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 70.935 1.105 71.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 70.525 1.105 70.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 70.115 1.105 70.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 69.705 1.105 70.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 69.295 1.105 69.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 68.885 1.105 69.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 68.475 1.105 68.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.785 68.065 1.105 68.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 92.635 0.995 92.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 92.225 0.995 92.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 91.815 0.995 92.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 91.405 0.995 91.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 90.995 0.995 91.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 90.585 0.995 90.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 90.175 0.995 90.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 89.765 0.995 90.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 89.355 0.995 89.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 88.945 0.995 89.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 88.535 0.995 88.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 88.125 0.995 88.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 87.715 0.995 88.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 87.305 0.995 87.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 86.895 0.995 87.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 86.485 0.995 86.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 86.075 0.995 86.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 85.665 0.995 85.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 85.255 0.995 85.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 84.845 0.995 85.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 84.435 0.995 84.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 84.025 0.995 84.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 83.615 0.995 83.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 83.205 0.995 83.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.675 82.795 0.995 83.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 22.160 0.890 22.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 21.730 0.890 21.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 21.300 0.890 21.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 20.870 0.890 21.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 20.440 0.890 20.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 20.010 0.890 20.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 19.580 0.890 19.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 19.150 0.890 19.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 18.720 0.890 18.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 18.290 0.890 18.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.690 17.860 0.890 18.060 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
  END VCCHIB
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
  END VSWITCH
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
  END VSSIO_Q
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
  END VSSIO
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.595 92.135 59.430 92.955 ;
        RECT 0.595 91.245 58.540 92.135 ;
        RECT 61.455 91.335 74.660 92.465 ;
        RECT 0.595 89.955 57.250 91.245 ;
        RECT 60.230 90.445 74.660 91.335 ;
        RECT 0.595 88.565 55.860 89.955 ;
        RECT 59.340 89.155 74.660 90.445 ;
        RECT 0.595 87.440 54.735 88.565 ;
        RECT 58.050 87.765 74.660 89.155 ;
        RECT 0.595 86.015 53.310 87.440 ;
        RECT 56.660 86.640 74.660 87.765 ;
        RECT 0.595 84.710 52.005 86.015 ;
        RECT 55.535 85.215 74.660 86.640 ;
        RECT 0.595 67.635 50.360 84.710 ;
        RECT 54.110 83.910 74.660 85.215 ;
        RECT 52.805 83.065 74.660 83.910 ;
        RECT 0.595 66.930 74.660 67.635 ;
        RECT 0.595 62.090 50.355 66.930 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 92.110 73.330 93.400 ;
        RECT 1.670 90.550 13.855 92.110 ;
        RECT 15.765 91.220 59.490 92.110 ;
        RECT 1.670 87.945 13.870 90.550 ;
        RECT 16.650 89.930 58.605 91.220 ;
        RECT 61.400 90.550 73.330 92.110 ;
        RECT 17.925 88.540 57.330 89.930 ;
        RECT 1.670 82.590 13.975 87.945 ;
        RECT 19.255 87.415 56.000 88.540 ;
        RECT 61.385 87.945 73.330 90.550 ;
        RECT 20.465 85.990 54.790 87.415 ;
        RECT 21.850 84.685 53.405 85.990 ;
        RECT 1.670 82.545 18.770 82.590 ;
        RECT 1.670 82.455 21.250 82.545 ;
        RECT 23.170 82.455 52.085 84.685 ;
        RECT 61.280 82.590 73.330 87.945 ;
        RECT 56.485 82.545 73.330 82.590 ;
        RECT 54.005 82.455 73.330 82.545 ;
        RECT 1.670 67.635 73.330 82.455 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 94.585 75.000 172.185 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__overlay_vddio_lvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vssa_hvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vssa_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
  END VCCD
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
  END VSWITCH
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
  END VCCHIB
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 1.270 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 1.270 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 47.740 24.395 48.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 56.410 24.395 56.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.970 36.740 24.395 40.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 36.740 74.290 40.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 47.740 74.290 48.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 51.650 74.290 52.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 56.410 74.290 56.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 56.470 74.200 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 52.555 74.200 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 52.135 74.200 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 51.715 74.200 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 47.800 74.200 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 39.900 74.200 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 39.460 74.200 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 39.020 74.200 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 38.580 74.200 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 38.140 74.200 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 37.700 74.200 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 37.260 74.200 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 36.820 74.200 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 52.555 73.795 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 52.135 73.795 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 51.715 73.795 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 39.900 73.795 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 39.460 73.795 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 39.020 73.795 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 38.580 73.795 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 38.140 73.795 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 37.700 73.795 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 37.260 73.795 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 36.820 73.795 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590 56.470 73.790 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.590 47.800 73.790 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 52.555 73.390 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 52.135 73.390 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 51.715 73.390 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 39.900 73.390 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 39.460 73.390 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 39.020 73.390 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 38.580 73.390 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 38.140 73.390 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 37.700 73.390 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 37.260 73.390 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 36.820 73.390 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.180 56.470 73.380 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.180 47.800 73.380 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 52.555 72.985 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 52.135 72.985 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 51.715 72.985 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 39.900 72.985 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 39.460 72.985 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 39.020 72.985 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 38.580 72.985 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 38.140 72.985 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 37.700 72.985 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 37.260 72.985 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 36.820 72.985 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.770 56.470 72.970 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.770 47.800 72.970 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 52.555 72.580 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 52.135 72.580 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 51.715 72.580 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 39.900 72.580 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 39.460 72.580 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 39.020 72.580 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 38.580 72.580 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 38.140 72.580 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 37.700 72.580 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 37.260 72.580 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 36.820 72.580 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.360 56.470 72.560 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.360 47.800 72.560 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 52.555 72.175 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 52.135 72.175 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 51.715 72.175 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 39.900 72.175 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 39.460 72.175 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 39.020 72.175 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 38.580 72.175 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 38.140 72.175 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 37.700 72.175 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 37.260 72.175 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 36.820 72.175 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.950 56.470 72.150 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.950 47.800 72.150 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 52.555 71.770 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 52.135 71.770 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 51.715 71.770 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 39.900 71.770 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 39.460 71.770 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 39.020 71.770 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 38.580 71.770 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 38.140 71.770 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 37.700 71.770 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 37.260 71.770 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 36.820 71.770 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.540 56.470 71.740 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.540 47.800 71.740 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 52.555 71.365 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 52.135 71.365 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 51.715 71.365 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 39.900 71.365 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 39.460 71.365 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 39.020 71.365 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 38.580 71.365 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 38.140 71.365 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 37.700 71.365 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 37.260 71.365 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 36.820 71.365 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.135 56.470 71.335 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.135 47.800 71.335 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 52.555 70.960 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 52.135 70.960 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 51.715 70.960 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 39.900 70.960 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 39.460 70.960 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 39.020 70.960 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 38.580 70.960 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 38.140 70.960 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 37.700 70.960 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 37.260 70.960 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 36.820 70.960 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 56.470 70.930 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 47.800 70.930 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 52.555 70.555 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 52.135 70.555 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 51.715 70.555 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 39.900 70.555 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 39.460 70.555 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 39.020 70.555 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 38.580 70.555 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 38.140 70.555 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 37.700 70.555 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 37.260 70.555 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 36.820 70.555 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.325 56.470 70.525 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.325 47.800 70.525 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 52.555 70.150 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 52.135 70.150 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 51.715 70.150 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 39.900 70.150 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 39.460 70.150 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 39.020 70.150 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 38.580 70.150 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 38.140 70.150 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 37.700 70.150 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 37.260 70.150 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 36.820 70.150 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.920 56.470 70.120 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.920 47.800 70.120 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 52.555 69.745 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 52.135 69.745 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 51.715 69.745 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 39.900 69.745 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 39.460 69.745 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 39.020 69.745 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 38.580 69.745 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 38.140 69.745 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 37.700 69.745 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 37.260 69.745 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 36.820 69.745 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.515 56.470 69.715 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.515 47.800 69.715 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 52.555 69.340 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 52.135 69.340 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 51.715 69.340 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 39.900 69.340 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 39.460 69.340 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 39.020 69.340 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 38.580 69.340 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 38.140 69.340 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 37.700 69.340 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 37.260 69.340 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 36.820 69.340 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 56.470 69.310 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 47.800 69.310 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 52.555 68.935 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 52.135 68.935 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 51.715 68.935 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 39.900 68.935 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 39.460 68.935 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 39.020 68.935 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 38.580 68.935 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 38.140 68.935 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 37.700 68.935 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 37.260 68.935 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 36.820 68.935 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.705 56.470 68.905 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.705 47.800 68.905 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 52.555 68.530 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 52.135 68.530 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 51.715 68.530 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 39.900 68.530 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 39.460 68.530 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 39.020 68.530 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 38.580 68.530 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 38.140 68.530 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 37.700 68.530 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 37.260 68.530 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 36.820 68.530 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.300 56.470 68.500 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.300 47.800 68.500 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 52.555 68.125 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 52.135 68.125 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 51.715 68.125 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 39.900 68.125 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 39.460 68.125 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 39.020 68.125 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 38.580 68.125 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 38.140 68.125 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 37.700 68.125 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 37.260 68.125 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 36.820 68.125 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.895 56.470 68.095 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.895 47.800 68.095 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 52.555 67.720 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 52.135 67.720 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 51.715 67.720 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 39.900 67.720 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 39.460 67.720 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 39.020 67.720 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 38.580 67.720 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 38.140 67.720 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 37.700 67.720 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 37.260 67.720 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 36.820 67.720 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.490 56.470 67.690 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.490 47.800 67.690 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 52.555 67.315 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 52.135 67.315 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 51.715 67.315 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 39.900 67.315 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 39.460 67.315 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 39.020 67.315 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 38.580 67.315 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 38.140 67.315 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 37.700 67.315 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 37.260 67.315 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 36.820 67.315 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.085 56.470 67.285 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.085 47.800 67.285 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 52.555 66.910 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 52.135 66.910 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 51.715 66.910 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 39.900 66.910 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 39.460 66.910 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 39.020 66.910 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 38.580 66.910 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 38.140 66.910 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 37.700 66.910 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 37.260 66.910 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 36.820 66.910 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.680 56.470 66.880 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.680 47.800 66.880 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 52.555 66.505 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 52.135 66.505 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 51.715 66.505 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 39.900 66.505 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 39.460 66.505 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 39.020 66.505 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 38.580 66.505 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 38.140 66.505 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 37.700 66.505 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 37.260 66.505 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 36.820 66.505 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.275 56.470 66.475 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.275 47.800 66.475 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 52.555 66.100 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 52.135 66.100 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 51.715 66.100 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 39.900 66.100 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 39.460 66.100 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 39.020 66.100 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 38.580 66.100 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 38.140 66.100 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 37.700 66.100 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 37.260 66.100 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 36.820 66.100 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.870 56.470 66.070 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.870 47.800 66.070 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 52.555 65.695 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 52.135 65.695 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 51.715 65.695 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 39.900 65.695 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 39.460 65.695 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 39.020 65.695 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 38.580 65.695 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 38.140 65.695 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 37.700 65.695 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 37.260 65.695 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 36.820 65.695 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.465 56.470 65.665 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.465 47.800 65.665 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 52.555 65.290 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 52.135 65.290 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 51.715 65.290 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 39.900 65.290 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 39.460 65.290 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 39.020 65.290 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 38.580 65.290 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 38.140 65.290 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 37.700 65.290 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 37.260 65.290 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 36.820 65.290 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.060 56.470 65.260 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.060 47.800 65.260 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 52.555 64.885 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 52.135 64.885 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 51.715 64.885 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 39.900 64.885 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 39.460 64.885 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 39.020 64.885 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 38.580 64.885 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 38.140 64.885 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 37.700 64.885 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 37.260 64.885 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 36.820 64.885 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.655 56.470 64.855 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.655 47.800 64.855 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 52.555 64.480 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 52.135 64.480 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 51.715 64.480 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 39.900 64.480 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 39.460 64.480 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 39.020 64.480 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 38.580 64.480 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 38.140 64.480 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 37.700 64.480 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 37.260 64.480 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 36.820 64.480 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.250 56.470 64.450 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.250 47.800 64.450 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 52.555 64.075 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 52.135 64.075 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 51.715 64.075 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 39.900 64.075 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 39.460 64.075 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 39.020 64.075 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 38.580 64.075 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 38.140 64.075 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 37.700 64.075 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 37.260 64.075 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 36.820 64.075 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.845 56.470 64.045 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.845 47.800 64.045 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 52.555 63.670 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 52.135 63.670 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 51.715 63.670 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 39.900 63.670 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 39.460 63.670 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 39.020 63.670 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 38.580 63.670 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 38.140 63.670 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 37.700 63.670 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 37.260 63.670 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 36.820 63.670 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.440 56.470 63.640 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.440 47.800 63.640 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 52.555 63.265 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 52.135 63.265 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 51.715 63.265 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 39.900 63.265 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 39.460 63.265 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 39.020 63.265 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 38.580 63.265 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 38.140 63.265 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 37.700 63.265 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 37.260 63.265 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 36.820 63.265 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.035 56.470 63.235 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.035 47.800 63.235 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 52.555 62.860 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 52.135 62.860 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 51.715 62.860 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 39.900 62.860 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 39.460 62.860 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 39.020 62.860 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 38.580 62.860 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 38.140 62.860 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 37.700 62.860 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 37.260 62.860 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 36.820 62.860 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.630 56.470 62.830 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.630 47.800 62.830 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 52.555 62.455 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 52.135 62.455 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 51.715 62.455 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 39.900 62.455 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 39.460 62.455 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 39.020 62.455 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 38.580 62.455 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 38.140 62.455 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 37.700 62.455 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 37.260 62.455 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 36.820 62.455 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.225 56.470 62.425 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.225 47.800 62.425 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 52.555 62.050 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 52.135 62.050 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 51.715 62.050 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 39.900 62.050 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 39.460 62.050 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 39.020 62.050 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 38.580 62.050 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 38.140 62.050 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 37.700 62.050 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 37.260 62.050 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 36.820 62.050 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.820 56.470 62.020 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.820 47.800 62.020 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 52.555 61.645 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 52.135 61.645 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 51.715 61.645 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 39.900 61.645 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 39.460 61.645 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 39.020 61.645 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 38.580 61.645 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 38.140 61.645 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 37.700 61.645 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 37.260 61.645 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 36.820 61.645 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.415 56.470 61.615 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.415 47.800 61.615 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 52.555 61.240 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 52.135 61.240 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 51.715 61.240 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 39.900 61.240 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 39.460 61.240 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 39.020 61.240 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 38.580 61.240 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 38.140 61.240 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 37.700 61.240 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 37.260 61.240 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 36.820 61.240 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 56.470 61.210 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.010 47.800 61.210 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 52.555 60.835 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 52.135 60.835 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 51.715 60.835 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 39.900 60.835 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 39.460 60.835 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 39.020 60.835 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 38.580 60.835 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 38.140 60.835 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 37.700 60.835 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 37.260 60.835 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 36.820 60.835 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.605 56.470 60.805 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.605 47.800 60.805 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 52.555 60.430 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 52.135 60.430 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 51.715 60.430 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 39.900 60.430 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 39.460 60.430 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 39.020 60.430 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 38.580 60.430 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 38.140 60.430 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 37.700 60.430 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 37.260 60.430 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 36.820 60.430 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.200 56.470 60.400 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.200 47.800 60.400 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 52.555 60.025 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 52.135 60.025 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 51.715 60.025 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 39.900 60.025 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 39.460 60.025 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 39.020 60.025 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 38.580 60.025 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 38.140 60.025 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 37.700 60.025 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 37.260 60.025 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 36.820 60.025 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.795 56.470 59.995 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.795 47.800 59.995 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 52.555 59.620 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 52.135 59.620 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 51.715 59.620 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 39.900 59.620 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 39.460 59.620 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 39.020 59.620 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 38.580 59.620 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 38.140 59.620 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 37.700 59.620 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 37.260 59.620 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 36.820 59.620 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.390 56.470 59.590 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.390 47.800 59.590 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 52.555 59.215 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 52.135 59.215 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 51.715 59.215 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 39.900 59.215 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 39.460 59.215 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 39.020 59.215 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 38.580 59.215 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 38.140 59.215 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 37.700 59.215 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 37.260 59.215 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 36.820 59.215 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.985 56.470 59.185 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.985 47.800 59.185 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 52.555 58.810 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 52.135 58.810 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 51.715 58.810 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 39.900 58.810 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 39.460 58.810 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 39.020 58.810 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 38.580 58.810 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 38.140 58.810 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 37.700 58.810 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 37.260 58.810 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 36.820 58.810 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.580 56.470 58.780 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.580 47.800 58.780 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 52.555 58.405 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 52.135 58.405 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 51.715 58.405 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 39.900 58.405 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 39.460 58.405 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 39.020 58.405 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 38.580 58.405 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 38.140 58.405 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 37.700 58.405 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 37.260 58.405 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 36.820 58.405 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.175 56.470 58.375 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.175 47.800 58.375 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 52.555 58.000 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 52.135 58.000 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 51.715 58.000 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 39.900 58.000 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 39.460 58.000 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 39.020 58.000 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 38.580 58.000 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 38.140 58.000 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 37.700 58.000 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 37.260 58.000 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 36.820 58.000 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.770 56.470 57.970 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.770 47.800 57.970 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 52.555 57.595 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 52.135 57.595 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 51.715 57.595 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 39.900 57.595 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 39.460 57.595 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 39.020 57.595 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 38.580 57.595 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 38.140 57.595 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 37.700 57.595 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 37.260 57.595 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 36.820 57.595 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.365 56.470 57.565 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.365 47.800 57.565 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 52.555 57.190 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 52.135 57.190 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 51.715 57.190 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 39.900 57.190 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 39.460 57.190 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 39.020 57.190 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 38.580 57.190 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 38.140 57.190 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 37.700 57.190 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 37.260 57.190 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 36.820 57.190 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.960 56.470 57.160 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.960 47.800 57.160 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 52.555 56.785 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 52.135 56.785 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 51.715 56.785 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 39.900 56.785 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 39.460 56.785 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 39.020 56.785 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 38.580 56.785 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 38.140 56.785 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 37.700 56.785 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 37.260 56.785 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 36.820 56.785 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.555 56.470 56.755 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.555 47.800 56.755 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 52.555 56.380 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 52.135 56.380 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 51.715 56.380 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 39.900 56.380 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 39.460 56.380 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 39.020 56.380 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 38.580 56.380 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 38.140 56.380 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 37.700 56.380 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 37.260 56.380 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 36.820 56.380 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150 56.470 56.350 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.150 47.800 56.350 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 52.555 55.975 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 52.135 55.975 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 51.715 55.975 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 39.900 55.975 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 39.460 55.975 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 39.020 55.975 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 38.580 55.975 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 38.140 55.975 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 37.700 55.975 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 37.260 55.975 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 36.820 55.975 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 56.470 55.945 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.745 47.800 55.945 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 52.555 55.570 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 52.135 55.570 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 51.715 55.570 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 39.900 55.570 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 39.460 55.570 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 39.020 55.570 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 38.580 55.570 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 38.140 55.570 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 37.700 55.570 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 37.260 55.570 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 36.820 55.570 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.340 56.470 55.540 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.340 47.800 55.540 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 52.555 55.165 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 52.135 55.165 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 51.715 55.165 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 39.900 55.165 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 39.460 55.165 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 39.020 55.165 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 38.580 55.165 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 38.140 55.165 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 37.700 55.165 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 37.260 55.165 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 36.820 55.165 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.935 56.470 55.135 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.935 47.800 55.135 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 52.555 54.760 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 52.135 54.760 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 51.715 54.760 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 39.900 54.760 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 39.460 54.760 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 39.020 54.760 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 38.580 54.760 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 38.140 54.760 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 37.700 54.760 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 37.260 54.760 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 36.820 54.760 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.530 56.470 54.730 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.530 47.800 54.730 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 52.555 54.355 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 52.135 54.355 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 51.715 54.355 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 39.900 54.355 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 39.460 54.355 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 39.020 54.355 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 38.580 54.355 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 38.140 54.355 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 37.700 54.355 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 37.260 54.355 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 36.820 54.355 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 56.470 54.325 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 47.800 54.325 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 52.555 53.950 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 52.135 53.950 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 51.715 53.950 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 39.900 53.950 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 39.460 53.950 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 39.020 53.950 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 38.580 53.950 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 38.140 53.950 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 37.700 53.950 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 37.260 53.950 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 36.820 53.950 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.720 56.470 53.920 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.720 47.800 53.920 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 52.555 53.545 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 52.135 53.545 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 51.715 53.545 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 39.900 53.545 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 39.460 53.545 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 39.020 53.545 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 38.580 53.545 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 38.140 53.545 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 37.700 53.545 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 37.260 53.545 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 36.820 53.545 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.315 56.470 53.515 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.315 47.800 53.515 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 52.555 53.140 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 52.135 53.140 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 51.715 53.140 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 39.900 53.140 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 39.460 53.140 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 39.020 53.140 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 38.580 53.140 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 38.140 53.140 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 37.700 53.140 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 37.260 53.140 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 36.820 53.140 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.910 56.470 53.110 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.910 47.800 53.110 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 52.555 52.730 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 52.135 52.730 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 51.715 52.730 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 39.900 52.730 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 39.460 52.730 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 39.020 52.730 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 38.580 52.730 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 38.140 52.730 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 37.700 52.730 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 37.260 52.730 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 36.820 52.730 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.505 56.470 52.705 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.505 47.800 52.705 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 52.555 52.320 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 52.135 52.320 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 51.715 52.320 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 39.900 52.320 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 39.460 52.320 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 39.020 52.320 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 38.580 52.320 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 38.140 52.320 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 37.700 52.320 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 37.260 52.320 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 36.820 52.320 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.100 56.470 52.300 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.100 47.800 52.300 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 52.555 51.910 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 52.135 51.910 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 51.715 51.910 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 39.900 51.910 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 39.460 51.910 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 39.020 51.910 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 38.580 51.910 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 38.140 51.910 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 37.700 51.910 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 37.260 51.910 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 36.820 51.910 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.695 56.470 51.895 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.695 47.800 51.895 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 52.555 51.500 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 52.135 51.500 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 51.715 51.500 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 39.900 51.500 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 39.460 51.500 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 39.020 51.500 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 38.580 51.500 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 38.140 51.500 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 37.700 51.500 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 37.260 51.500 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 36.820 51.500 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.290 56.470 51.490 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.290 47.800 51.490 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 52.555 51.090 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 52.135 51.090 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 51.715 51.090 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 39.900 51.090 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 39.460 51.090 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 39.020 51.090 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 38.580 51.090 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 38.140 51.090 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 37.700 51.090 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 37.260 51.090 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 36.820 51.090 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.885 56.470 51.085 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.885 47.800 51.085 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 56.470 50.680 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 52.555 50.680 52.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 52.135 50.680 52.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 51.715 50.680 51.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 47.800 50.680 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 39.900 50.680 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 39.460 50.680 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 39.020 50.680 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 38.580 50.680 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 38.140 50.680 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 37.700 50.680 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 37.260 50.680 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 36.820 50.680 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 56.470 24.305 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 52.495 24.365 52.815 ;
      LAYER met4 ;
        RECT 24.045 52.495 24.365 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 52.075 24.365 52.395 ;
      LAYER met4 ;
        RECT 24.045 52.075 24.365 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 51.655 24.365 51.975 ;
      LAYER met4 ;
        RECT 24.045 51.655 24.365 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 47.800 24.305 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 39.900 24.305 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 39.460 24.305 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 39.020 24.305 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 38.580 24.305 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 38.140 24.305 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 37.700 24.305 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 37.260 24.305 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 36.820 24.305 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 56.470 23.905 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 47.800 23.905 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 39.900 23.905 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 39.460 23.905 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 39.020 23.905 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 38.580 23.905 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 38.140 23.905 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 37.700 23.905 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 37.260 23.905 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 36.820 23.905 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 52.495 23.960 52.815 ;
      LAYER met4 ;
        RECT 23.640 52.495 23.960 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 52.075 23.960 52.395 ;
      LAYER met4 ;
        RECT 23.640 52.075 23.960 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 51.655 23.960 51.975 ;
      LAYER met4 ;
        RECT 23.640 51.655 23.960 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 39.900 23.505 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 39.460 23.505 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 39.020 23.505 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 38.580 23.505 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 38.140 23.505 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 37.700 23.505 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 37.260 23.505 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.305 36.820 23.505 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 56.470 23.500 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 47.800 23.500 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 52.495 23.555 52.815 ;
      LAYER met4 ;
        RECT 23.235 52.495 23.555 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 52.075 23.555 52.395 ;
      LAYER met4 ;
        RECT 23.235 52.075 23.555 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 51.655 23.555 51.975 ;
      LAYER met4 ;
        RECT 23.235 51.655 23.555 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 39.900 23.105 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 39.460 23.105 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 39.020 23.105 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 38.580 23.105 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 38.140 23.105 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 37.700 23.105 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 37.260 23.105 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.905 36.820 23.105 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 56.470 23.095 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 47.800 23.095 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 52.495 23.150 52.815 ;
      LAYER met4 ;
        RECT 22.830 52.495 23.150 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 52.075 23.150 52.395 ;
      LAYER met4 ;
        RECT 22.830 52.075 23.150 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 51.655 23.150 51.975 ;
      LAYER met4 ;
        RECT 22.830 51.655 23.150 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 39.900 22.705 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 39.460 22.705 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 39.020 22.705 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 38.580 22.705 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 38.140 22.705 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 37.700 22.705 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 37.260 22.705 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.505 36.820 22.705 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 56.470 22.690 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 47.800 22.690 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 52.495 22.745 52.815 ;
      LAYER met4 ;
        RECT 22.425 52.495 22.745 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 52.075 22.745 52.395 ;
      LAYER met4 ;
        RECT 22.425 52.075 22.745 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 51.655 22.745 51.975 ;
      LAYER met4 ;
        RECT 22.425 51.655 22.745 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 39.900 22.305 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 39.460 22.305 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 39.020 22.305 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 38.580 22.305 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 38.140 22.305 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 37.700 22.305 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 37.260 22.305 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.105 36.820 22.305 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 56.470 22.285 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 47.800 22.285 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 52.495 22.340 52.815 ;
      LAYER met4 ;
        RECT 22.020 52.495 22.340 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 52.075 22.340 52.395 ;
      LAYER met4 ;
        RECT 22.020 52.075 22.340 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 51.655 22.340 51.975 ;
      LAYER met4 ;
        RECT 22.020 51.655 22.340 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 39.900 21.905 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 39.460 21.905 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 39.020 21.905 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 38.580 21.905 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 38.140 21.905 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 37.700 21.905 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 37.260 21.905 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.705 36.820 21.905 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 56.470 21.880 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 47.800 21.880 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 52.495 21.935 52.815 ;
      LAYER met4 ;
        RECT 21.615 52.495 21.935 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 52.075 21.935 52.395 ;
      LAYER met4 ;
        RECT 21.615 52.075 21.935 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 51.655 21.935 51.975 ;
      LAYER met4 ;
        RECT 21.615 51.655 21.935 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 39.900 21.505 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 39.460 21.505 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 39.020 21.505 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 38.580 21.505 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 38.140 21.505 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 37.700 21.505 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 37.260 21.505 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.305 36.820 21.505 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 56.470 21.475 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 47.800 21.475 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 52.495 21.530 52.815 ;
      LAYER met4 ;
        RECT 21.210 52.495 21.530 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 52.075 21.530 52.395 ;
      LAYER met4 ;
        RECT 21.210 52.075 21.530 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 51.655 21.530 51.975 ;
      LAYER met4 ;
        RECT 21.210 51.655 21.530 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 39.900 21.105 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 39.460 21.105 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 39.020 21.105 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 38.580 21.105 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 38.140 21.105 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 37.700 21.105 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 37.260 21.105 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.905 36.820 21.105 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 56.470 21.070 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 47.800 21.070 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 52.495 21.125 52.815 ;
      LAYER met4 ;
        RECT 20.805 52.495 21.125 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 52.075 21.125 52.395 ;
      LAYER met4 ;
        RECT 20.805 52.075 21.125 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 51.655 21.125 51.975 ;
      LAYER met4 ;
        RECT 20.805 51.655 21.125 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 39.900 20.700 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 39.460 20.700 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 39.020 20.700 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 38.580 20.700 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 38.140 20.700 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 37.700 20.700 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 37.260 20.700 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.500 36.820 20.700 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 56.470 20.665 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 47.800 20.665 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 52.495 20.720 52.815 ;
      LAYER met4 ;
        RECT 20.400 52.495 20.720 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 52.075 20.720 52.395 ;
      LAYER met4 ;
        RECT 20.400 52.075 20.720 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 51.655 20.720 51.975 ;
      LAYER met4 ;
        RECT 20.400 51.655 20.720 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 39.900 20.295 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 39.460 20.295 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 39.020 20.295 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 38.580 20.295 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 38.140 20.295 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 37.700 20.295 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 37.260 20.295 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.095 36.820 20.295 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 56.470 20.260 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 47.800 20.260 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 52.495 20.315 52.815 ;
      LAYER met4 ;
        RECT 19.995 52.495 20.315 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 52.075 20.315 52.395 ;
      LAYER met4 ;
        RECT 19.995 52.075 20.315 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 51.655 20.315 51.975 ;
      LAYER met4 ;
        RECT 19.995 51.655 20.315 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 39.900 19.890 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 39.460 19.890 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 39.020 19.890 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 38.580 19.890 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 38.140 19.890 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 37.700 19.890 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 37.260 19.890 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.690 36.820 19.890 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 56.470 19.855 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 47.800 19.855 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 52.495 19.910 52.815 ;
      LAYER met4 ;
        RECT 19.590 52.495 19.910 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 52.075 19.910 52.395 ;
      LAYER met4 ;
        RECT 19.590 52.075 19.910 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 51.655 19.910 51.975 ;
      LAYER met4 ;
        RECT 19.590 51.655 19.910 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 39.900 19.485 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 39.460 19.485 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 39.020 19.485 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 38.580 19.485 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 38.140 19.485 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 37.700 19.485 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 37.260 19.485 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.285 36.820 19.485 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 56.470 19.450 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 47.800 19.450 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 52.495 19.505 52.815 ;
      LAYER met4 ;
        RECT 19.185 52.495 19.505 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 52.075 19.505 52.395 ;
      LAYER met4 ;
        RECT 19.185 52.075 19.505 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 51.655 19.505 51.975 ;
      LAYER met4 ;
        RECT 19.185 51.655 19.505 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 39.900 19.080 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 39.460 19.080 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 39.020 19.080 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 38.580 19.080 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 38.140 19.080 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 37.700 19.080 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 37.260 19.080 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.880 36.820 19.080 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 56.470 19.045 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 47.800 19.045 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 52.495 19.100 52.815 ;
      LAYER met4 ;
        RECT 18.780 52.495 19.100 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 52.075 19.100 52.395 ;
      LAYER met4 ;
        RECT 18.780 52.075 19.100 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 51.655 19.100 51.975 ;
      LAYER met4 ;
        RECT 18.780 51.655 19.100 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 39.900 18.675 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 39.460 18.675 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 39.020 18.675 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 38.580 18.675 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 38.140 18.675 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 37.700 18.675 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 37.260 18.675 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.475 36.820 18.675 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 56.470 18.640 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 47.800 18.640 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 52.495 18.695 52.815 ;
      LAYER met4 ;
        RECT 18.375 52.495 18.695 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 52.075 18.695 52.395 ;
      LAYER met4 ;
        RECT 18.375 52.075 18.695 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 51.655 18.695 51.975 ;
      LAYER met4 ;
        RECT 18.375 51.655 18.695 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 39.900 18.270 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 39.460 18.270 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 39.020 18.270 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 38.580 18.270 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 38.140 18.270 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 37.700 18.270 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 37.260 18.270 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.070 36.820 18.270 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 56.470 18.235 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 47.800 18.235 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 52.495 18.290 52.815 ;
      LAYER met4 ;
        RECT 17.970 52.495 18.290 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 52.075 18.290 52.395 ;
      LAYER met4 ;
        RECT 17.970 52.075 18.290 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 51.655 18.290 51.975 ;
      LAYER met4 ;
        RECT 17.970 51.655 18.290 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 39.900 17.865 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 39.460 17.865 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 39.020 17.865 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 38.580 17.865 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 38.140 17.865 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 37.700 17.865 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 37.260 17.865 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.665 36.820 17.865 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 56.470 17.830 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 47.800 17.830 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 52.495 17.885 52.815 ;
      LAYER met4 ;
        RECT 17.565 52.495 17.885 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 52.075 17.885 52.395 ;
      LAYER met4 ;
        RECT 17.565 52.075 17.885 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 51.655 17.885 51.975 ;
      LAYER met4 ;
        RECT 17.565 51.655 17.885 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 39.900 17.460 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 39.460 17.460 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 39.020 17.460 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 38.580 17.460 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 38.140 17.460 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 37.700 17.460 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 37.260 17.460 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.260 36.820 17.460 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 56.470 17.425 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 47.800 17.425 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 52.495 17.480 52.815 ;
      LAYER met4 ;
        RECT 17.160 52.495 17.480 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 52.075 17.480 52.395 ;
      LAYER met4 ;
        RECT 17.160 52.075 17.480 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 51.655 17.480 51.975 ;
      LAYER met4 ;
        RECT 17.160 51.655 17.480 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 39.900 17.055 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 39.460 17.055 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 39.020 17.055 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 38.580 17.055 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 38.140 17.055 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 37.700 17.055 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 37.260 17.055 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.855 36.820 17.055 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 56.470 17.020 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 47.800 17.020 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 52.495 17.075 52.815 ;
      LAYER met4 ;
        RECT 16.755 52.495 17.075 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 52.075 17.075 52.395 ;
      LAYER met4 ;
        RECT 16.755 52.075 17.075 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 51.655 17.075 51.975 ;
      LAYER met4 ;
        RECT 16.755 51.655 17.075 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 39.900 16.650 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 39.460 16.650 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 39.020 16.650 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 38.580 16.650 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 38.140 16.650 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 37.700 16.650 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 37.260 16.650 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.450 36.820 16.650 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 56.470 16.615 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 47.800 16.615 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 52.495 16.670 52.815 ;
      LAYER met4 ;
        RECT 16.350 52.495 16.670 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 52.075 16.670 52.395 ;
      LAYER met4 ;
        RECT 16.350 52.075 16.670 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 51.655 16.670 51.975 ;
      LAYER met4 ;
        RECT 16.350 51.655 16.670 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 39.900 16.245 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 39.460 16.245 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 39.020 16.245 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 38.580 16.245 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 38.140 16.245 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 37.700 16.245 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 37.260 16.245 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.045 36.820 16.245 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 56.470 16.210 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 47.800 16.210 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 52.495 16.265 52.815 ;
      LAYER met4 ;
        RECT 15.945 52.495 16.265 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 52.075 16.265 52.395 ;
      LAYER met4 ;
        RECT 15.945 52.075 16.265 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 51.655 16.265 51.975 ;
      LAYER met4 ;
        RECT 15.945 51.655 16.265 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 39.900 15.840 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 39.460 15.840 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 39.020 15.840 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 38.580 15.840 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 38.140 15.840 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 37.700 15.840 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 37.260 15.840 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.640 36.820 15.840 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 56.470 15.805 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 47.800 15.805 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 52.495 15.860 52.815 ;
      LAYER met4 ;
        RECT 15.540 52.495 15.860 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 52.075 15.860 52.395 ;
      LAYER met4 ;
        RECT 15.540 52.075 15.860 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 51.655 15.860 51.975 ;
      LAYER met4 ;
        RECT 15.540 51.655 15.860 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 39.900 15.435 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 39.460 15.435 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 39.020 15.435 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 38.580 15.435 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 38.140 15.435 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 37.700 15.435 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 37.260 15.435 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.235 36.820 15.435 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 56.470 15.400 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 47.800 15.400 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 52.495 15.455 52.815 ;
      LAYER met4 ;
        RECT 15.135 52.495 15.455 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 52.075 15.455 52.395 ;
      LAYER met4 ;
        RECT 15.135 52.075 15.455 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 51.655 15.455 51.975 ;
      LAYER met4 ;
        RECT 15.135 51.655 15.455 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 39.900 15.030 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 39.460 15.030 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 39.020 15.030 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 38.580 15.030 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 38.140 15.030 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 37.700 15.030 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 37.260 15.030 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.830 36.820 15.030 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 56.470 14.995 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 47.800 14.995 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 52.495 15.050 52.815 ;
      LAYER met4 ;
        RECT 14.730 52.495 15.050 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 52.075 15.050 52.395 ;
      LAYER met4 ;
        RECT 14.730 52.075 15.050 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 51.655 15.050 51.975 ;
      LAYER met4 ;
        RECT 14.730 51.655 15.050 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 39.900 14.625 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 39.460 14.625 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 39.020 14.625 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 38.580 14.625 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 38.140 14.625 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 37.700 14.625 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 37.260 14.625 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.425 36.820 14.625 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 56.470 14.590 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 47.800 14.590 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 52.495 14.645 52.815 ;
      LAYER met4 ;
        RECT 14.325 52.495 14.645 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 52.075 14.645 52.395 ;
      LAYER met4 ;
        RECT 14.325 52.075 14.645 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 51.655 14.645 51.975 ;
      LAYER met4 ;
        RECT 14.325 51.655 14.645 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 39.900 14.220 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 39.460 14.220 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 39.020 14.220 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 38.580 14.220 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 38.140 14.220 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 37.700 14.220 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 37.260 14.220 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.020 36.820 14.220 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 56.470 14.185 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 47.800 14.185 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 52.495 14.240 52.815 ;
      LAYER met4 ;
        RECT 13.920 52.495 14.240 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 52.075 14.240 52.395 ;
      LAYER met4 ;
        RECT 13.920 52.075 14.240 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 51.655 14.240 51.975 ;
      LAYER met4 ;
        RECT 13.920 51.655 14.240 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 39.900 13.815 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 39.460 13.815 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 39.020 13.815 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 38.580 13.815 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 38.140 13.815 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 37.700 13.815 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 37.260 13.815 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.615 36.820 13.815 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 56.470 13.780 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 47.800 13.780 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 52.495 13.835 52.815 ;
      LAYER met4 ;
        RECT 13.515 52.495 13.835 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 52.075 13.835 52.395 ;
      LAYER met4 ;
        RECT 13.515 52.075 13.835 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 51.655 13.835 51.975 ;
      LAYER met4 ;
        RECT 13.515 51.655 13.835 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 39.900 13.410 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 39.460 13.410 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 39.020 13.410 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 38.580 13.410 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 38.140 13.410 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 37.700 13.410 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 37.260 13.410 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.210 36.820 13.410 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 56.470 13.375 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 47.800 13.375 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 52.495 13.430 52.815 ;
      LAYER met4 ;
        RECT 13.110 52.495 13.430 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 52.075 13.430 52.395 ;
      LAYER met4 ;
        RECT 13.110 52.075 13.430 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 51.655 13.430 51.975 ;
      LAYER met4 ;
        RECT 13.110 51.655 13.430 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 39.900 13.005 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 39.460 13.005 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 39.020 13.005 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 38.580 13.005 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 38.140 13.005 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 37.700 13.005 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 37.260 13.005 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.805 36.820 13.005 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 56.470 12.970 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 47.800 12.970 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 52.495 13.025 52.815 ;
      LAYER met4 ;
        RECT 12.705 52.495 13.025 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 52.075 13.025 52.395 ;
      LAYER met4 ;
        RECT 12.705 52.075 13.025 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 51.655 13.025 51.975 ;
      LAYER met4 ;
        RECT 12.705 51.655 13.025 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 39.900 12.600 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 39.460 12.600 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 39.020 12.600 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 38.580 12.600 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 38.140 12.600 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 37.700 12.600 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 37.260 12.600 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.400 36.820 12.600 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 56.470 12.565 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 47.800 12.565 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 52.495 12.620 52.815 ;
      LAYER met4 ;
        RECT 12.300 52.495 12.620 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 52.075 12.620 52.395 ;
      LAYER met4 ;
        RECT 12.300 52.075 12.620 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 51.655 12.620 51.975 ;
      LAYER met4 ;
        RECT 12.300 51.655 12.620 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 39.900 12.195 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 39.460 12.195 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 39.020 12.195 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 38.580 12.195 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 38.140 12.195 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 37.700 12.195 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 37.260 12.195 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.995 36.820 12.195 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 56.470 12.160 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 47.800 12.160 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 52.495 12.215 52.815 ;
      LAYER met4 ;
        RECT 11.895 52.495 12.215 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 52.075 12.215 52.395 ;
      LAYER met4 ;
        RECT 11.895 52.075 12.215 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 51.655 12.215 51.975 ;
      LAYER met4 ;
        RECT 11.895 51.655 12.215 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 39.900 11.790 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 39.460 11.790 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 39.020 11.790 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 38.580 11.790 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 38.140 11.790 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 37.700 11.790 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 37.260 11.790 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.590 36.820 11.790 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 56.470 11.755 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 47.800 11.755 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 52.495 11.810 52.815 ;
      LAYER met4 ;
        RECT 11.490 52.495 11.810 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 52.075 11.810 52.395 ;
      LAYER met4 ;
        RECT 11.490 52.075 11.810 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 51.655 11.810 51.975 ;
      LAYER met4 ;
        RECT 11.490 51.655 11.810 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 39.900 11.385 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 39.460 11.385 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 39.020 11.385 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 38.580 11.385 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 38.140 11.385 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 37.700 11.385 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 37.260 11.385 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.185 36.820 11.385 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 56.470 11.350 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 47.800 11.350 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 52.495 11.405 52.815 ;
      LAYER met4 ;
        RECT 11.085 52.495 11.405 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 52.075 11.405 52.395 ;
      LAYER met4 ;
        RECT 11.085 52.075 11.405 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 51.655 11.405 51.975 ;
      LAYER met4 ;
        RECT 11.085 51.655 11.405 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 39.900 10.980 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 39.460 10.980 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 39.020 10.980 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 38.580 10.980 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 38.140 10.980 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 37.700 10.980 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 37.260 10.980 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.780 36.820 10.980 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 56.470 10.945 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 47.800 10.945 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 52.495 11.000 52.815 ;
      LAYER met4 ;
        RECT 10.680 52.495 11.000 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 52.075 11.000 52.395 ;
      LAYER met4 ;
        RECT 10.680 52.075 11.000 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 51.655 11.000 51.975 ;
      LAYER met4 ;
        RECT 10.680 51.655 11.000 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 39.900 10.575 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 39.460 10.575 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 39.020 10.575 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 38.580 10.575 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 38.140 10.575 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 37.700 10.575 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 37.260 10.575 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.375 36.820 10.575 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 56.470 10.540 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 47.800 10.540 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 52.495 10.595 52.815 ;
      LAYER met4 ;
        RECT 10.275 52.495 10.595 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 52.075 10.595 52.395 ;
      LAYER met4 ;
        RECT 10.275 52.075 10.595 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 51.655 10.595 51.975 ;
      LAYER met4 ;
        RECT 10.275 51.655 10.595 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 39.900 10.170 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 39.460 10.170 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 39.020 10.170 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 38.580 10.170 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 38.140 10.170 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 37.700 10.170 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 37.260 10.170 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.970 36.820 10.170 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 56.470 10.135 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 47.800 10.135 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 52.495 10.190 52.815 ;
      LAYER met4 ;
        RECT 9.870 52.495 10.190 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 52.075 10.190 52.395 ;
      LAYER met4 ;
        RECT 9.870 52.075 10.190 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 51.655 10.190 51.975 ;
      LAYER met4 ;
        RECT 9.870 51.655 10.190 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 39.900 9.765 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 39.460 9.765 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 39.020 9.765 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 38.580 9.765 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 38.140 9.765 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 37.700 9.765 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 37.260 9.765 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.565 36.820 9.765 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 56.470 9.730 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 47.800 9.730 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 52.495 9.785 52.815 ;
      LAYER met4 ;
        RECT 9.465 52.495 9.785 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 52.075 9.785 52.395 ;
      LAYER met4 ;
        RECT 9.465 52.075 9.785 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 51.655 9.785 51.975 ;
      LAYER met4 ;
        RECT 9.465 51.655 9.785 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 39.900 9.360 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 39.460 9.360 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 39.020 9.360 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 38.580 9.360 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 38.140 9.360 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 37.700 9.360 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 37.260 9.360 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.160 36.820 9.360 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 56.470 9.325 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 47.800 9.325 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 52.495 9.380 52.815 ;
      LAYER met4 ;
        RECT 9.060 52.495 9.380 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 52.075 9.380 52.395 ;
      LAYER met4 ;
        RECT 9.060 52.075 9.380 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 51.655 9.380 51.975 ;
      LAYER met4 ;
        RECT 9.060 51.655 9.380 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 39.900 8.955 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 39.460 8.955 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 39.020 8.955 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 38.580 8.955 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 38.140 8.955 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 37.700 8.955 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 37.260 8.955 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.755 36.820 8.955 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 56.470 8.920 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 47.800 8.920 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 52.495 8.975 52.815 ;
      LAYER met4 ;
        RECT 8.655 52.495 8.975 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 52.075 8.975 52.395 ;
      LAYER met4 ;
        RECT 8.655 52.075 8.975 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 51.655 8.975 51.975 ;
      LAYER met4 ;
        RECT 8.655 51.655 8.975 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 39.900 8.550 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 39.460 8.550 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 39.020 8.550 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 38.580 8.550 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 38.140 8.550 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 37.700 8.550 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 37.260 8.550 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.350 36.820 8.550 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 56.470 8.515 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 47.800 8.515 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 52.495 8.570 52.815 ;
      LAYER met4 ;
        RECT 8.250 52.495 8.570 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 52.075 8.570 52.395 ;
      LAYER met4 ;
        RECT 8.250 52.075 8.570 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 51.655 8.570 51.975 ;
      LAYER met4 ;
        RECT 8.250 51.655 8.570 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 39.900 8.145 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 39.460 8.145 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 39.020 8.145 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 38.580 8.145 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 38.140 8.145 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 37.700 8.145 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 37.260 8.145 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.945 36.820 8.145 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 56.470 8.110 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 47.800 8.110 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 52.495 8.165 52.815 ;
      LAYER met4 ;
        RECT 7.845 52.495 8.165 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 52.075 8.165 52.395 ;
      LAYER met4 ;
        RECT 7.845 52.075 8.165 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 51.655 8.165 51.975 ;
      LAYER met4 ;
        RECT 7.845 51.655 8.165 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 39.900 7.740 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 39.460 7.740 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 39.020 7.740 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 38.580 7.740 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 38.140 7.740 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 37.700 7.740 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 37.260 7.740 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.540 36.820 7.740 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 56.470 7.705 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 47.800 7.705 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 52.495 7.760 52.815 ;
      LAYER met4 ;
        RECT 7.440 52.495 7.760 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 52.075 7.760 52.395 ;
      LAYER met4 ;
        RECT 7.440 52.075 7.760 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 51.655 7.760 51.975 ;
      LAYER met4 ;
        RECT 7.440 51.655 7.760 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 39.900 7.335 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 39.460 7.335 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 39.020 7.335 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 38.580 7.335 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 38.140 7.335 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 37.700 7.335 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 37.260 7.335 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.135 36.820 7.335 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 56.470 7.300 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 47.800 7.300 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 52.495 7.355 52.815 ;
      LAYER met4 ;
        RECT 7.035 52.495 7.355 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 52.075 7.355 52.395 ;
      LAYER met4 ;
        RECT 7.035 52.075 7.355 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 51.655 7.355 51.975 ;
      LAYER met4 ;
        RECT 7.035 51.655 7.355 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 39.900 6.930 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 39.460 6.930 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 39.020 6.930 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 38.580 6.930 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 38.140 6.930 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 37.700 6.930 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 37.260 6.930 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.730 36.820 6.930 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 56.470 6.895 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 47.800 6.895 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 52.495 6.950 52.815 ;
      LAYER met4 ;
        RECT 6.630 52.495 6.950 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 52.075 6.950 52.395 ;
      LAYER met4 ;
        RECT 6.630 52.075 6.950 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 51.655 6.950 51.975 ;
      LAYER met4 ;
        RECT 6.630 51.655 6.950 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 39.900 6.525 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 39.460 6.525 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 39.020 6.525 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 38.580 6.525 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 38.140 6.525 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 37.700 6.525 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 37.260 6.525 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.325 36.820 6.525 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 56.470 6.490 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 47.800 6.490 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 52.495 6.545 52.815 ;
      LAYER met4 ;
        RECT 6.225 52.495 6.545 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 52.075 6.545 52.395 ;
      LAYER met4 ;
        RECT 6.225 52.075 6.545 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 51.655 6.545 51.975 ;
      LAYER met4 ;
        RECT 6.225 51.655 6.545 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 39.900 6.120 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 39.460 6.120 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 39.020 6.120 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 38.580 6.120 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 38.140 6.120 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 37.700 6.120 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 37.260 6.120 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.920 36.820 6.120 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 56.470 6.085 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 47.800 6.085 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 52.495 6.140 52.815 ;
      LAYER met4 ;
        RECT 5.820 52.495 6.140 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 52.075 6.140 52.395 ;
      LAYER met4 ;
        RECT 5.820 52.075 6.140 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 51.655 6.140 51.975 ;
      LAYER met4 ;
        RECT 5.820 51.655 6.140 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 39.900 5.715 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 39.460 5.715 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 39.020 5.715 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 38.580 5.715 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 38.140 5.715 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 37.700 5.715 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 37.260 5.715 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.515 36.820 5.715 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 56.470 5.680 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 47.800 5.680 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 52.495 5.735 52.815 ;
      LAYER met4 ;
        RECT 5.415 52.495 5.735 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 52.075 5.735 52.395 ;
      LAYER met4 ;
        RECT 5.415 52.075 5.735 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 51.655 5.735 51.975 ;
      LAYER met4 ;
        RECT 5.415 51.655 5.735 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 39.900 5.310 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 39.460 5.310 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 39.020 5.310 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 38.580 5.310 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 38.140 5.310 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 37.700 5.310 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 37.260 5.310 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.110 36.820 5.310 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 56.470 5.275 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 47.800 5.275 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 52.495 5.330 52.815 ;
      LAYER met4 ;
        RECT 5.010 52.495 5.330 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 52.075 5.330 52.395 ;
      LAYER met4 ;
        RECT 5.010 52.075 5.330 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 51.655 5.330 51.975 ;
      LAYER met4 ;
        RECT 5.010 51.655 5.330 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 39.900 4.905 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 39.460 4.905 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 39.020 4.905 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 38.580 4.905 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 38.140 4.905 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 37.700 4.905 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 37.260 4.905 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.705 36.820 4.905 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 56.470 4.870 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 47.800 4.870 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 52.495 4.925 52.815 ;
      LAYER met4 ;
        RECT 4.605 52.495 4.925 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 52.075 4.925 52.395 ;
      LAYER met4 ;
        RECT 4.605 52.075 4.925 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 51.655 4.925 51.975 ;
      LAYER met4 ;
        RECT 4.605 51.655 4.925 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 39.900 4.500 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 39.460 4.500 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 39.020 4.500 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 38.580 4.500 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 38.140 4.500 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 37.700 4.500 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 37.260 4.500 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.300 36.820 4.500 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 56.470 4.465 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 47.800 4.465 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 52.495 4.520 52.815 ;
      LAYER met4 ;
        RECT 4.200 52.495 4.520 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 52.075 4.520 52.395 ;
      LAYER met4 ;
        RECT 4.200 52.075 4.520 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 51.655 4.520 51.975 ;
      LAYER met4 ;
        RECT 4.200 51.655 4.520 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 39.900 4.095 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 39.460 4.095 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 39.020 4.095 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 38.580 4.095 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 38.140 4.095 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 37.700 4.095 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 37.260 4.095 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.895 36.820 4.095 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 56.470 4.060 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 47.800 4.060 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 52.495 4.115 52.815 ;
      LAYER met4 ;
        RECT 3.795 52.495 4.115 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 52.075 4.115 52.395 ;
      LAYER met4 ;
        RECT 3.795 52.075 4.115 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 51.655 4.115 51.975 ;
      LAYER met4 ;
        RECT 3.795 51.655 4.115 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 39.900 3.690 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 39.460 3.690 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 39.020 3.690 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 38.580 3.690 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 38.140 3.690 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 37.700 3.690 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 37.260 3.690 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.490 36.820 3.690 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 56.470 3.655 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 47.800 3.655 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 52.495 3.710 52.815 ;
      LAYER met4 ;
        RECT 3.390 52.495 3.710 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 52.075 3.710 52.395 ;
      LAYER met4 ;
        RECT 3.390 52.075 3.710 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 51.655 3.710 51.975 ;
      LAYER met4 ;
        RECT 3.390 51.655 3.710 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 39.900 3.285 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 39.460 3.285 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 39.020 3.285 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 38.580 3.285 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 38.140 3.285 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 37.700 3.285 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 37.260 3.285 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.085 36.820 3.285 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 56.470 3.250 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 47.800 3.250 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 52.495 3.305 52.815 ;
      LAYER met4 ;
        RECT 2.985 52.495 3.305 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 52.075 3.305 52.395 ;
      LAYER met4 ;
        RECT 2.985 52.075 3.305 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 51.655 3.305 51.975 ;
      LAYER met4 ;
        RECT 2.985 51.655 3.305 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 39.900 2.880 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 39.460 2.880 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 39.020 2.880 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 38.580 2.880 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 38.140 2.880 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 37.700 2.880 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 37.260 2.880 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.680 36.820 2.880 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.645 56.470 2.845 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.645 47.800 2.845 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 52.495 2.895 52.815 ;
      LAYER met4 ;
        RECT 2.575 52.495 2.895 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 52.075 2.895 52.395 ;
      LAYER met4 ;
        RECT 2.575 52.075 2.895 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 51.655 2.895 51.975 ;
      LAYER met4 ;
        RECT 2.575 51.655 2.895 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 39.900 2.475 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 39.460 2.475 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 39.020 2.475 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 38.580 2.475 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 38.140 2.475 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 37.700 2.475 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 37.260 2.475 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.275 36.820 2.475 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.240 56.470 2.440 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.240 47.800 2.440 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 52.495 2.485 52.815 ;
      LAYER met4 ;
        RECT 2.165 52.495 2.485 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 52.075 2.485 52.395 ;
      LAYER met4 ;
        RECT 2.165 52.075 2.485 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 51.655 2.485 51.975 ;
      LAYER met4 ;
        RECT 2.165 51.655 2.485 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 39.900 2.070 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 39.460 2.070 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 39.020 2.070 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 38.580 2.070 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 38.140 2.070 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 37.700 2.070 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 37.260 2.070 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.870 36.820 2.070 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.835 56.470 2.035 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.835 47.800 2.035 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 52.495 2.075 52.815 ;
      LAYER met4 ;
        RECT 1.755 52.495 2.075 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 52.075 2.075 52.395 ;
      LAYER met4 ;
        RECT 1.755 52.075 2.075 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 51.655 2.075 51.975 ;
      LAYER met4 ;
        RECT 1.755 51.655 2.075 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 39.900 1.665 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 39.460 1.665 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 39.020 1.665 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 38.580 1.665 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 38.140 1.665 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 37.700 1.665 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 37.260 1.665 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.465 36.820 1.665 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.430 56.470 1.630 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.430 47.800 1.630 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 52.495 1.665 52.815 ;
      LAYER met4 ;
        RECT 1.345 52.495 1.665 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 52.075 1.665 52.395 ;
      LAYER met4 ;
        RECT 1.345 52.075 1.665 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 51.655 1.665 51.975 ;
      LAYER met4 ;
        RECT 1.345 51.655 1.665 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 39.900 1.260 40.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 39.460 1.260 39.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 39.020 1.260 39.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 38.580 1.260 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 38.140 1.260 38.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 37.700 1.260 37.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 37.260 1.260 37.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.060 36.820 1.260 37.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 56.470 1.225 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 47.800 1.225 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 52.495 1.255 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 52.075 1.255 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 51.655 1.255 51.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.620 56.470 0.820 56.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.620 47.800 0.820 48.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 52.495 0.845 52.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 52.075 0.845 52.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 51.655 0.845 51.975 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
  END VSSD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  OBS
      LAYER met3 ;
        RECT 0.495 51.650 24.395 52.820 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 56.505 73.330 57.135 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 1.670 47.335 73.330 47.965 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 96.585 75.000 174.185 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__overlay_vssa_hvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vssa_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vssa_lvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
  END VDDIO_Q
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
  END VCCD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 49.650 24.400 50.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 34.740 74.655 38.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 49.650 74.655 50.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 50.555 74.565 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 50.135 74.565 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 49.715 74.565 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 37.900 74.565 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 37.460 74.565 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 37.020 74.565 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 36.580 74.565 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 36.140 74.565 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 35.700 74.565 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 35.260 74.565 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.365 34.820 74.565 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 50.555 74.160 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 50.135 74.160 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 49.715 74.160 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 37.900 74.160 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 37.460 74.160 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 37.020 74.160 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 36.580 74.160 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 36.140 74.160 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 35.700 74.160 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 35.260 74.160 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.960 34.820 74.160 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 50.555 73.755 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 50.135 73.755 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 49.715 73.755 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 37.900 73.755 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 37.460 73.755 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 37.020 73.755 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 36.580 73.755 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 36.140 73.755 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 35.700 73.755 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 35.260 73.755 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.555 34.820 73.755 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 50.555 73.350 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 50.135 73.350 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 49.715 73.350 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 37.900 73.350 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 37.460 73.350 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 37.020 73.350 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 36.580 73.350 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 36.140 73.350 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 35.700 73.350 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 35.260 73.350 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.150 34.820 73.350 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 50.555 72.945 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 50.135 72.945 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 49.715 72.945 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 37.900 72.945 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 37.460 72.945 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 37.020 72.945 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 36.580 72.945 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 36.140 72.945 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 35.700 72.945 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 35.260 72.945 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.745 34.820 72.945 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 50.555 72.540 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 50.135 72.540 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 49.715 72.540 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 37.900 72.540 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 37.460 72.540 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 37.020 72.540 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 36.580 72.540 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 36.140 72.540 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 35.700 72.540 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 35.260 72.540 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.340 34.820 72.540 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 50.555 72.135 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 50.135 72.135 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 49.715 72.135 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 37.900 72.135 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 37.460 72.135 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 37.020 72.135 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 36.580 72.135 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 36.140 72.135 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 35.700 72.135 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 35.260 72.135 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.935 34.820 72.135 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 50.555 71.730 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 50.135 71.730 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 49.715 71.730 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 37.900 71.730 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 37.460 71.730 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 37.020 71.730 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 36.580 71.730 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 36.140 71.730 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 35.700 71.730 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 35.260 71.730 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 34.820 71.730 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 50.555 71.325 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 50.135 71.325 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 49.715 71.325 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 37.900 71.325 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 37.460 71.325 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 37.020 71.325 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 36.580 71.325 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 36.140 71.325 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 35.700 71.325 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 35.260 71.325 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.125 34.820 71.325 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 50.555 70.920 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 50.135 70.920 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 49.715 70.920 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 37.900 70.920 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 37.460 70.920 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 37.020 70.920 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 36.580 70.920 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 36.140 70.920 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 35.700 70.920 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 35.260 70.920 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.720 34.820 70.920 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 50.555 70.515 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 50.135 70.515 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 49.715 70.515 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 37.900 70.515 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 37.460 70.515 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 37.020 70.515 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 36.580 70.515 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 36.140 70.515 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 35.700 70.515 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 35.260 70.515 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.315 34.820 70.515 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 50.555 70.110 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 50.135 70.110 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 49.715 70.110 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 37.900 70.110 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 37.460 70.110 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 37.020 70.110 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 36.580 70.110 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 36.140 70.110 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 35.700 70.110 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 35.260 70.110 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.910 34.820 70.110 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 50.555 69.705 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 50.135 69.705 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 49.715 69.705 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 37.900 69.705 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 37.460 69.705 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 37.020 69.705 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 36.580 69.705 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 36.140 69.705 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 35.700 69.705 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 35.260 69.705 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.505 34.820 69.705 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 50.555 69.300 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 50.135 69.300 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 49.715 69.300 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 37.900 69.300 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 37.460 69.300 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 37.020 69.300 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 36.580 69.300 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 36.140 69.300 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 35.700 69.300 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 35.260 69.300 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.100 34.820 69.300 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 50.555 68.895 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 50.135 68.895 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 49.715 68.895 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 37.900 68.895 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 37.460 68.895 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 37.020 68.895 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 36.580 68.895 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 36.140 68.895 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 35.700 68.895 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 35.260 68.895 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.695 34.820 68.895 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 50.555 68.490 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 50.135 68.490 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 49.715 68.490 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 37.900 68.490 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 37.460 68.490 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 37.020 68.490 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 36.580 68.490 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 36.140 68.490 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 35.700 68.490 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 35.260 68.490 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 34.820 68.490 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 50.555 68.085 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 50.135 68.085 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 49.715 68.085 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 37.900 68.085 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 37.460 68.085 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 37.020 68.085 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 36.580 68.085 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 36.140 68.085 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 35.700 68.085 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 35.260 68.085 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.885 34.820 68.085 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 50.555 67.680 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 50.135 67.680 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 49.715 67.680 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 37.900 67.680 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 37.460 67.680 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 37.020 67.680 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 36.580 67.680 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 36.140 67.680 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 35.700 67.680 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 35.260 67.680 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.480 34.820 67.680 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 50.555 67.275 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 50.135 67.275 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 49.715 67.275 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 37.900 67.275 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 37.460 67.275 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 37.020 67.275 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 36.580 67.275 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 36.140 67.275 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 35.700 67.275 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 35.260 67.275 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.075 34.820 67.275 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 50.555 66.870 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 50.135 66.870 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 49.715 66.870 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 37.900 66.870 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 37.460 66.870 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 37.020 66.870 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 36.580 66.870 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 36.140 66.870 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 35.700 66.870 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 35.260 66.870 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.670 34.820 66.870 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 50.555 66.465 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 50.135 66.465 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 49.715 66.465 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 37.900 66.465 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 37.460 66.465 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 37.020 66.465 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 36.580 66.465 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 36.140 66.465 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 35.700 66.465 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 35.260 66.465 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.265 34.820 66.465 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 50.555 66.060 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 50.135 66.060 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 49.715 66.060 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 37.900 66.060 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 37.460 66.060 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 37.020 66.060 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 36.580 66.060 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 36.140 66.060 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 35.700 66.060 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 35.260 66.060 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.860 34.820 66.060 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 50.555 65.655 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 50.135 65.655 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 49.715 65.655 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 37.900 65.655 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 37.460 65.655 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 37.020 65.655 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 36.580 65.655 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 36.140 65.655 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 35.700 65.655 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 35.260 65.655 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.455 34.820 65.655 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 50.555 65.250 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 50.135 65.250 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 49.715 65.250 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 37.900 65.250 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 37.460 65.250 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 37.020 65.250 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 36.580 65.250 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 36.140 65.250 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 35.700 65.250 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 35.260 65.250 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.050 34.820 65.250 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 50.555 64.845 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 50.135 64.845 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 49.715 64.845 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 37.900 64.845 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 37.460 64.845 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 37.020 64.845 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 36.580 64.845 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 36.140 64.845 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 35.700 64.845 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 35.260 64.845 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.645 34.820 64.845 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 50.555 64.440 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 50.135 64.440 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 49.715 64.440 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 37.900 64.440 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 37.460 64.440 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 37.020 64.440 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 36.580 64.440 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 36.140 64.440 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 35.700 64.440 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 35.260 64.440 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.240 34.820 64.440 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 50.555 64.035 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 50.135 64.035 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 49.715 64.035 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 37.900 64.035 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 37.460 64.035 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 37.020 64.035 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 36.580 64.035 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 36.140 64.035 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 35.700 64.035 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 35.260 64.035 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.835 34.820 64.035 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 50.555 63.630 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 50.135 63.630 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 49.715 63.630 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 37.900 63.630 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 37.460 63.630 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 37.020 63.630 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 36.580 63.630 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 36.140 63.630 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 35.700 63.630 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 35.260 63.630 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.430 34.820 63.630 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 50.555 63.225 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 50.135 63.225 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 49.715 63.225 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 37.900 63.225 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 37.460 63.225 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 37.020 63.225 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 36.580 63.225 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 36.140 63.225 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 35.700 63.225 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 35.260 63.225 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.025 34.820 63.225 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 50.555 62.820 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 50.135 62.820 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 49.715 62.820 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 37.900 62.820 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 37.460 62.820 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 37.020 62.820 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 36.580 62.820 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 36.140 62.820 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 35.700 62.820 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 35.260 62.820 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.620 34.820 62.820 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 50.555 62.415 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 50.135 62.415 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 49.715 62.415 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 37.900 62.415 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 37.460 62.415 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 37.020 62.415 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 36.580 62.415 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 36.140 62.415 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 35.700 62.415 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 35.260 62.415 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.215 34.820 62.415 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 50.555 62.010 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 50.135 62.010 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 49.715 62.010 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 37.900 62.010 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 37.460 62.010 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 37.020 62.010 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 36.580 62.010 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 36.140 62.010 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 35.700 62.010 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 35.260 62.010 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.810 34.820 62.010 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 50.555 61.605 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 50.135 61.605 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 49.715 61.605 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 37.900 61.605 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 37.460 61.605 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 37.020 61.605 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 36.580 61.605 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 36.140 61.605 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 35.700 61.605 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 35.260 61.605 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.405 34.820 61.605 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 50.555 61.200 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 50.135 61.200 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 49.715 61.200 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 37.900 61.200 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 37.460 61.200 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 37.020 61.200 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 36.580 61.200 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 36.140 61.200 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 35.700 61.200 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 35.260 61.200 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.000 34.820 61.200 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 50.555 60.795 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 50.135 60.795 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 49.715 60.795 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 37.900 60.795 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 37.460 60.795 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 37.020 60.795 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 36.580 60.795 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 36.140 60.795 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 35.700 60.795 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 35.260 60.795 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.595 34.820 60.795 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 50.555 60.390 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 50.135 60.390 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 49.715 60.390 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 37.900 60.390 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 37.460 60.390 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 37.020 60.390 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 36.580 60.390 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 36.140 60.390 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 35.700 60.390 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 35.260 60.390 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.190 34.820 60.390 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 50.555 59.985 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 50.135 59.985 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 49.715 59.985 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 37.900 59.985 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 37.460 59.985 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 37.020 59.985 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 36.580 59.985 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 36.140 59.985 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 35.700 59.985 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 35.260 59.985 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.785 34.820 59.985 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 50.555 59.580 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 50.135 59.580 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 49.715 59.580 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 37.900 59.580 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 37.460 59.580 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 37.020 59.580 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 36.580 59.580 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 36.140 59.580 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 35.700 59.580 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 35.260 59.580 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.380 34.820 59.580 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 50.555 59.175 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 50.135 59.175 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 49.715 59.175 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 37.900 59.175 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 37.460 59.175 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 37.020 59.175 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 36.580 59.175 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 36.140 59.175 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 35.700 59.175 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 35.260 59.175 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.975 34.820 59.175 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 50.555 58.770 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 50.135 58.770 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 49.715 58.770 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 37.900 58.770 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 37.460 58.770 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 37.020 58.770 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 36.580 58.770 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 36.140 58.770 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 35.700 58.770 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 35.260 58.770 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.570 34.820 58.770 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 50.555 58.365 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 50.135 58.365 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 49.715 58.365 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 37.900 58.365 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 37.460 58.365 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 37.020 58.365 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 36.580 58.365 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 36.140 58.365 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 35.700 58.365 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 35.260 58.365 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.165 34.820 58.365 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 50.555 57.960 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 50.135 57.960 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 49.715 57.960 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 37.900 57.960 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 37.460 57.960 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 37.020 57.960 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 36.580 57.960 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 36.140 57.960 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 35.700 57.960 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 35.260 57.960 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.760 34.820 57.960 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 50.555 57.555 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 50.135 57.555 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 49.715 57.555 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 37.900 57.555 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 37.460 57.555 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 37.020 57.555 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 36.580 57.555 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 36.140 57.555 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 35.700 57.555 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 35.260 57.555 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.355 34.820 57.555 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 50.555 57.150 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 50.135 57.150 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 49.715 57.150 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 37.900 57.150 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 37.460 57.150 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 37.020 57.150 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 36.580 57.150 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 36.140 57.150 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 35.700 57.150 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 35.260 57.150 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.950 34.820 57.150 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 50.555 56.745 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 50.135 56.745 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 49.715 56.745 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 37.900 56.745 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 37.460 56.745 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 37.020 56.745 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 36.580 56.745 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 36.140 56.745 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 35.700 56.745 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 35.260 56.745 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.545 34.820 56.745 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 50.555 56.340 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 50.135 56.340 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 49.715 56.340 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 37.900 56.340 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 37.460 56.340 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 37.020 56.340 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 36.580 56.340 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 36.140 56.340 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 35.700 56.340 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 35.260 56.340 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.140 34.820 56.340 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 50.555 55.935 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 50.135 55.935 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 49.715 55.935 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 37.900 55.935 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 37.460 55.935 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 37.020 55.935 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 36.580 55.935 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 36.140 55.935 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 35.700 55.935 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 35.260 55.935 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.735 34.820 55.935 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 50.555 55.530 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 50.135 55.530 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 49.715 55.530 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 37.900 55.530 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 37.460 55.530 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 37.020 55.530 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 36.580 55.530 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 36.140 55.530 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 35.700 55.530 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 35.260 55.530 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.330 34.820 55.530 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 50.555 55.125 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 50.135 55.125 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 49.715 55.125 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 37.900 55.125 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 37.460 55.125 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 37.020 55.125 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 36.580 55.125 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 36.140 55.125 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 35.700 55.125 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 35.260 55.125 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.925 34.820 55.125 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 50.555 54.720 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 50.135 54.720 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 49.715 54.720 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 37.900 54.720 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 37.460 54.720 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 37.020 54.720 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 36.580 54.720 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 36.140 54.720 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 35.700 54.720 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 35.260 54.720 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.520 34.820 54.720 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 50.555 54.315 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 50.135 54.315 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 49.715 54.315 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 37.900 54.315 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 37.460 54.315 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 37.020 54.315 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 36.580 54.315 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 36.140 54.315 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 35.700 54.315 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 35.260 54.315 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.115 34.820 54.315 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 50.555 53.910 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 50.135 53.910 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 49.715 53.910 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 37.900 53.910 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 37.460 53.910 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 37.020 53.910 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 36.580 53.910 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 36.140 53.910 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 35.700 53.910 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 35.260 53.910 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.710 34.820 53.910 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 50.555 53.505 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 50.135 53.505 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 49.715 53.505 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 37.900 53.505 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 37.460 53.505 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 37.020 53.505 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 36.580 53.505 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 36.140 53.505 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 35.700 53.505 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 35.260 53.505 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 34.820 53.505 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 50.555 53.095 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 50.135 53.095 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 49.715 53.095 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 37.900 53.095 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 37.460 53.095 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 37.020 53.095 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 36.580 53.095 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 36.140 53.095 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 35.700 53.095 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 35.260 53.095 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 34.820 53.095 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 50.555 52.685 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 50.135 52.685 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 49.715 52.685 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 37.900 52.685 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 37.460 52.685 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 37.020 52.685 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 36.580 52.685 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 36.140 52.685 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 35.700 52.685 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 35.260 52.685 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 34.820 52.685 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 50.555 52.275 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 50.135 52.275 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 49.715 52.275 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 37.900 52.275 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 37.460 52.275 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 37.020 52.275 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 36.580 52.275 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 36.140 52.275 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 35.700 52.275 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 35.260 52.275 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 34.820 52.275 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 50.555 51.865 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 50.135 51.865 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 49.715 51.865 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 37.900 51.865 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 37.460 51.865 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 37.020 51.865 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 36.580 51.865 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 36.140 51.865 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 35.700 51.865 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 35.260 51.865 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 34.820 51.865 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 50.555 51.455 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 50.135 51.455 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 49.715 51.455 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 37.900 51.455 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 37.460 51.455 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 37.020 51.455 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 36.580 51.455 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 36.140 51.455 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 35.700 51.455 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 35.260 51.455 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 34.820 51.455 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 50.555 51.045 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 50.135 51.045 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 49.715 51.045 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 37.900 51.045 38.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 37.460 51.045 37.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 37.020 51.045 37.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 36.580 51.045 36.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 36.140 51.045 36.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 35.700 51.045 35.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 35.260 51.045 35.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 34.820 51.045 35.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 50.555 24.310 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 50.135 24.310 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 49.715 24.310 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 37.840 24.370 38.160 ;
      LAYER met4 ;
        RECT 24.050 37.840 24.370 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 37.400 24.370 37.720 ;
      LAYER met4 ;
        RECT 24.050 37.400 24.370 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 36.960 24.370 37.280 ;
      LAYER met4 ;
        RECT 24.050 36.960 24.370 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 36.520 24.370 36.840 ;
      LAYER met4 ;
        RECT 24.050 36.520 24.370 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 36.080 24.370 36.400 ;
      LAYER met4 ;
        RECT 24.050 36.080 24.370 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 35.640 24.370 35.960 ;
      LAYER met4 ;
        RECT 24.050 35.640 24.370 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 35.200 24.370 35.520 ;
      LAYER met4 ;
        RECT 24.050 35.200 24.370 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 34.760 24.370 35.080 ;
      LAYER met4 ;
        RECT 24.050 34.760 24.370 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 50.555 23.905 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 50.135 23.905 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 49.715 23.905 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 37.840 23.965 38.160 ;
      LAYER met4 ;
        RECT 23.645 37.840 23.965 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 37.400 23.965 37.720 ;
      LAYER met4 ;
        RECT 23.645 37.400 23.965 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 36.960 23.965 37.280 ;
      LAYER met4 ;
        RECT 23.645 36.960 23.965 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 36.520 23.965 36.840 ;
      LAYER met4 ;
        RECT 23.645 36.520 23.965 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 36.080 23.965 36.400 ;
      LAYER met4 ;
        RECT 23.645 36.080 23.965 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 35.640 23.965 35.960 ;
      LAYER met4 ;
        RECT 23.645 35.640 23.965 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 35.200 23.965 35.520 ;
      LAYER met4 ;
        RECT 23.645 35.200 23.965 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 34.760 23.965 35.080 ;
      LAYER met4 ;
        RECT 23.645 34.760 23.965 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 50.555 23.500 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 50.135 23.500 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 49.715 23.500 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 37.840 23.560 38.160 ;
      LAYER met4 ;
        RECT 23.240 37.840 23.560 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 37.400 23.560 37.720 ;
      LAYER met4 ;
        RECT 23.240 37.400 23.560 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 36.960 23.560 37.280 ;
      LAYER met4 ;
        RECT 23.240 36.960 23.560 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 36.520 23.560 36.840 ;
      LAYER met4 ;
        RECT 23.240 36.520 23.560 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 36.080 23.560 36.400 ;
      LAYER met4 ;
        RECT 23.240 36.080 23.560 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 35.640 23.560 35.960 ;
      LAYER met4 ;
        RECT 23.240 35.640 23.560 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 35.200 23.560 35.520 ;
      LAYER met4 ;
        RECT 23.240 35.200 23.560 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 34.760 23.560 35.080 ;
      LAYER met4 ;
        RECT 23.240 34.760 23.560 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 50.555 23.095 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 50.135 23.095 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 49.715 23.095 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 37.840 23.155 38.160 ;
      LAYER met4 ;
        RECT 22.835 37.840 23.155 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 37.400 23.155 37.720 ;
      LAYER met4 ;
        RECT 22.835 37.400 23.155 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 36.960 23.155 37.280 ;
      LAYER met4 ;
        RECT 22.835 36.960 23.155 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 36.520 23.155 36.840 ;
      LAYER met4 ;
        RECT 22.835 36.520 23.155 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 36.080 23.155 36.400 ;
      LAYER met4 ;
        RECT 22.835 36.080 23.155 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 35.640 23.155 35.960 ;
      LAYER met4 ;
        RECT 22.835 35.640 23.155 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 35.200 23.155 35.520 ;
      LAYER met4 ;
        RECT 22.835 35.200 23.155 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 34.760 23.155 35.080 ;
      LAYER met4 ;
        RECT 22.835 34.760 23.155 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 50.555 22.690 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 50.135 22.690 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 49.715 22.690 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 37.840 22.750 38.160 ;
      LAYER met4 ;
        RECT 22.430 37.840 22.750 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 37.400 22.750 37.720 ;
      LAYER met4 ;
        RECT 22.430 37.400 22.750 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 36.960 22.750 37.280 ;
      LAYER met4 ;
        RECT 22.430 36.960 22.750 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 36.520 22.750 36.840 ;
      LAYER met4 ;
        RECT 22.430 36.520 22.750 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 36.080 22.750 36.400 ;
      LAYER met4 ;
        RECT 22.430 36.080 22.750 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 35.640 22.750 35.960 ;
      LAYER met4 ;
        RECT 22.430 35.640 22.750 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 35.200 22.750 35.520 ;
      LAYER met4 ;
        RECT 22.430 35.200 22.750 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 34.760 22.750 35.080 ;
      LAYER met4 ;
        RECT 22.430 34.760 22.750 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 50.555 22.285 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 50.135 22.285 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 49.715 22.285 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 37.840 22.345 38.160 ;
      LAYER met4 ;
        RECT 22.025 37.840 22.345 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 37.400 22.345 37.720 ;
      LAYER met4 ;
        RECT 22.025 37.400 22.345 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 36.960 22.345 37.280 ;
      LAYER met4 ;
        RECT 22.025 36.960 22.345 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 36.520 22.345 36.840 ;
      LAYER met4 ;
        RECT 22.025 36.520 22.345 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 36.080 22.345 36.400 ;
      LAYER met4 ;
        RECT 22.025 36.080 22.345 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 35.640 22.345 35.960 ;
      LAYER met4 ;
        RECT 22.025 35.640 22.345 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 35.200 22.345 35.520 ;
      LAYER met4 ;
        RECT 22.025 35.200 22.345 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 34.760 22.345 35.080 ;
      LAYER met4 ;
        RECT 22.025 34.760 22.345 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 50.555 21.880 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 50.135 21.880 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 49.715 21.880 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 37.840 21.940 38.160 ;
      LAYER met4 ;
        RECT 21.620 37.840 21.940 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 37.400 21.940 37.720 ;
      LAYER met4 ;
        RECT 21.620 37.400 21.940 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 36.960 21.940 37.280 ;
      LAYER met4 ;
        RECT 21.620 36.960 21.940 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 36.520 21.940 36.840 ;
      LAYER met4 ;
        RECT 21.620 36.520 21.940 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 36.080 21.940 36.400 ;
      LAYER met4 ;
        RECT 21.620 36.080 21.940 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 35.640 21.940 35.960 ;
      LAYER met4 ;
        RECT 21.620 35.640 21.940 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 35.200 21.940 35.520 ;
      LAYER met4 ;
        RECT 21.620 35.200 21.940 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 34.760 21.940 35.080 ;
      LAYER met4 ;
        RECT 21.620 34.760 21.940 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 50.555 21.475 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 50.135 21.475 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 49.715 21.475 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 37.840 21.535 38.160 ;
      LAYER met4 ;
        RECT 21.215 37.840 21.535 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 37.400 21.535 37.720 ;
      LAYER met4 ;
        RECT 21.215 37.400 21.535 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 36.960 21.535 37.280 ;
      LAYER met4 ;
        RECT 21.215 36.960 21.535 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 36.520 21.535 36.840 ;
      LAYER met4 ;
        RECT 21.215 36.520 21.535 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 36.080 21.535 36.400 ;
      LAYER met4 ;
        RECT 21.215 36.080 21.535 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 35.640 21.535 35.960 ;
      LAYER met4 ;
        RECT 21.215 35.640 21.535 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 35.200 21.535 35.520 ;
      LAYER met4 ;
        RECT 21.215 35.200 21.535 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 34.760 21.535 35.080 ;
      LAYER met4 ;
        RECT 21.215 34.760 21.535 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 50.555 21.070 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 50.135 21.070 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 49.715 21.070 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 37.840 21.130 38.160 ;
      LAYER met4 ;
        RECT 20.810 37.840 21.130 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 37.400 21.130 37.720 ;
      LAYER met4 ;
        RECT 20.810 37.400 21.130 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 36.960 21.130 37.280 ;
      LAYER met4 ;
        RECT 20.810 36.960 21.130 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 36.520 21.130 36.840 ;
      LAYER met4 ;
        RECT 20.810 36.520 21.130 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 36.080 21.130 36.400 ;
      LAYER met4 ;
        RECT 20.810 36.080 21.130 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 35.640 21.130 35.960 ;
      LAYER met4 ;
        RECT 20.810 35.640 21.130 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 35.200 21.130 35.520 ;
      LAYER met4 ;
        RECT 20.810 35.200 21.130 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 34.760 21.130 35.080 ;
      LAYER met4 ;
        RECT 20.810 34.760 21.130 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 50.555 20.665 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 50.135 20.665 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 49.715 20.665 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 37.840 20.725 38.160 ;
      LAYER met4 ;
        RECT 20.405 37.840 20.725 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 37.400 20.725 37.720 ;
      LAYER met4 ;
        RECT 20.405 37.400 20.725 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 36.960 20.725 37.280 ;
      LAYER met4 ;
        RECT 20.405 36.960 20.725 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 36.520 20.725 36.840 ;
      LAYER met4 ;
        RECT 20.405 36.520 20.725 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 36.080 20.725 36.400 ;
      LAYER met4 ;
        RECT 20.405 36.080 20.725 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 35.640 20.725 35.960 ;
      LAYER met4 ;
        RECT 20.405 35.640 20.725 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 35.200 20.725 35.520 ;
      LAYER met4 ;
        RECT 20.405 35.200 20.725 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 34.760 20.725 35.080 ;
      LAYER met4 ;
        RECT 20.405 34.760 20.725 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 50.555 20.260 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 50.135 20.260 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 49.715 20.260 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 37.840 20.320 38.160 ;
      LAYER met4 ;
        RECT 20.000 37.840 20.320 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 37.400 20.320 37.720 ;
      LAYER met4 ;
        RECT 20.000 37.400 20.320 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 36.960 20.320 37.280 ;
      LAYER met4 ;
        RECT 20.000 36.960 20.320 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 36.520 20.320 36.840 ;
      LAYER met4 ;
        RECT 20.000 36.520 20.320 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 36.080 20.320 36.400 ;
      LAYER met4 ;
        RECT 20.000 36.080 20.320 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 35.640 20.320 35.960 ;
      LAYER met4 ;
        RECT 20.000 35.640 20.320 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 35.200 20.320 35.520 ;
      LAYER met4 ;
        RECT 20.000 35.200 20.320 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 34.760 20.320 35.080 ;
      LAYER met4 ;
        RECT 20.000 34.760 20.320 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 50.555 19.855 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 50.135 19.855 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 49.715 19.855 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 37.840 19.915 38.160 ;
      LAYER met4 ;
        RECT 19.595 37.840 19.915 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 37.400 19.915 37.720 ;
      LAYER met4 ;
        RECT 19.595 37.400 19.915 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 36.960 19.915 37.280 ;
      LAYER met4 ;
        RECT 19.595 36.960 19.915 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 36.520 19.915 36.840 ;
      LAYER met4 ;
        RECT 19.595 36.520 19.915 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 36.080 19.915 36.400 ;
      LAYER met4 ;
        RECT 19.595 36.080 19.915 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 35.640 19.915 35.960 ;
      LAYER met4 ;
        RECT 19.595 35.640 19.915 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 35.200 19.915 35.520 ;
      LAYER met4 ;
        RECT 19.595 35.200 19.915 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 34.760 19.915 35.080 ;
      LAYER met4 ;
        RECT 19.595 34.760 19.915 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 50.555 19.450 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 50.135 19.450 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 49.715 19.450 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 37.840 19.510 38.160 ;
      LAYER met4 ;
        RECT 19.190 37.840 19.510 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 37.400 19.510 37.720 ;
      LAYER met4 ;
        RECT 19.190 37.400 19.510 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 36.960 19.510 37.280 ;
      LAYER met4 ;
        RECT 19.190 36.960 19.510 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 36.520 19.510 36.840 ;
      LAYER met4 ;
        RECT 19.190 36.520 19.510 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 36.080 19.510 36.400 ;
      LAYER met4 ;
        RECT 19.190 36.080 19.510 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 35.640 19.510 35.960 ;
      LAYER met4 ;
        RECT 19.190 35.640 19.510 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 35.200 19.510 35.520 ;
      LAYER met4 ;
        RECT 19.190 35.200 19.510 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 34.760 19.510 35.080 ;
      LAYER met4 ;
        RECT 19.190 34.760 19.510 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 50.555 19.045 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 50.135 19.045 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 49.715 19.045 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 37.840 19.105 38.160 ;
      LAYER met4 ;
        RECT 18.785 37.840 19.105 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 37.400 19.105 37.720 ;
      LAYER met4 ;
        RECT 18.785 37.400 19.105 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 36.960 19.105 37.280 ;
      LAYER met4 ;
        RECT 18.785 36.960 19.105 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 36.520 19.105 36.840 ;
      LAYER met4 ;
        RECT 18.785 36.520 19.105 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 36.080 19.105 36.400 ;
      LAYER met4 ;
        RECT 18.785 36.080 19.105 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 35.640 19.105 35.960 ;
      LAYER met4 ;
        RECT 18.785 35.640 19.105 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 35.200 19.105 35.520 ;
      LAYER met4 ;
        RECT 18.785 35.200 19.105 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 34.760 19.105 35.080 ;
      LAYER met4 ;
        RECT 18.785 34.760 19.105 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 50.555 18.640 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 50.135 18.640 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 49.715 18.640 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 37.840 18.700 38.160 ;
      LAYER met4 ;
        RECT 18.380 37.840 18.700 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 37.400 18.700 37.720 ;
      LAYER met4 ;
        RECT 18.380 37.400 18.700 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 36.960 18.700 37.280 ;
      LAYER met4 ;
        RECT 18.380 36.960 18.700 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 36.520 18.700 36.840 ;
      LAYER met4 ;
        RECT 18.380 36.520 18.700 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 36.080 18.700 36.400 ;
      LAYER met4 ;
        RECT 18.380 36.080 18.700 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 35.640 18.700 35.960 ;
      LAYER met4 ;
        RECT 18.380 35.640 18.700 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 35.200 18.700 35.520 ;
      LAYER met4 ;
        RECT 18.380 35.200 18.700 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 34.760 18.700 35.080 ;
      LAYER met4 ;
        RECT 18.380 34.760 18.700 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 50.555 18.235 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 50.135 18.235 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 49.715 18.235 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 37.840 18.295 38.160 ;
      LAYER met4 ;
        RECT 17.975 37.840 18.295 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 37.400 18.295 37.720 ;
      LAYER met4 ;
        RECT 17.975 37.400 18.295 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 36.960 18.295 37.280 ;
      LAYER met4 ;
        RECT 17.975 36.960 18.295 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 36.520 18.295 36.840 ;
      LAYER met4 ;
        RECT 17.975 36.520 18.295 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 36.080 18.295 36.400 ;
      LAYER met4 ;
        RECT 17.975 36.080 18.295 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 35.640 18.295 35.960 ;
      LAYER met4 ;
        RECT 17.975 35.640 18.295 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 35.200 18.295 35.520 ;
      LAYER met4 ;
        RECT 17.975 35.200 18.295 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 34.760 18.295 35.080 ;
      LAYER met4 ;
        RECT 17.975 34.760 18.295 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 50.555 17.830 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 50.135 17.830 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 49.715 17.830 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 37.840 17.890 38.160 ;
      LAYER met4 ;
        RECT 17.570 37.840 17.890 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 37.400 17.890 37.720 ;
      LAYER met4 ;
        RECT 17.570 37.400 17.890 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 36.960 17.890 37.280 ;
      LAYER met4 ;
        RECT 17.570 36.960 17.890 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 36.520 17.890 36.840 ;
      LAYER met4 ;
        RECT 17.570 36.520 17.890 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 36.080 17.890 36.400 ;
      LAYER met4 ;
        RECT 17.570 36.080 17.890 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 35.640 17.890 35.960 ;
      LAYER met4 ;
        RECT 17.570 35.640 17.890 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 35.200 17.890 35.520 ;
      LAYER met4 ;
        RECT 17.570 35.200 17.890 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 34.760 17.890 35.080 ;
      LAYER met4 ;
        RECT 17.570 34.760 17.890 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 50.555 17.425 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 50.135 17.425 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 49.715 17.425 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 37.840 17.485 38.160 ;
      LAYER met4 ;
        RECT 17.165 37.840 17.485 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 37.400 17.485 37.720 ;
      LAYER met4 ;
        RECT 17.165 37.400 17.485 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 36.960 17.485 37.280 ;
      LAYER met4 ;
        RECT 17.165 36.960 17.485 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 36.520 17.485 36.840 ;
      LAYER met4 ;
        RECT 17.165 36.520 17.485 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 36.080 17.485 36.400 ;
      LAYER met4 ;
        RECT 17.165 36.080 17.485 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 35.640 17.485 35.960 ;
      LAYER met4 ;
        RECT 17.165 35.640 17.485 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 35.200 17.485 35.520 ;
      LAYER met4 ;
        RECT 17.165 35.200 17.485 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 34.760 17.485 35.080 ;
      LAYER met4 ;
        RECT 17.165 34.760 17.485 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 50.555 17.020 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 50.135 17.020 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 49.715 17.020 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 37.840 17.080 38.160 ;
      LAYER met4 ;
        RECT 16.760 37.840 17.080 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 37.400 17.080 37.720 ;
      LAYER met4 ;
        RECT 16.760 37.400 17.080 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 36.960 17.080 37.280 ;
      LAYER met4 ;
        RECT 16.760 36.960 17.080 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 36.520 17.080 36.840 ;
      LAYER met4 ;
        RECT 16.760 36.520 17.080 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 36.080 17.080 36.400 ;
      LAYER met4 ;
        RECT 16.760 36.080 17.080 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 35.640 17.080 35.960 ;
      LAYER met4 ;
        RECT 16.760 35.640 17.080 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 35.200 17.080 35.520 ;
      LAYER met4 ;
        RECT 16.760 35.200 17.080 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 34.760 17.080 35.080 ;
      LAYER met4 ;
        RECT 16.760 34.760 17.080 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 50.555 16.615 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 50.135 16.615 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 49.715 16.615 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 37.840 16.675 38.160 ;
      LAYER met4 ;
        RECT 16.355 37.840 16.675 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 37.400 16.675 37.720 ;
      LAYER met4 ;
        RECT 16.355 37.400 16.675 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 36.960 16.675 37.280 ;
      LAYER met4 ;
        RECT 16.355 36.960 16.675 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 36.520 16.675 36.840 ;
      LAYER met4 ;
        RECT 16.355 36.520 16.675 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 36.080 16.675 36.400 ;
      LAYER met4 ;
        RECT 16.355 36.080 16.675 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 35.640 16.675 35.960 ;
      LAYER met4 ;
        RECT 16.355 35.640 16.675 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 35.200 16.675 35.520 ;
      LAYER met4 ;
        RECT 16.355 35.200 16.675 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 34.760 16.675 35.080 ;
      LAYER met4 ;
        RECT 16.355 34.760 16.675 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 50.555 16.210 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 50.135 16.210 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 49.715 16.210 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 37.840 16.270 38.160 ;
      LAYER met4 ;
        RECT 15.950 37.840 16.270 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 37.400 16.270 37.720 ;
      LAYER met4 ;
        RECT 15.950 37.400 16.270 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 36.960 16.270 37.280 ;
      LAYER met4 ;
        RECT 15.950 36.960 16.270 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 36.520 16.270 36.840 ;
      LAYER met4 ;
        RECT 15.950 36.520 16.270 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 36.080 16.270 36.400 ;
      LAYER met4 ;
        RECT 15.950 36.080 16.270 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 35.640 16.270 35.960 ;
      LAYER met4 ;
        RECT 15.950 35.640 16.270 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 35.200 16.270 35.520 ;
      LAYER met4 ;
        RECT 15.950 35.200 16.270 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 34.760 16.270 35.080 ;
      LAYER met4 ;
        RECT 15.950 34.760 16.270 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 50.555 15.805 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 50.135 15.805 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 49.715 15.805 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 37.840 15.865 38.160 ;
      LAYER met4 ;
        RECT 15.545 37.840 15.865 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 37.400 15.865 37.720 ;
      LAYER met4 ;
        RECT 15.545 37.400 15.865 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 36.960 15.865 37.280 ;
      LAYER met4 ;
        RECT 15.545 36.960 15.865 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 36.520 15.865 36.840 ;
      LAYER met4 ;
        RECT 15.545 36.520 15.865 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 36.080 15.865 36.400 ;
      LAYER met4 ;
        RECT 15.545 36.080 15.865 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 35.640 15.865 35.960 ;
      LAYER met4 ;
        RECT 15.545 35.640 15.865 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 35.200 15.865 35.520 ;
      LAYER met4 ;
        RECT 15.545 35.200 15.865 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 34.760 15.865 35.080 ;
      LAYER met4 ;
        RECT 15.545 34.760 15.865 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 50.555 15.400 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 50.135 15.400 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 49.715 15.400 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 37.840 15.460 38.160 ;
      LAYER met4 ;
        RECT 15.140 37.840 15.460 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 37.400 15.460 37.720 ;
      LAYER met4 ;
        RECT 15.140 37.400 15.460 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 36.960 15.460 37.280 ;
      LAYER met4 ;
        RECT 15.140 36.960 15.460 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 36.520 15.460 36.840 ;
      LAYER met4 ;
        RECT 15.140 36.520 15.460 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 36.080 15.460 36.400 ;
      LAYER met4 ;
        RECT 15.140 36.080 15.460 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 35.640 15.460 35.960 ;
      LAYER met4 ;
        RECT 15.140 35.640 15.460 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 35.200 15.460 35.520 ;
      LAYER met4 ;
        RECT 15.140 35.200 15.460 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 34.760 15.460 35.080 ;
      LAYER met4 ;
        RECT 15.140 34.760 15.460 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 50.555 14.995 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 50.135 14.995 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 49.715 14.995 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 37.840 15.055 38.160 ;
      LAYER met4 ;
        RECT 14.735 37.840 15.055 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 37.400 15.055 37.720 ;
      LAYER met4 ;
        RECT 14.735 37.400 15.055 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 36.960 15.055 37.280 ;
      LAYER met4 ;
        RECT 14.735 36.960 15.055 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 36.520 15.055 36.840 ;
      LAYER met4 ;
        RECT 14.735 36.520 15.055 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 36.080 15.055 36.400 ;
      LAYER met4 ;
        RECT 14.735 36.080 15.055 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 35.640 15.055 35.960 ;
      LAYER met4 ;
        RECT 14.735 35.640 15.055 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 35.200 15.055 35.520 ;
      LAYER met4 ;
        RECT 14.735 35.200 15.055 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 34.760 15.055 35.080 ;
      LAYER met4 ;
        RECT 14.735 34.760 15.055 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 50.555 14.590 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 50.135 14.590 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 49.715 14.590 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 37.840 14.650 38.160 ;
      LAYER met4 ;
        RECT 14.330 37.840 14.650 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 37.400 14.650 37.720 ;
      LAYER met4 ;
        RECT 14.330 37.400 14.650 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 36.960 14.650 37.280 ;
      LAYER met4 ;
        RECT 14.330 36.960 14.650 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 36.520 14.650 36.840 ;
      LAYER met4 ;
        RECT 14.330 36.520 14.650 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 36.080 14.650 36.400 ;
      LAYER met4 ;
        RECT 14.330 36.080 14.650 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 35.640 14.650 35.960 ;
      LAYER met4 ;
        RECT 14.330 35.640 14.650 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 35.200 14.650 35.520 ;
      LAYER met4 ;
        RECT 14.330 35.200 14.650 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 34.760 14.650 35.080 ;
      LAYER met4 ;
        RECT 14.330 34.760 14.650 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 50.555 14.185 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 50.135 14.185 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 49.715 14.185 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 37.840 14.245 38.160 ;
      LAYER met4 ;
        RECT 13.925 37.840 14.245 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 37.400 14.245 37.720 ;
      LAYER met4 ;
        RECT 13.925 37.400 14.245 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 36.960 14.245 37.280 ;
      LAYER met4 ;
        RECT 13.925 36.960 14.245 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 36.520 14.245 36.840 ;
      LAYER met4 ;
        RECT 13.925 36.520 14.245 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 36.080 14.245 36.400 ;
      LAYER met4 ;
        RECT 13.925 36.080 14.245 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 35.640 14.245 35.960 ;
      LAYER met4 ;
        RECT 13.925 35.640 14.245 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 35.200 14.245 35.520 ;
      LAYER met4 ;
        RECT 13.925 35.200 14.245 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 34.760 14.245 35.080 ;
      LAYER met4 ;
        RECT 13.925 34.760 14.245 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 50.555 13.780 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 50.135 13.780 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 49.715 13.780 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 37.840 13.840 38.160 ;
      LAYER met4 ;
        RECT 13.520 37.840 13.840 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 37.400 13.840 37.720 ;
      LAYER met4 ;
        RECT 13.520 37.400 13.840 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 36.960 13.840 37.280 ;
      LAYER met4 ;
        RECT 13.520 36.960 13.840 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 36.520 13.840 36.840 ;
      LAYER met4 ;
        RECT 13.520 36.520 13.840 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 36.080 13.840 36.400 ;
      LAYER met4 ;
        RECT 13.520 36.080 13.840 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 35.640 13.840 35.960 ;
      LAYER met4 ;
        RECT 13.520 35.640 13.840 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 35.200 13.840 35.520 ;
      LAYER met4 ;
        RECT 13.520 35.200 13.840 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 34.760 13.840 35.080 ;
      LAYER met4 ;
        RECT 13.520 34.760 13.840 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 50.555 13.375 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 50.135 13.375 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 49.715 13.375 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 37.840 13.435 38.160 ;
      LAYER met4 ;
        RECT 13.115 37.840 13.435 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 37.400 13.435 37.720 ;
      LAYER met4 ;
        RECT 13.115 37.400 13.435 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 36.960 13.435 37.280 ;
      LAYER met4 ;
        RECT 13.115 36.960 13.435 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 36.520 13.435 36.840 ;
      LAYER met4 ;
        RECT 13.115 36.520 13.435 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 36.080 13.435 36.400 ;
      LAYER met4 ;
        RECT 13.115 36.080 13.435 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 35.640 13.435 35.960 ;
      LAYER met4 ;
        RECT 13.115 35.640 13.435 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 35.200 13.435 35.520 ;
      LAYER met4 ;
        RECT 13.115 35.200 13.435 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 34.760 13.435 35.080 ;
      LAYER met4 ;
        RECT 13.115 34.760 13.435 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 50.555 12.970 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 50.135 12.970 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 49.715 12.970 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 37.840 13.030 38.160 ;
      LAYER met4 ;
        RECT 12.710 37.840 13.030 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 37.400 13.030 37.720 ;
      LAYER met4 ;
        RECT 12.710 37.400 13.030 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 36.960 13.030 37.280 ;
      LAYER met4 ;
        RECT 12.710 36.960 13.030 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 36.520 13.030 36.840 ;
      LAYER met4 ;
        RECT 12.710 36.520 13.030 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 36.080 13.030 36.400 ;
      LAYER met4 ;
        RECT 12.710 36.080 13.030 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 35.640 13.030 35.960 ;
      LAYER met4 ;
        RECT 12.710 35.640 13.030 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 35.200 13.030 35.520 ;
      LAYER met4 ;
        RECT 12.710 35.200 13.030 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 34.760 13.030 35.080 ;
      LAYER met4 ;
        RECT 12.710 34.760 13.030 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 50.555 12.565 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 50.135 12.565 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 49.715 12.565 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 37.840 12.625 38.160 ;
      LAYER met4 ;
        RECT 12.305 37.840 12.625 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 37.400 12.625 37.720 ;
      LAYER met4 ;
        RECT 12.305 37.400 12.625 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 36.960 12.625 37.280 ;
      LAYER met4 ;
        RECT 12.305 36.960 12.625 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 36.520 12.625 36.840 ;
      LAYER met4 ;
        RECT 12.305 36.520 12.625 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 36.080 12.625 36.400 ;
      LAYER met4 ;
        RECT 12.305 36.080 12.625 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 35.640 12.625 35.960 ;
      LAYER met4 ;
        RECT 12.305 35.640 12.625 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 35.200 12.625 35.520 ;
      LAYER met4 ;
        RECT 12.305 35.200 12.625 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 34.760 12.625 35.080 ;
      LAYER met4 ;
        RECT 12.305 34.760 12.625 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 50.555 12.160 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 50.135 12.160 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 49.715 12.160 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 37.840 12.220 38.160 ;
      LAYER met4 ;
        RECT 11.900 37.840 12.220 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 37.400 12.220 37.720 ;
      LAYER met4 ;
        RECT 11.900 37.400 12.220 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 36.960 12.220 37.280 ;
      LAYER met4 ;
        RECT 11.900 36.960 12.220 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 36.520 12.220 36.840 ;
      LAYER met4 ;
        RECT 11.900 36.520 12.220 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 36.080 12.220 36.400 ;
      LAYER met4 ;
        RECT 11.900 36.080 12.220 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 35.640 12.220 35.960 ;
      LAYER met4 ;
        RECT 11.900 35.640 12.220 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 35.200 12.220 35.520 ;
      LAYER met4 ;
        RECT 11.900 35.200 12.220 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 34.760 12.220 35.080 ;
      LAYER met4 ;
        RECT 11.900 34.760 12.220 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 50.555 11.755 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 50.135 11.755 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 49.715 11.755 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 37.840 11.815 38.160 ;
      LAYER met4 ;
        RECT 11.495 37.840 11.815 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 37.400 11.815 37.720 ;
      LAYER met4 ;
        RECT 11.495 37.400 11.815 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 36.960 11.815 37.280 ;
      LAYER met4 ;
        RECT 11.495 36.960 11.815 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 36.520 11.815 36.840 ;
      LAYER met4 ;
        RECT 11.495 36.520 11.815 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 36.080 11.815 36.400 ;
      LAYER met4 ;
        RECT 11.495 36.080 11.815 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 35.640 11.815 35.960 ;
      LAYER met4 ;
        RECT 11.495 35.640 11.815 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 35.200 11.815 35.520 ;
      LAYER met4 ;
        RECT 11.495 35.200 11.815 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 34.760 11.815 35.080 ;
      LAYER met4 ;
        RECT 11.495 34.760 11.815 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 50.555 11.350 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 50.135 11.350 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 49.715 11.350 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 37.840 11.410 38.160 ;
      LAYER met4 ;
        RECT 11.090 37.840 11.410 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 37.400 11.410 37.720 ;
      LAYER met4 ;
        RECT 11.090 37.400 11.410 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 36.960 11.410 37.280 ;
      LAYER met4 ;
        RECT 11.090 36.960 11.410 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 36.520 11.410 36.840 ;
      LAYER met4 ;
        RECT 11.090 36.520 11.410 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 36.080 11.410 36.400 ;
      LAYER met4 ;
        RECT 11.090 36.080 11.410 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 35.640 11.410 35.960 ;
      LAYER met4 ;
        RECT 11.090 35.640 11.410 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 35.200 11.410 35.520 ;
      LAYER met4 ;
        RECT 11.090 35.200 11.410 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 34.760 11.410 35.080 ;
      LAYER met4 ;
        RECT 11.090 34.760 11.410 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 50.555 10.945 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 50.135 10.945 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 49.715 10.945 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 37.840 11.005 38.160 ;
      LAYER met4 ;
        RECT 10.685 37.840 11.005 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 37.400 11.005 37.720 ;
      LAYER met4 ;
        RECT 10.685 37.400 11.005 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 36.960 11.005 37.280 ;
      LAYER met4 ;
        RECT 10.685 36.960 11.005 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 36.520 11.005 36.840 ;
      LAYER met4 ;
        RECT 10.685 36.520 11.005 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 36.080 11.005 36.400 ;
      LAYER met4 ;
        RECT 10.685 36.080 11.005 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 35.640 11.005 35.960 ;
      LAYER met4 ;
        RECT 10.685 35.640 11.005 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 35.200 11.005 35.520 ;
      LAYER met4 ;
        RECT 10.685 35.200 11.005 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 34.760 11.005 35.080 ;
      LAYER met4 ;
        RECT 10.685 34.760 11.005 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 50.555 10.540 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 50.135 10.540 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 49.715 10.540 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 37.840 10.600 38.160 ;
      LAYER met4 ;
        RECT 10.280 37.840 10.600 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 37.400 10.600 37.720 ;
      LAYER met4 ;
        RECT 10.280 37.400 10.600 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 36.960 10.600 37.280 ;
      LAYER met4 ;
        RECT 10.280 36.960 10.600 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 36.520 10.600 36.840 ;
      LAYER met4 ;
        RECT 10.280 36.520 10.600 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 36.080 10.600 36.400 ;
      LAYER met4 ;
        RECT 10.280 36.080 10.600 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 35.640 10.600 35.960 ;
      LAYER met4 ;
        RECT 10.280 35.640 10.600 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 35.200 10.600 35.520 ;
      LAYER met4 ;
        RECT 10.280 35.200 10.600 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 34.760 10.600 35.080 ;
      LAYER met4 ;
        RECT 10.280 34.760 10.600 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 50.555 10.135 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 50.135 10.135 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 49.715 10.135 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 37.840 10.195 38.160 ;
      LAYER met4 ;
        RECT 9.875 37.840 10.195 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 37.400 10.195 37.720 ;
      LAYER met4 ;
        RECT 9.875 37.400 10.195 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 36.960 10.195 37.280 ;
      LAYER met4 ;
        RECT 9.875 36.960 10.195 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 36.520 10.195 36.840 ;
      LAYER met4 ;
        RECT 9.875 36.520 10.195 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 36.080 10.195 36.400 ;
      LAYER met4 ;
        RECT 9.875 36.080 10.195 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 35.640 10.195 35.960 ;
      LAYER met4 ;
        RECT 9.875 35.640 10.195 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 35.200 10.195 35.520 ;
      LAYER met4 ;
        RECT 9.875 35.200 10.195 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 34.760 10.195 35.080 ;
      LAYER met4 ;
        RECT 9.875 34.760 10.195 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 50.555 9.730 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 50.135 9.730 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 49.715 9.730 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 37.840 9.790 38.160 ;
      LAYER met4 ;
        RECT 9.470 37.840 9.790 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 37.400 9.790 37.720 ;
      LAYER met4 ;
        RECT 9.470 37.400 9.790 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 36.960 9.790 37.280 ;
      LAYER met4 ;
        RECT 9.470 36.960 9.790 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 36.520 9.790 36.840 ;
      LAYER met4 ;
        RECT 9.470 36.520 9.790 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 36.080 9.790 36.400 ;
      LAYER met4 ;
        RECT 9.470 36.080 9.790 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 35.640 9.790 35.960 ;
      LAYER met4 ;
        RECT 9.470 35.640 9.790 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 35.200 9.790 35.520 ;
      LAYER met4 ;
        RECT 9.470 35.200 9.790 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 34.760 9.790 35.080 ;
      LAYER met4 ;
        RECT 9.470 34.760 9.790 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 50.555 9.325 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 50.135 9.325 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 49.715 9.325 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 37.840 9.385 38.160 ;
      LAYER met4 ;
        RECT 9.065 37.840 9.385 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 37.400 9.385 37.720 ;
      LAYER met4 ;
        RECT 9.065 37.400 9.385 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 36.960 9.385 37.280 ;
      LAYER met4 ;
        RECT 9.065 36.960 9.385 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 36.520 9.385 36.840 ;
      LAYER met4 ;
        RECT 9.065 36.520 9.385 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 36.080 9.385 36.400 ;
      LAYER met4 ;
        RECT 9.065 36.080 9.385 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 35.640 9.385 35.960 ;
      LAYER met4 ;
        RECT 9.065 35.640 9.385 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 35.200 9.385 35.520 ;
      LAYER met4 ;
        RECT 9.065 35.200 9.385 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 34.760 9.385 35.080 ;
      LAYER met4 ;
        RECT 9.065 34.760 9.385 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 50.555 8.920 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 50.135 8.920 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 49.715 8.920 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 37.840 8.980 38.160 ;
      LAYER met4 ;
        RECT 8.660 37.840 8.980 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 37.400 8.980 37.720 ;
      LAYER met4 ;
        RECT 8.660 37.400 8.980 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 36.960 8.980 37.280 ;
      LAYER met4 ;
        RECT 8.660 36.960 8.980 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 36.520 8.980 36.840 ;
      LAYER met4 ;
        RECT 8.660 36.520 8.980 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 36.080 8.980 36.400 ;
      LAYER met4 ;
        RECT 8.660 36.080 8.980 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 35.640 8.980 35.960 ;
      LAYER met4 ;
        RECT 8.660 35.640 8.980 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 35.200 8.980 35.520 ;
      LAYER met4 ;
        RECT 8.660 35.200 8.980 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 34.760 8.980 35.080 ;
      LAYER met4 ;
        RECT 8.660 34.760 8.980 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 50.555 8.515 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 50.135 8.515 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 49.715 8.515 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 37.840 8.575 38.160 ;
      LAYER met4 ;
        RECT 8.255 37.840 8.575 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 37.400 8.575 37.720 ;
      LAYER met4 ;
        RECT 8.255 37.400 8.575 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 36.960 8.575 37.280 ;
      LAYER met4 ;
        RECT 8.255 36.960 8.575 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 36.520 8.575 36.840 ;
      LAYER met4 ;
        RECT 8.255 36.520 8.575 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 36.080 8.575 36.400 ;
      LAYER met4 ;
        RECT 8.255 36.080 8.575 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 35.640 8.575 35.960 ;
      LAYER met4 ;
        RECT 8.255 35.640 8.575 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 35.200 8.575 35.520 ;
      LAYER met4 ;
        RECT 8.255 35.200 8.575 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 34.760 8.575 35.080 ;
      LAYER met4 ;
        RECT 8.255 34.760 8.575 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 50.555 8.110 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 50.135 8.110 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 49.715 8.110 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 37.840 8.170 38.160 ;
      LAYER met4 ;
        RECT 7.850 37.840 8.170 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 37.400 8.170 37.720 ;
      LAYER met4 ;
        RECT 7.850 37.400 8.170 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 36.960 8.170 37.280 ;
      LAYER met4 ;
        RECT 7.850 36.960 8.170 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 36.520 8.170 36.840 ;
      LAYER met4 ;
        RECT 7.850 36.520 8.170 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 36.080 8.170 36.400 ;
      LAYER met4 ;
        RECT 7.850 36.080 8.170 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 35.640 8.170 35.960 ;
      LAYER met4 ;
        RECT 7.850 35.640 8.170 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 35.200 8.170 35.520 ;
      LAYER met4 ;
        RECT 7.850 35.200 8.170 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 34.760 8.170 35.080 ;
      LAYER met4 ;
        RECT 7.850 34.760 8.170 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 50.555 7.705 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 50.135 7.705 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 49.715 7.705 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 37.840 7.765 38.160 ;
      LAYER met4 ;
        RECT 7.445 37.840 7.765 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 37.400 7.765 37.720 ;
      LAYER met4 ;
        RECT 7.445 37.400 7.765 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 36.960 7.765 37.280 ;
      LAYER met4 ;
        RECT 7.445 36.960 7.765 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 36.520 7.765 36.840 ;
      LAYER met4 ;
        RECT 7.445 36.520 7.765 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 36.080 7.765 36.400 ;
      LAYER met4 ;
        RECT 7.445 36.080 7.765 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 35.640 7.765 35.960 ;
      LAYER met4 ;
        RECT 7.445 35.640 7.765 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 35.200 7.765 35.520 ;
      LAYER met4 ;
        RECT 7.445 35.200 7.765 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 34.760 7.765 35.080 ;
      LAYER met4 ;
        RECT 7.445 34.760 7.765 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 50.555 7.300 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 50.135 7.300 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 49.715 7.300 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 37.840 7.360 38.160 ;
      LAYER met4 ;
        RECT 7.040 37.840 7.360 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 37.400 7.360 37.720 ;
      LAYER met4 ;
        RECT 7.040 37.400 7.360 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 36.960 7.360 37.280 ;
      LAYER met4 ;
        RECT 7.040 36.960 7.360 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 36.520 7.360 36.840 ;
      LAYER met4 ;
        RECT 7.040 36.520 7.360 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 36.080 7.360 36.400 ;
      LAYER met4 ;
        RECT 7.040 36.080 7.360 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 35.640 7.360 35.960 ;
      LAYER met4 ;
        RECT 7.040 35.640 7.360 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 35.200 7.360 35.520 ;
      LAYER met4 ;
        RECT 7.040 35.200 7.360 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 34.760 7.360 35.080 ;
      LAYER met4 ;
        RECT 7.040 34.760 7.360 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 50.555 6.895 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 50.135 6.895 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 49.715 6.895 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 37.840 6.955 38.160 ;
      LAYER met4 ;
        RECT 6.635 37.840 6.955 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 37.400 6.955 37.720 ;
      LAYER met4 ;
        RECT 6.635 37.400 6.955 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 36.960 6.955 37.280 ;
      LAYER met4 ;
        RECT 6.635 36.960 6.955 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 36.520 6.955 36.840 ;
      LAYER met4 ;
        RECT 6.635 36.520 6.955 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 36.080 6.955 36.400 ;
      LAYER met4 ;
        RECT 6.635 36.080 6.955 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 35.640 6.955 35.960 ;
      LAYER met4 ;
        RECT 6.635 35.640 6.955 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 35.200 6.955 35.520 ;
      LAYER met4 ;
        RECT 6.635 35.200 6.955 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 34.760 6.955 35.080 ;
      LAYER met4 ;
        RECT 6.635 34.760 6.955 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 50.555 6.490 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 50.135 6.490 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 49.715 6.490 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 37.840 6.550 38.160 ;
      LAYER met4 ;
        RECT 6.230 37.840 6.550 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 37.400 6.550 37.720 ;
      LAYER met4 ;
        RECT 6.230 37.400 6.550 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 36.960 6.550 37.280 ;
      LAYER met4 ;
        RECT 6.230 36.960 6.550 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 36.520 6.550 36.840 ;
      LAYER met4 ;
        RECT 6.230 36.520 6.550 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 36.080 6.550 36.400 ;
      LAYER met4 ;
        RECT 6.230 36.080 6.550 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 35.640 6.550 35.960 ;
      LAYER met4 ;
        RECT 6.230 35.640 6.550 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 35.200 6.550 35.520 ;
      LAYER met4 ;
        RECT 6.230 35.200 6.550 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 34.760 6.550 35.080 ;
      LAYER met4 ;
        RECT 6.230 34.760 6.550 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 50.555 6.085 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 50.135 6.085 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 49.715 6.085 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 37.840 6.145 38.160 ;
      LAYER met4 ;
        RECT 5.825 37.840 6.145 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 37.400 6.145 37.720 ;
      LAYER met4 ;
        RECT 5.825 37.400 6.145 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 36.960 6.145 37.280 ;
      LAYER met4 ;
        RECT 5.825 36.960 6.145 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 36.520 6.145 36.840 ;
      LAYER met4 ;
        RECT 5.825 36.520 6.145 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 36.080 6.145 36.400 ;
      LAYER met4 ;
        RECT 5.825 36.080 6.145 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 35.640 6.145 35.960 ;
      LAYER met4 ;
        RECT 5.825 35.640 6.145 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 35.200 6.145 35.520 ;
      LAYER met4 ;
        RECT 5.825 35.200 6.145 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 34.760 6.145 35.080 ;
      LAYER met4 ;
        RECT 5.825 34.760 6.145 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 50.555 5.680 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 50.135 5.680 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 49.715 5.680 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 37.840 5.740 38.160 ;
      LAYER met4 ;
        RECT 5.420 37.840 5.740 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 37.400 5.740 37.720 ;
      LAYER met4 ;
        RECT 5.420 37.400 5.740 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 36.960 5.740 37.280 ;
      LAYER met4 ;
        RECT 5.420 36.960 5.740 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 36.520 5.740 36.840 ;
      LAYER met4 ;
        RECT 5.420 36.520 5.740 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 36.080 5.740 36.400 ;
      LAYER met4 ;
        RECT 5.420 36.080 5.740 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 35.640 5.740 35.960 ;
      LAYER met4 ;
        RECT 5.420 35.640 5.740 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 35.200 5.740 35.520 ;
      LAYER met4 ;
        RECT 5.420 35.200 5.740 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 34.760 5.740 35.080 ;
      LAYER met4 ;
        RECT 5.420 34.760 5.740 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 50.555 5.275 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 50.135 5.275 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 49.715 5.275 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 37.840 5.335 38.160 ;
      LAYER met4 ;
        RECT 5.015 37.840 5.335 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 37.400 5.335 37.720 ;
      LAYER met4 ;
        RECT 5.015 37.400 5.335 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 36.960 5.335 37.280 ;
      LAYER met4 ;
        RECT 5.015 36.960 5.335 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 36.520 5.335 36.840 ;
      LAYER met4 ;
        RECT 5.015 36.520 5.335 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 36.080 5.335 36.400 ;
      LAYER met4 ;
        RECT 5.015 36.080 5.335 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 35.640 5.335 35.960 ;
      LAYER met4 ;
        RECT 5.015 35.640 5.335 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 35.200 5.335 35.520 ;
      LAYER met4 ;
        RECT 5.015 35.200 5.335 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 34.760 5.335 35.080 ;
      LAYER met4 ;
        RECT 5.015 34.760 5.335 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 50.555 4.870 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 50.135 4.870 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 49.715 4.870 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 37.840 4.930 38.160 ;
      LAYER met4 ;
        RECT 4.610 37.840 4.930 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 37.400 4.930 37.720 ;
      LAYER met4 ;
        RECT 4.610 37.400 4.930 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 36.960 4.930 37.280 ;
      LAYER met4 ;
        RECT 4.610 36.960 4.930 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 36.520 4.930 36.840 ;
      LAYER met4 ;
        RECT 4.610 36.520 4.930 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 36.080 4.930 36.400 ;
      LAYER met4 ;
        RECT 4.610 36.080 4.930 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 35.640 4.930 35.960 ;
      LAYER met4 ;
        RECT 4.610 35.640 4.930 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 35.200 4.930 35.520 ;
      LAYER met4 ;
        RECT 4.610 35.200 4.930 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 34.760 4.930 35.080 ;
      LAYER met4 ;
        RECT 4.610 34.760 4.930 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 50.555 4.465 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 50.135 4.465 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 49.715 4.465 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 37.840 4.525 38.160 ;
      LAYER met4 ;
        RECT 4.205 37.840 4.525 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 37.400 4.525 37.720 ;
      LAYER met4 ;
        RECT 4.205 37.400 4.525 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 36.960 4.525 37.280 ;
      LAYER met4 ;
        RECT 4.205 36.960 4.525 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 36.520 4.525 36.840 ;
      LAYER met4 ;
        RECT 4.205 36.520 4.525 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 36.080 4.525 36.400 ;
      LAYER met4 ;
        RECT 4.205 36.080 4.525 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 35.640 4.525 35.960 ;
      LAYER met4 ;
        RECT 4.205 35.640 4.525 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 35.200 4.525 35.520 ;
      LAYER met4 ;
        RECT 4.205 35.200 4.525 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 34.760 4.525 35.080 ;
      LAYER met4 ;
        RECT 4.205 34.760 4.525 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 50.555 4.060 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 50.135 4.060 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 49.715 4.060 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 37.840 4.120 38.160 ;
      LAYER met4 ;
        RECT 3.800 37.840 4.120 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 37.400 4.120 37.720 ;
      LAYER met4 ;
        RECT 3.800 37.400 4.120 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 36.960 4.120 37.280 ;
      LAYER met4 ;
        RECT 3.800 36.960 4.120 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 36.520 4.120 36.840 ;
      LAYER met4 ;
        RECT 3.800 36.520 4.120 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 36.080 4.120 36.400 ;
      LAYER met4 ;
        RECT 3.800 36.080 4.120 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 35.640 4.120 35.960 ;
      LAYER met4 ;
        RECT 3.800 35.640 4.120 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 35.200 4.120 35.520 ;
      LAYER met4 ;
        RECT 3.800 35.200 4.120 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 34.760 4.120 35.080 ;
      LAYER met4 ;
        RECT 3.800 34.760 4.120 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 50.555 3.655 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 50.135 3.655 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 49.715 3.655 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 37.840 3.715 38.160 ;
      LAYER met4 ;
        RECT 3.395 37.840 3.715 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 37.400 3.715 37.720 ;
      LAYER met4 ;
        RECT 3.395 37.400 3.715 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 36.960 3.715 37.280 ;
      LAYER met4 ;
        RECT 3.395 36.960 3.715 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 36.520 3.715 36.840 ;
      LAYER met4 ;
        RECT 3.395 36.520 3.715 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 36.080 3.715 36.400 ;
      LAYER met4 ;
        RECT 3.395 36.080 3.715 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 35.640 3.715 35.960 ;
      LAYER met4 ;
        RECT 3.395 35.640 3.715 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 35.200 3.715 35.520 ;
      LAYER met4 ;
        RECT 3.395 35.200 3.715 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 34.760 3.715 35.080 ;
      LAYER met4 ;
        RECT 3.395 34.760 3.715 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 50.555 3.250 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 50.135 3.250 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 49.715 3.250 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 37.840 3.310 38.160 ;
      LAYER met4 ;
        RECT 2.990 37.840 3.310 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 37.400 3.310 37.720 ;
      LAYER met4 ;
        RECT 2.990 37.400 3.310 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 36.960 3.310 37.280 ;
      LAYER met4 ;
        RECT 2.990 36.960 3.310 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 36.520 3.310 36.840 ;
      LAYER met4 ;
        RECT 2.990 36.520 3.310 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 36.080 3.310 36.400 ;
      LAYER met4 ;
        RECT 2.990 36.080 3.310 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 35.640 3.310 35.960 ;
      LAYER met4 ;
        RECT 2.990 35.640 3.310 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 35.200 3.310 35.520 ;
      LAYER met4 ;
        RECT 2.990 35.200 3.310 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 34.760 3.310 35.080 ;
      LAYER met4 ;
        RECT 2.990 34.760 3.310 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 50.555 2.840 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 50.135 2.840 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 49.715 2.840 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 37.840 2.900 38.160 ;
      LAYER met4 ;
        RECT 2.580 37.840 2.900 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 37.400 2.900 37.720 ;
      LAYER met4 ;
        RECT 2.580 37.400 2.900 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 36.960 2.900 37.280 ;
      LAYER met4 ;
        RECT 2.580 36.960 2.900 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 36.520 2.900 36.840 ;
      LAYER met4 ;
        RECT 2.580 36.520 2.900 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 36.080 2.900 36.400 ;
      LAYER met4 ;
        RECT 2.580 36.080 2.900 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 35.640 2.900 35.960 ;
      LAYER met4 ;
        RECT 2.580 35.640 2.900 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 35.200 2.900 35.520 ;
      LAYER met4 ;
        RECT 2.580 35.200 2.900 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 34.760 2.900 35.080 ;
      LAYER met4 ;
        RECT 2.580 34.760 2.900 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 50.555 2.430 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 50.135 2.430 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 49.715 2.430 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 37.840 2.490 38.160 ;
      LAYER met4 ;
        RECT 2.170 37.840 2.490 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 37.400 2.490 37.720 ;
      LAYER met4 ;
        RECT 2.170 37.400 2.490 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 36.960 2.490 37.280 ;
      LAYER met4 ;
        RECT 2.170 36.960 2.490 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 36.520 2.490 36.840 ;
      LAYER met4 ;
        RECT 2.170 36.520 2.490 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 36.080 2.490 36.400 ;
      LAYER met4 ;
        RECT 2.170 36.080 2.490 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 35.640 2.490 35.960 ;
      LAYER met4 ;
        RECT 2.170 35.640 2.490 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 35.200 2.490 35.520 ;
      LAYER met4 ;
        RECT 2.170 35.200 2.490 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 34.760 2.490 35.080 ;
      LAYER met4 ;
        RECT 2.170 34.760 2.490 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 50.555 2.020 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 50.135 2.020 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 49.715 2.020 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 37.840 2.080 38.160 ;
      LAYER met4 ;
        RECT 1.760 37.840 2.080 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 37.400 2.080 37.720 ;
      LAYER met4 ;
        RECT 1.760 37.400 2.080 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 36.960 2.080 37.280 ;
      LAYER met4 ;
        RECT 1.760 36.960 2.080 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 36.520 2.080 36.840 ;
      LAYER met4 ;
        RECT 1.760 36.520 2.080 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 36.080 2.080 36.400 ;
      LAYER met4 ;
        RECT 1.760 36.080 2.080 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 35.640 2.080 35.960 ;
      LAYER met4 ;
        RECT 1.760 35.640 2.080 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 35.200 2.080 35.520 ;
      LAYER met4 ;
        RECT 1.760 35.200 2.080 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 34.760 2.080 35.080 ;
      LAYER met4 ;
        RECT 1.760 34.760 2.080 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 50.555 1.610 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 50.135 1.610 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 49.715 1.610 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 37.840 1.670 38.160 ;
      LAYER met4 ;
        RECT 1.350 37.840 1.670 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 37.400 1.670 37.720 ;
      LAYER met4 ;
        RECT 1.350 37.400 1.670 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 36.960 1.670 37.280 ;
      LAYER met4 ;
        RECT 1.350 36.960 1.670 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 36.520 1.670 36.840 ;
      LAYER met4 ;
        RECT 1.350 36.520 1.670 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 36.080 1.670 36.400 ;
      LAYER met4 ;
        RECT 1.350 36.080 1.670 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 35.640 1.670 35.960 ;
      LAYER met4 ;
        RECT 1.350 35.640 1.670 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 35.200 1.670 35.520 ;
      LAYER met4 ;
        RECT 1.350 35.200 1.670 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 34.760 1.670 35.080 ;
      LAYER met4 ;
        RECT 1.350 34.760 1.670 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 50.555 1.200 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 50.135 1.200 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 49.715 1.200 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 37.840 1.260 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 37.400 1.260 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 36.960 1.260 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 36.520 1.260 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 36.080 1.260 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 35.640 1.260 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 35.200 1.260 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 34.760 1.260 35.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 50.555 0.790 50.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 50.135 0.790 50.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 49.715 0.790 49.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 37.840 0.850 38.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 37.400 0.850 37.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 36.960 0.850 37.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 36.520 0.850 36.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 36.080 0.850 36.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 35.640 0.850 35.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 35.200 0.850 35.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 34.760 0.850 35.080 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
  END VSSIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
  END VDDIO
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  OBS
      LAYER met3 ;
        RECT 0.500 34.740 24.400 38.180 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 94.585 75.000 172.185 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__overlay_vssa_lvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vssd_hvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vssd_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
  END VCCD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
  END VDDA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 41.590 74.290 46.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 45.960 74.200 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 45.530 74.200 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 45.100 74.200 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 44.670 74.200 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 44.240 74.200 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 43.810 74.200 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 43.380 74.200 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 42.950 74.200 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 42.520 74.200 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 42.090 74.200 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 41.660 74.200 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 45.960 73.795 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 45.530 73.795 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 45.100 73.795 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 44.670 73.795 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 44.240 73.795 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 43.810 73.795 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 43.380 73.795 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 42.950 73.795 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 42.520 73.795 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 42.090 73.795 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 41.660 73.795 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 45.960 73.390 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 45.530 73.390 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 45.100 73.390 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 44.670 73.390 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 44.240 73.390 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 43.810 73.390 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 43.380 73.390 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 42.950 73.390 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 42.520 73.390 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 42.090 73.390 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 41.660 73.390 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 45.960 72.985 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 45.530 72.985 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 45.100 72.985 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 44.670 72.985 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 44.240 72.985 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 43.810 72.985 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 43.380 72.985 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 42.950 72.985 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 42.520 72.985 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 42.090 72.985 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 41.660 72.985 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 45.960 72.580 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 45.530 72.580 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 45.100 72.580 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 44.670 72.580 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 44.240 72.580 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 43.810 72.580 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 43.380 72.580 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 42.950 72.580 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 42.520 72.580 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 42.090 72.580 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 41.660 72.580 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 45.960 72.175 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 45.530 72.175 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 45.100 72.175 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 44.670 72.175 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 44.240 72.175 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 43.810 72.175 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 43.380 72.175 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 42.950 72.175 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 42.520 72.175 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 42.090 72.175 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 41.660 72.175 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 45.960 71.770 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 45.530 71.770 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 45.100 71.770 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 44.670 71.770 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 44.240 71.770 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 43.810 71.770 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 43.380 71.770 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 42.950 71.770 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 42.520 71.770 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 42.090 71.770 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 41.660 71.770 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 45.960 71.365 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 45.530 71.365 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 45.100 71.365 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 44.670 71.365 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 44.240 71.365 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 43.810 71.365 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 43.380 71.365 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 42.950 71.365 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 42.520 71.365 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 42.090 71.365 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 41.660 71.365 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 45.960 70.960 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 45.530 70.960 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 45.100 70.960 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 44.670 70.960 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 44.240 70.960 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 43.810 70.960 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 43.380 70.960 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 42.950 70.960 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 42.520 70.960 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 42.090 70.960 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 41.660 70.960 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 45.960 70.555 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 45.530 70.555 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 45.100 70.555 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 44.670 70.555 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 44.240 70.555 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 43.810 70.555 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 43.380 70.555 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 42.950 70.555 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 42.520 70.555 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 42.090 70.555 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 41.660 70.555 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 45.960 70.150 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 45.530 70.150 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 45.100 70.150 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 44.670 70.150 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 44.240 70.150 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 43.810 70.150 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 43.380 70.150 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 42.950 70.150 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 42.520 70.150 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 42.090 70.150 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 41.660 70.150 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 45.960 69.745 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 45.530 69.745 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 45.100 69.745 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 44.670 69.745 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 44.240 69.745 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 43.810 69.745 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 43.380 69.745 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 42.950 69.745 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 42.520 69.745 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 42.090 69.745 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 41.660 69.745 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 45.960 69.340 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 45.530 69.340 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 45.100 69.340 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 44.670 69.340 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 44.240 69.340 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 43.810 69.340 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 43.380 69.340 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 42.950 69.340 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 42.520 69.340 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 42.090 69.340 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 41.660 69.340 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 45.960 68.935 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 45.530 68.935 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 45.100 68.935 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 44.670 68.935 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 44.240 68.935 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 43.810 68.935 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 43.380 68.935 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 42.950 68.935 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 42.520 68.935 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 42.090 68.935 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 41.660 68.935 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 45.960 68.530 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 45.530 68.530 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 45.100 68.530 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 44.670 68.530 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 44.240 68.530 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 43.810 68.530 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 43.380 68.530 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 42.950 68.530 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 42.520 68.530 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 42.090 68.530 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 41.660 68.530 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 45.960 68.125 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 45.530 68.125 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 45.100 68.125 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 44.670 68.125 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 44.240 68.125 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 43.810 68.125 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 43.380 68.125 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 42.950 68.125 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 42.520 68.125 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 42.090 68.125 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 41.660 68.125 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 45.960 67.720 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 45.530 67.720 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 45.100 67.720 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 44.670 67.720 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 44.240 67.720 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 43.810 67.720 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 43.380 67.720 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 42.950 67.720 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 42.520 67.720 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 42.090 67.720 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 41.660 67.720 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 45.960 67.315 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 45.530 67.315 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 45.100 67.315 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 44.670 67.315 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 44.240 67.315 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 43.810 67.315 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 43.380 67.315 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 42.950 67.315 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 42.520 67.315 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 42.090 67.315 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 41.660 67.315 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 45.960 66.910 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 45.530 66.910 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 45.100 66.910 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 44.670 66.910 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 44.240 66.910 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 43.810 66.910 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 43.380 66.910 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 42.950 66.910 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 42.520 66.910 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 42.090 66.910 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 41.660 66.910 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 45.960 66.505 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 45.530 66.505 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 45.100 66.505 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 44.670 66.505 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 44.240 66.505 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 43.810 66.505 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 43.380 66.505 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 42.950 66.505 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 42.520 66.505 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 42.090 66.505 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 41.660 66.505 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 45.960 66.100 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 45.530 66.100 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 45.100 66.100 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 44.670 66.100 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 44.240 66.100 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 43.810 66.100 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 43.380 66.100 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 42.950 66.100 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 42.520 66.100 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 42.090 66.100 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 41.660 66.100 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 45.960 65.695 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 45.530 65.695 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 45.100 65.695 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 44.670 65.695 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 44.240 65.695 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 43.810 65.695 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 43.380 65.695 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 42.950 65.695 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 42.520 65.695 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 42.090 65.695 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 41.660 65.695 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 45.960 65.290 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 45.530 65.290 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 45.100 65.290 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 44.670 65.290 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 44.240 65.290 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 43.810 65.290 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 43.380 65.290 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 42.950 65.290 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 42.520 65.290 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 42.090 65.290 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 41.660 65.290 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 45.960 64.885 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 45.530 64.885 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 45.100 64.885 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 44.670 64.885 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 44.240 64.885 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 43.810 64.885 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 43.380 64.885 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 42.950 64.885 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 42.520 64.885 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 42.090 64.885 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 41.660 64.885 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 45.960 64.480 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 45.530 64.480 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 45.100 64.480 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 44.670 64.480 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 44.240 64.480 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 43.810 64.480 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 43.380 64.480 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 42.950 64.480 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 42.520 64.480 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 42.090 64.480 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 41.660 64.480 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 45.960 64.075 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 45.530 64.075 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 45.100 64.075 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 44.670 64.075 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 44.240 64.075 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 43.810 64.075 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 43.380 64.075 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 42.950 64.075 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 42.520 64.075 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 42.090 64.075 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 41.660 64.075 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 45.960 63.670 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 45.530 63.670 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 45.100 63.670 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 44.670 63.670 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 44.240 63.670 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 43.810 63.670 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 43.380 63.670 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 42.950 63.670 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 42.520 63.670 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 42.090 63.670 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 41.660 63.670 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 45.960 63.265 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 45.530 63.265 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 45.100 63.265 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 44.670 63.265 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 44.240 63.265 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 43.810 63.265 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 43.380 63.265 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 42.950 63.265 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 42.520 63.265 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 42.090 63.265 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 41.660 63.265 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 45.960 62.860 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 45.530 62.860 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 45.100 62.860 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 44.670 62.860 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 44.240 62.860 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 43.810 62.860 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 43.380 62.860 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 42.950 62.860 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 42.520 62.860 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 42.090 62.860 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 41.660 62.860 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 45.960 62.455 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 45.530 62.455 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 45.100 62.455 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 44.670 62.455 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 44.240 62.455 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 43.810 62.455 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 43.380 62.455 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 42.950 62.455 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 42.520 62.455 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 42.090 62.455 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 41.660 62.455 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 45.960 62.050 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 45.530 62.050 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 45.100 62.050 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 44.670 62.050 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 44.240 62.050 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 43.810 62.050 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 43.380 62.050 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 42.950 62.050 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 42.520 62.050 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 42.090 62.050 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 41.660 62.050 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 45.960 61.645 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 45.530 61.645 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 45.100 61.645 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 44.670 61.645 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 44.240 61.645 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 43.810 61.645 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 43.380 61.645 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 42.950 61.645 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 42.520 61.645 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 42.090 61.645 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 41.660 61.645 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 45.960 61.240 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 45.530 61.240 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 45.100 61.240 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 44.670 61.240 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 44.240 61.240 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 43.810 61.240 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 43.380 61.240 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 42.950 61.240 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 42.520 61.240 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 42.090 61.240 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 41.660 61.240 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 45.960 60.835 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 45.530 60.835 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 45.100 60.835 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 44.670 60.835 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 44.240 60.835 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 43.810 60.835 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 43.380 60.835 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 42.950 60.835 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 42.520 60.835 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 42.090 60.835 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 41.660 60.835 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 45.960 60.430 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 45.530 60.430 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 45.100 60.430 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 44.670 60.430 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 44.240 60.430 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 43.810 60.430 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 43.380 60.430 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 42.950 60.430 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 42.520 60.430 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 42.090 60.430 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 41.660 60.430 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 45.960 60.025 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 45.530 60.025 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 45.100 60.025 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 44.670 60.025 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 44.240 60.025 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 43.810 60.025 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 43.380 60.025 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 42.950 60.025 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 42.520 60.025 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 42.090 60.025 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 41.660 60.025 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 45.960 59.620 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 45.530 59.620 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 45.100 59.620 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 44.670 59.620 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 44.240 59.620 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 43.810 59.620 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 43.380 59.620 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 42.950 59.620 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 42.520 59.620 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 42.090 59.620 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 41.660 59.620 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 45.960 59.215 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 45.530 59.215 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 45.100 59.215 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 44.670 59.215 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 44.240 59.215 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 43.810 59.215 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 43.380 59.215 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 42.950 59.215 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 42.520 59.215 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 42.090 59.215 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 41.660 59.215 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 45.960 58.810 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 45.530 58.810 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 45.100 58.810 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 44.670 58.810 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 44.240 58.810 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 43.810 58.810 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 43.380 58.810 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 42.950 58.810 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 42.520 58.810 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 42.090 58.810 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 41.660 58.810 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 45.960 58.405 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 45.530 58.405 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 45.100 58.405 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 44.670 58.405 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 44.240 58.405 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 43.810 58.405 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 43.380 58.405 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 42.950 58.405 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 42.520 58.405 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 42.090 58.405 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 41.660 58.405 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 45.960 58.000 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 45.530 58.000 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 45.100 58.000 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 44.670 58.000 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 44.240 58.000 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 43.810 58.000 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 43.380 58.000 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 42.950 58.000 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 42.520 58.000 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 42.090 58.000 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 41.660 58.000 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 45.960 57.595 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 45.530 57.595 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 45.100 57.595 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 44.670 57.595 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 44.240 57.595 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 43.810 57.595 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 43.380 57.595 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 42.950 57.595 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 42.520 57.595 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 42.090 57.595 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 41.660 57.595 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 45.960 57.190 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 45.530 57.190 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 45.100 57.190 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 44.670 57.190 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 44.240 57.190 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 43.810 57.190 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 43.380 57.190 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 42.950 57.190 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 42.520 57.190 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 42.090 57.190 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 41.660 57.190 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 45.960 56.785 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 45.530 56.785 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 45.100 56.785 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 44.670 56.785 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 44.240 56.785 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 43.810 56.785 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 43.380 56.785 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 42.950 56.785 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 42.520 56.785 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 42.090 56.785 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 41.660 56.785 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 45.960 56.380 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 45.530 56.380 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 45.100 56.380 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 44.670 56.380 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 44.240 56.380 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 43.810 56.380 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 43.380 56.380 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 42.950 56.380 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 42.520 56.380 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 42.090 56.380 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 41.660 56.380 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 45.960 55.975 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 45.530 55.975 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 45.100 55.975 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 44.670 55.975 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 44.240 55.975 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 43.810 55.975 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 43.380 55.975 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 42.950 55.975 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 42.520 55.975 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 42.090 55.975 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 41.660 55.975 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 45.960 55.570 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 45.530 55.570 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 45.100 55.570 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 44.670 55.570 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 44.240 55.570 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 43.810 55.570 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 43.380 55.570 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 42.950 55.570 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 42.520 55.570 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 42.090 55.570 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 41.660 55.570 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 45.960 55.165 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 45.530 55.165 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 45.100 55.165 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 44.670 55.165 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 44.240 55.165 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 43.810 55.165 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 43.380 55.165 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 42.950 55.165 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 42.520 55.165 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 42.090 55.165 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 41.660 55.165 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 45.960 54.760 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 45.530 54.760 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 45.100 54.760 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 44.670 54.760 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 44.240 54.760 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 43.810 54.760 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 43.380 54.760 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 42.950 54.760 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 42.520 54.760 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 42.090 54.760 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 41.660 54.760 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 45.960 54.355 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 45.530 54.355 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 45.100 54.355 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 44.670 54.355 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 44.240 54.355 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 43.810 54.355 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 43.380 54.355 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 42.950 54.355 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 42.520 54.355 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 42.090 54.355 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 41.660 54.355 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 45.960 53.950 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 45.530 53.950 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 45.100 53.950 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 44.670 53.950 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 44.240 53.950 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 43.810 53.950 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 43.380 53.950 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 42.950 53.950 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 42.520 53.950 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 42.090 53.950 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 41.660 53.950 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 45.960 53.545 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 45.530 53.545 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 45.100 53.545 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 44.670 53.545 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 44.240 53.545 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 43.810 53.545 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 43.380 53.545 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 42.950 53.545 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 42.520 53.545 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 42.090 53.545 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 41.660 53.545 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 45.960 53.140 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 45.530 53.140 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 45.100 53.140 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 44.670 53.140 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 44.240 53.140 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 43.810 53.140 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 43.380 53.140 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 42.950 53.140 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 42.520 53.140 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 42.090 53.140 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 41.660 53.140 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 45.960 52.730 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 45.530 52.730 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 45.100 52.730 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 44.670 52.730 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 44.240 52.730 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 43.810 52.730 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 43.380 52.730 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 42.950 52.730 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 42.520 52.730 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 42.090 52.730 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 41.660 52.730 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 45.960 52.320 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 45.530 52.320 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 45.100 52.320 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 44.670 52.320 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 44.240 52.320 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 43.810 52.320 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 43.380 52.320 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 42.950 52.320 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 42.520 52.320 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 42.090 52.320 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 41.660 52.320 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 45.960 51.910 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 45.530 51.910 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 45.100 51.910 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 44.670 51.910 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 44.240 51.910 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 43.810 51.910 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 43.380 51.910 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 42.950 51.910 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 42.520 51.910 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 42.090 51.910 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 41.660 51.910 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 45.960 51.500 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 45.530 51.500 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 45.100 51.500 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 44.670 51.500 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 44.240 51.500 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 43.810 51.500 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 43.380 51.500 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 42.950 51.500 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 42.520 51.500 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 42.090 51.500 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 41.660 51.500 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 45.960 51.090 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 45.530 51.090 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 45.100 51.090 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 44.670 51.090 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 44.240 51.090 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 43.810 51.090 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 43.380 51.090 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 42.950 51.090 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 42.520 51.090 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 42.090 51.090 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 41.660 51.090 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 45.960 50.680 46.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 45.530 50.680 45.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 45.100 50.680 45.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 44.670 50.680 44.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 44.240 50.680 44.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 43.810 50.680 44.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 43.380 50.680 43.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 42.950 50.680 43.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 42.520 50.680 42.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 42.090 50.680 42.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 41.660 50.680 41.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 45.900 24.365 46.220 ;
      LAYER met4 ;
        RECT 24.045 45.900 24.365 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 45.470 24.365 45.790 ;
      LAYER met4 ;
        RECT 24.045 45.470 24.365 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 45.040 24.365 45.360 ;
      LAYER met4 ;
        RECT 24.045 45.040 24.365 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 44.610 24.365 44.930 ;
      LAYER met4 ;
        RECT 24.045 44.610 24.365 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 44.180 24.365 44.500 ;
      LAYER met4 ;
        RECT 24.045 44.180 24.365 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 43.750 24.365 44.070 ;
      LAYER met4 ;
        RECT 24.045 43.750 24.365 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 43.320 24.365 43.640 ;
      LAYER met4 ;
        RECT 24.045 43.320 24.365 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 42.890 24.365 43.210 ;
      LAYER met4 ;
        RECT 24.045 42.890 24.365 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 42.460 24.365 42.780 ;
      LAYER met4 ;
        RECT 24.045 42.460 24.365 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 42.030 24.365 42.350 ;
      LAYER met4 ;
        RECT 24.045 42.030 24.365 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 41.600 24.365 41.920 ;
      LAYER met4 ;
        RECT 24.045 41.600 24.365 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 45.900 23.965 46.220 ;
      LAYER met4 ;
        RECT 23.645 45.900 23.965 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 45.470 23.965 45.790 ;
      LAYER met4 ;
        RECT 23.645 45.470 23.965 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 45.040 23.965 45.360 ;
      LAYER met4 ;
        RECT 23.645 45.040 23.965 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 44.610 23.965 44.930 ;
      LAYER met4 ;
        RECT 23.645 44.610 23.965 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 44.180 23.965 44.500 ;
      LAYER met4 ;
        RECT 23.645 44.180 23.965 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 43.750 23.965 44.070 ;
      LAYER met4 ;
        RECT 23.645 43.750 23.965 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 43.320 23.965 43.640 ;
      LAYER met4 ;
        RECT 23.645 43.320 23.965 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 42.890 23.965 43.210 ;
      LAYER met4 ;
        RECT 23.645 42.890 23.965 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 42.460 23.965 42.780 ;
      LAYER met4 ;
        RECT 23.645 42.460 23.965 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 42.030 23.965 42.350 ;
      LAYER met4 ;
        RECT 23.645 42.030 23.965 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 41.600 23.965 41.920 ;
      LAYER met4 ;
        RECT 23.645 41.600 23.965 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 45.900 23.565 46.220 ;
      LAYER met4 ;
        RECT 23.245 45.900 23.565 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 45.470 23.565 45.790 ;
      LAYER met4 ;
        RECT 23.245 45.470 23.565 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 45.040 23.565 45.360 ;
      LAYER met4 ;
        RECT 23.245 45.040 23.565 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 44.610 23.565 44.930 ;
      LAYER met4 ;
        RECT 23.245 44.610 23.565 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 44.180 23.565 44.500 ;
      LAYER met4 ;
        RECT 23.245 44.180 23.565 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 43.750 23.565 44.070 ;
      LAYER met4 ;
        RECT 23.245 43.750 23.565 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 43.320 23.565 43.640 ;
      LAYER met4 ;
        RECT 23.245 43.320 23.565 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 42.890 23.565 43.210 ;
      LAYER met4 ;
        RECT 23.245 42.890 23.565 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 42.460 23.565 42.780 ;
      LAYER met4 ;
        RECT 23.245 42.460 23.565 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 42.030 23.565 42.350 ;
      LAYER met4 ;
        RECT 23.245 42.030 23.565 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.245 41.600 23.565 41.920 ;
      LAYER met4 ;
        RECT 23.245 41.600 23.565 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 45.900 23.165 46.220 ;
      LAYER met4 ;
        RECT 22.845 45.900 23.165 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 45.470 23.165 45.790 ;
      LAYER met4 ;
        RECT 22.845 45.470 23.165 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 45.040 23.165 45.360 ;
      LAYER met4 ;
        RECT 22.845 45.040 23.165 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 44.610 23.165 44.930 ;
      LAYER met4 ;
        RECT 22.845 44.610 23.165 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 44.180 23.165 44.500 ;
      LAYER met4 ;
        RECT 22.845 44.180 23.165 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 43.750 23.165 44.070 ;
      LAYER met4 ;
        RECT 22.845 43.750 23.165 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 43.320 23.165 43.640 ;
      LAYER met4 ;
        RECT 22.845 43.320 23.165 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 42.890 23.165 43.210 ;
      LAYER met4 ;
        RECT 22.845 42.890 23.165 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 42.460 23.165 42.780 ;
      LAYER met4 ;
        RECT 22.845 42.460 23.165 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 42.030 23.165 42.350 ;
      LAYER met4 ;
        RECT 22.845 42.030 23.165 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.845 41.600 23.165 41.920 ;
      LAYER met4 ;
        RECT 22.845 41.600 23.165 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 45.900 22.765 46.220 ;
      LAYER met4 ;
        RECT 22.445 45.900 22.765 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 45.470 22.765 45.790 ;
      LAYER met4 ;
        RECT 22.445 45.470 22.765 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 45.040 22.765 45.360 ;
      LAYER met4 ;
        RECT 22.445 45.040 22.765 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 44.610 22.765 44.930 ;
      LAYER met4 ;
        RECT 22.445 44.610 22.765 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 44.180 22.765 44.500 ;
      LAYER met4 ;
        RECT 22.445 44.180 22.765 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 43.750 22.765 44.070 ;
      LAYER met4 ;
        RECT 22.445 43.750 22.765 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 43.320 22.765 43.640 ;
      LAYER met4 ;
        RECT 22.445 43.320 22.765 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 42.890 22.765 43.210 ;
      LAYER met4 ;
        RECT 22.445 42.890 22.765 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 42.460 22.765 42.780 ;
      LAYER met4 ;
        RECT 22.445 42.460 22.765 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 42.030 22.765 42.350 ;
      LAYER met4 ;
        RECT 22.445 42.030 22.765 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.445 41.600 22.765 41.920 ;
      LAYER met4 ;
        RECT 22.445 41.600 22.765 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 45.900 22.365 46.220 ;
      LAYER met4 ;
        RECT 22.045 45.900 22.365 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 45.470 22.365 45.790 ;
      LAYER met4 ;
        RECT 22.045 45.470 22.365 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 45.040 22.365 45.360 ;
      LAYER met4 ;
        RECT 22.045 45.040 22.365 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 44.610 22.365 44.930 ;
      LAYER met4 ;
        RECT 22.045 44.610 22.365 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 44.180 22.365 44.500 ;
      LAYER met4 ;
        RECT 22.045 44.180 22.365 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 43.750 22.365 44.070 ;
      LAYER met4 ;
        RECT 22.045 43.750 22.365 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 43.320 22.365 43.640 ;
      LAYER met4 ;
        RECT 22.045 43.320 22.365 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 42.890 22.365 43.210 ;
      LAYER met4 ;
        RECT 22.045 42.890 22.365 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 42.460 22.365 42.780 ;
      LAYER met4 ;
        RECT 22.045 42.460 22.365 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 42.030 22.365 42.350 ;
      LAYER met4 ;
        RECT 22.045 42.030 22.365 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.045 41.600 22.365 41.920 ;
      LAYER met4 ;
        RECT 22.045 41.600 22.365 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 45.900 21.965 46.220 ;
      LAYER met4 ;
        RECT 21.645 45.900 21.965 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 45.470 21.965 45.790 ;
      LAYER met4 ;
        RECT 21.645 45.470 21.965 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 45.040 21.965 45.360 ;
      LAYER met4 ;
        RECT 21.645 45.040 21.965 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 44.610 21.965 44.930 ;
      LAYER met4 ;
        RECT 21.645 44.610 21.965 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 44.180 21.965 44.500 ;
      LAYER met4 ;
        RECT 21.645 44.180 21.965 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 43.750 21.965 44.070 ;
      LAYER met4 ;
        RECT 21.645 43.750 21.965 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 43.320 21.965 43.640 ;
      LAYER met4 ;
        RECT 21.645 43.320 21.965 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 42.890 21.965 43.210 ;
      LAYER met4 ;
        RECT 21.645 42.890 21.965 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 42.460 21.965 42.780 ;
      LAYER met4 ;
        RECT 21.645 42.460 21.965 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 42.030 21.965 42.350 ;
      LAYER met4 ;
        RECT 21.645 42.030 21.965 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.645 41.600 21.965 41.920 ;
      LAYER met4 ;
        RECT 21.645 41.600 21.965 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 45.900 21.565 46.220 ;
      LAYER met4 ;
        RECT 21.245 45.900 21.565 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 45.470 21.565 45.790 ;
      LAYER met4 ;
        RECT 21.245 45.470 21.565 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 45.040 21.565 45.360 ;
      LAYER met4 ;
        RECT 21.245 45.040 21.565 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 44.610 21.565 44.930 ;
      LAYER met4 ;
        RECT 21.245 44.610 21.565 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 44.180 21.565 44.500 ;
      LAYER met4 ;
        RECT 21.245 44.180 21.565 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 43.750 21.565 44.070 ;
      LAYER met4 ;
        RECT 21.245 43.750 21.565 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 43.320 21.565 43.640 ;
      LAYER met4 ;
        RECT 21.245 43.320 21.565 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 42.890 21.565 43.210 ;
      LAYER met4 ;
        RECT 21.245 42.890 21.565 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 42.460 21.565 42.780 ;
      LAYER met4 ;
        RECT 21.245 42.460 21.565 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 42.030 21.565 42.350 ;
      LAYER met4 ;
        RECT 21.245 42.030 21.565 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.245 41.600 21.565 41.920 ;
      LAYER met4 ;
        RECT 21.245 41.600 21.565 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 45.900 21.165 46.220 ;
      LAYER met4 ;
        RECT 20.845 45.900 21.165 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 45.470 21.165 45.790 ;
      LAYER met4 ;
        RECT 20.845 45.470 21.165 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 45.040 21.165 45.360 ;
      LAYER met4 ;
        RECT 20.845 45.040 21.165 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 44.610 21.165 44.930 ;
      LAYER met4 ;
        RECT 20.845 44.610 21.165 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 44.180 21.165 44.500 ;
      LAYER met4 ;
        RECT 20.845 44.180 21.165 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 43.750 21.165 44.070 ;
      LAYER met4 ;
        RECT 20.845 43.750 21.165 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 43.320 21.165 43.640 ;
      LAYER met4 ;
        RECT 20.845 43.320 21.165 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 42.890 21.165 43.210 ;
      LAYER met4 ;
        RECT 20.845 42.890 21.165 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 42.460 21.165 42.780 ;
      LAYER met4 ;
        RECT 20.845 42.460 21.165 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 42.030 21.165 42.350 ;
      LAYER met4 ;
        RECT 20.845 42.030 21.165 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.845 41.600 21.165 41.920 ;
      LAYER met4 ;
        RECT 20.845 41.600 21.165 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 45.900 20.760 46.220 ;
      LAYER met4 ;
        RECT 20.440 45.900 20.760 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 45.470 20.760 45.790 ;
      LAYER met4 ;
        RECT 20.440 45.470 20.760 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 45.040 20.760 45.360 ;
      LAYER met4 ;
        RECT 20.440 45.040 20.760 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 44.610 20.760 44.930 ;
      LAYER met4 ;
        RECT 20.440 44.610 20.760 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 44.180 20.760 44.500 ;
      LAYER met4 ;
        RECT 20.440 44.180 20.760 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 43.750 20.760 44.070 ;
      LAYER met4 ;
        RECT 20.440 43.750 20.760 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 43.320 20.760 43.640 ;
      LAYER met4 ;
        RECT 20.440 43.320 20.760 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 42.890 20.760 43.210 ;
      LAYER met4 ;
        RECT 20.440 42.890 20.760 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 42.460 20.760 42.780 ;
      LAYER met4 ;
        RECT 20.440 42.460 20.760 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 42.030 20.760 42.350 ;
      LAYER met4 ;
        RECT 20.440 42.030 20.760 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.440 41.600 20.760 41.920 ;
      LAYER met4 ;
        RECT 20.440 41.600 20.760 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 45.900 20.355 46.220 ;
      LAYER met4 ;
        RECT 20.035 45.900 20.355 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 45.470 20.355 45.790 ;
      LAYER met4 ;
        RECT 20.035 45.470 20.355 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 45.040 20.355 45.360 ;
      LAYER met4 ;
        RECT 20.035 45.040 20.355 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 44.610 20.355 44.930 ;
      LAYER met4 ;
        RECT 20.035 44.610 20.355 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 44.180 20.355 44.500 ;
      LAYER met4 ;
        RECT 20.035 44.180 20.355 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 43.750 20.355 44.070 ;
      LAYER met4 ;
        RECT 20.035 43.750 20.355 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 43.320 20.355 43.640 ;
      LAYER met4 ;
        RECT 20.035 43.320 20.355 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 42.890 20.355 43.210 ;
      LAYER met4 ;
        RECT 20.035 42.890 20.355 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 42.460 20.355 42.780 ;
      LAYER met4 ;
        RECT 20.035 42.460 20.355 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 42.030 20.355 42.350 ;
      LAYER met4 ;
        RECT 20.035 42.030 20.355 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.035 41.600 20.355 41.920 ;
      LAYER met4 ;
        RECT 20.035 41.600 20.355 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 45.900 19.950 46.220 ;
      LAYER met4 ;
        RECT 19.630 45.900 19.950 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 45.470 19.950 45.790 ;
      LAYER met4 ;
        RECT 19.630 45.470 19.950 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 45.040 19.950 45.360 ;
      LAYER met4 ;
        RECT 19.630 45.040 19.950 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 44.610 19.950 44.930 ;
      LAYER met4 ;
        RECT 19.630 44.610 19.950 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 44.180 19.950 44.500 ;
      LAYER met4 ;
        RECT 19.630 44.180 19.950 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 43.750 19.950 44.070 ;
      LAYER met4 ;
        RECT 19.630 43.750 19.950 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 43.320 19.950 43.640 ;
      LAYER met4 ;
        RECT 19.630 43.320 19.950 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 42.890 19.950 43.210 ;
      LAYER met4 ;
        RECT 19.630 42.890 19.950 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 42.460 19.950 42.780 ;
      LAYER met4 ;
        RECT 19.630 42.460 19.950 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 42.030 19.950 42.350 ;
      LAYER met4 ;
        RECT 19.630 42.030 19.950 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.630 41.600 19.950 41.920 ;
      LAYER met4 ;
        RECT 19.630 41.600 19.950 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 45.900 19.545 46.220 ;
      LAYER met4 ;
        RECT 19.225 45.900 19.545 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 45.470 19.545 45.790 ;
      LAYER met4 ;
        RECT 19.225 45.470 19.545 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 45.040 19.545 45.360 ;
      LAYER met4 ;
        RECT 19.225 45.040 19.545 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 44.610 19.545 44.930 ;
      LAYER met4 ;
        RECT 19.225 44.610 19.545 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 44.180 19.545 44.500 ;
      LAYER met4 ;
        RECT 19.225 44.180 19.545 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 43.750 19.545 44.070 ;
      LAYER met4 ;
        RECT 19.225 43.750 19.545 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 43.320 19.545 43.640 ;
      LAYER met4 ;
        RECT 19.225 43.320 19.545 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 42.890 19.545 43.210 ;
      LAYER met4 ;
        RECT 19.225 42.890 19.545 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 42.460 19.545 42.780 ;
      LAYER met4 ;
        RECT 19.225 42.460 19.545 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 42.030 19.545 42.350 ;
      LAYER met4 ;
        RECT 19.225 42.030 19.545 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.225 41.600 19.545 41.920 ;
      LAYER met4 ;
        RECT 19.225 41.600 19.545 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 45.900 19.140 46.220 ;
      LAYER met4 ;
        RECT 18.820 45.900 19.140 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 45.470 19.140 45.790 ;
      LAYER met4 ;
        RECT 18.820 45.470 19.140 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 45.040 19.140 45.360 ;
      LAYER met4 ;
        RECT 18.820 45.040 19.140 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 44.610 19.140 44.930 ;
      LAYER met4 ;
        RECT 18.820 44.610 19.140 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 44.180 19.140 44.500 ;
      LAYER met4 ;
        RECT 18.820 44.180 19.140 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 43.750 19.140 44.070 ;
      LAYER met4 ;
        RECT 18.820 43.750 19.140 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 43.320 19.140 43.640 ;
      LAYER met4 ;
        RECT 18.820 43.320 19.140 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 42.890 19.140 43.210 ;
      LAYER met4 ;
        RECT 18.820 42.890 19.140 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 42.460 19.140 42.780 ;
      LAYER met4 ;
        RECT 18.820 42.460 19.140 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 42.030 19.140 42.350 ;
      LAYER met4 ;
        RECT 18.820 42.030 19.140 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.820 41.600 19.140 41.920 ;
      LAYER met4 ;
        RECT 18.820 41.600 19.140 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 45.900 18.735 46.220 ;
      LAYER met4 ;
        RECT 18.415 45.900 18.735 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 45.470 18.735 45.790 ;
      LAYER met4 ;
        RECT 18.415 45.470 18.735 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 45.040 18.735 45.360 ;
      LAYER met4 ;
        RECT 18.415 45.040 18.735 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 44.610 18.735 44.930 ;
      LAYER met4 ;
        RECT 18.415 44.610 18.735 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 44.180 18.735 44.500 ;
      LAYER met4 ;
        RECT 18.415 44.180 18.735 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 43.750 18.735 44.070 ;
      LAYER met4 ;
        RECT 18.415 43.750 18.735 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 43.320 18.735 43.640 ;
      LAYER met4 ;
        RECT 18.415 43.320 18.735 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 42.890 18.735 43.210 ;
      LAYER met4 ;
        RECT 18.415 42.890 18.735 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 42.460 18.735 42.780 ;
      LAYER met4 ;
        RECT 18.415 42.460 18.735 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 42.030 18.735 42.350 ;
      LAYER met4 ;
        RECT 18.415 42.030 18.735 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.415 41.600 18.735 41.920 ;
      LAYER met4 ;
        RECT 18.415 41.600 18.735 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 45.900 18.330 46.220 ;
      LAYER met4 ;
        RECT 18.010 45.900 18.330 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 45.470 18.330 45.790 ;
      LAYER met4 ;
        RECT 18.010 45.470 18.330 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 45.040 18.330 45.360 ;
      LAYER met4 ;
        RECT 18.010 45.040 18.330 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 44.610 18.330 44.930 ;
      LAYER met4 ;
        RECT 18.010 44.610 18.330 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 44.180 18.330 44.500 ;
      LAYER met4 ;
        RECT 18.010 44.180 18.330 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 43.750 18.330 44.070 ;
      LAYER met4 ;
        RECT 18.010 43.750 18.330 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 43.320 18.330 43.640 ;
      LAYER met4 ;
        RECT 18.010 43.320 18.330 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 42.890 18.330 43.210 ;
      LAYER met4 ;
        RECT 18.010 42.890 18.330 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 42.460 18.330 42.780 ;
      LAYER met4 ;
        RECT 18.010 42.460 18.330 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 42.030 18.330 42.350 ;
      LAYER met4 ;
        RECT 18.010 42.030 18.330 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.010 41.600 18.330 41.920 ;
      LAYER met4 ;
        RECT 18.010 41.600 18.330 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 45.900 17.925 46.220 ;
      LAYER met4 ;
        RECT 17.605 45.900 17.925 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 45.470 17.925 45.790 ;
      LAYER met4 ;
        RECT 17.605 45.470 17.925 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 45.040 17.925 45.360 ;
      LAYER met4 ;
        RECT 17.605 45.040 17.925 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 44.610 17.925 44.930 ;
      LAYER met4 ;
        RECT 17.605 44.610 17.925 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 44.180 17.925 44.500 ;
      LAYER met4 ;
        RECT 17.605 44.180 17.925 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 43.750 17.925 44.070 ;
      LAYER met4 ;
        RECT 17.605 43.750 17.925 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 43.320 17.925 43.640 ;
      LAYER met4 ;
        RECT 17.605 43.320 17.925 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 42.890 17.925 43.210 ;
      LAYER met4 ;
        RECT 17.605 42.890 17.925 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 42.460 17.925 42.780 ;
      LAYER met4 ;
        RECT 17.605 42.460 17.925 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 42.030 17.925 42.350 ;
      LAYER met4 ;
        RECT 17.605 42.030 17.925 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.605 41.600 17.925 41.920 ;
      LAYER met4 ;
        RECT 17.605 41.600 17.925 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 45.900 17.520 46.220 ;
      LAYER met4 ;
        RECT 17.200 45.900 17.520 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 45.470 17.520 45.790 ;
      LAYER met4 ;
        RECT 17.200 45.470 17.520 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 45.040 17.520 45.360 ;
      LAYER met4 ;
        RECT 17.200 45.040 17.520 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 44.610 17.520 44.930 ;
      LAYER met4 ;
        RECT 17.200 44.610 17.520 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 44.180 17.520 44.500 ;
      LAYER met4 ;
        RECT 17.200 44.180 17.520 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 43.750 17.520 44.070 ;
      LAYER met4 ;
        RECT 17.200 43.750 17.520 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 43.320 17.520 43.640 ;
      LAYER met4 ;
        RECT 17.200 43.320 17.520 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 42.890 17.520 43.210 ;
      LAYER met4 ;
        RECT 17.200 42.890 17.520 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 42.460 17.520 42.780 ;
      LAYER met4 ;
        RECT 17.200 42.460 17.520 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 42.030 17.520 42.350 ;
      LAYER met4 ;
        RECT 17.200 42.030 17.520 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.200 41.600 17.520 41.920 ;
      LAYER met4 ;
        RECT 17.200 41.600 17.520 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 45.900 17.115 46.220 ;
      LAYER met4 ;
        RECT 16.795 45.900 17.115 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 45.470 17.115 45.790 ;
      LAYER met4 ;
        RECT 16.795 45.470 17.115 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 45.040 17.115 45.360 ;
      LAYER met4 ;
        RECT 16.795 45.040 17.115 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 44.610 17.115 44.930 ;
      LAYER met4 ;
        RECT 16.795 44.610 17.115 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 44.180 17.115 44.500 ;
      LAYER met4 ;
        RECT 16.795 44.180 17.115 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 43.750 17.115 44.070 ;
      LAYER met4 ;
        RECT 16.795 43.750 17.115 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 43.320 17.115 43.640 ;
      LAYER met4 ;
        RECT 16.795 43.320 17.115 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 42.890 17.115 43.210 ;
      LAYER met4 ;
        RECT 16.795 42.890 17.115 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 42.460 17.115 42.780 ;
      LAYER met4 ;
        RECT 16.795 42.460 17.115 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 42.030 17.115 42.350 ;
      LAYER met4 ;
        RECT 16.795 42.030 17.115 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.795 41.600 17.115 41.920 ;
      LAYER met4 ;
        RECT 16.795 41.600 17.115 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 45.900 16.710 46.220 ;
      LAYER met4 ;
        RECT 16.390 45.900 16.710 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 45.470 16.710 45.790 ;
      LAYER met4 ;
        RECT 16.390 45.470 16.710 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 45.040 16.710 45.360 ;
      LAYER met4 ;
        RECT 16.390 45.040 16.710 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 44.610 16.710 44.930 ;
      LAYER met4 ;
        RECT 16.390 44.610 16.710 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 44.180 16.710 44.500 ;
      LAYER met4 ;
        RECT 16.390 44.180 16.710 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 43.750 16.710 44.070 ;
      LAYER met4 ;
        RECT 16.390 43.750 16.710 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 43.320 16.710 43.640 ;
      LAYER met4 ;
        RECT 16.390 43.320 16.710 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 42.890 16.710 43.210 ;
      LAYER met4 ;
        RECT 16.390 42.890 16.710 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 42.460 16.710 42.780 ;
      LAYER met4 ;
        RECT 16.390 42.460 16.710 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 42.030 16.710 42.350 ;
      LAYER met4 ;
        RECT 16.390 42.030 16.710 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.390 41.600 16.710 41.920 ;
      LAYER met4 ;
        RECT 16.390 41.600 16.710 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 45.900 16.305 46.220 ;
      LAYER met4 ;
        RECT 15.985 45.900 16.305 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 45.470 16.305 45.790 ;
      LAYER met4 ;
        RECT 15.985 45.470 16.305 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 45.040 16.305 45.360 ;
      LAYER met4 ;
        RECT 15.985 45.040 16.305 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 44.610 16.305 44.930 ;
      LAYER met4 ;
        RECT 15.985 44.610 16.305 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 44.180 16.305 44.500 ;
      LAYER met4 ;
        RECT 15.985 44.180 16.305 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 43.750 16.305 44.070 ;
      LAYER met4 ;
        RECT 15.985 43.750 16.305 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 43.320 16.305 43.640 ;
      LAYER met4 ;
        RECT 15.985 43.320 16.305 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 42.890 16.305 43.210 ;
      LAYER met4 ;
        RECT 15.985 42.890 16.305 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 42.460 16.305 42.780 ;
      LAYER met4 ;
        RECT 15.985 42.460 16.305 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 42.030 16.305 42.350 ;
      LAYER met4 ;
        RECT 15.985 42.030 16.305 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.985 41.600 16.305 41.920 ;
      LAYER met4 ;
        RECT 15.985 41.600 16.305 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 45.900 15.900 46.220 ;
      LAYER met4 ;
        RECT 15.580 45.900 15.900 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 45.470 15.900 45.790 ;
      LAYER met4 ;
        RECT 15.580 45.470 15.900 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 45.040 15.900 45.360 ;
      LAYER met4 ;
        RECT 15.580 45.040 15.900 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 44.610 15.900 44.930 ;
      LAYER met4 ;
        RECT 15.580 44.610 15.900 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 44.180 15.900 44.500 ;
      LAYER met4 ;
        RECT 15.580 44.180 15.900 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 43.750 15.900 44.070 ;
      LAYER met4 ;
        RECT 15.580 43.750 15.900 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 43.320 15.900 43.640 ;
      LAYER met4 ;
        RECT 15.580 43.320 15.900 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 42.890 15.900 43.210 ;
      LAYER met4 ;
        RECT 15.580 42.890 15.900 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 42.460 15.900 42.780 ;
      LAYER met4 ;
        RECT 15.580 42.460 15.900 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 42.030 15.900 42.350 ;
      LAYER met4 ;
        RECT 15.580 42.030 15.900 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.580 41.600 15.900 41.920 ;
      LAYER met4 ;
        RECT 15.580 41.600 15.900 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 45.900 15.495 46.220 ;
      LAYER met4 ;
        RECT 15.175 45.900 15.495 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 45.470 15.495 45.790 ;
      LAYER met4 ;
        RECT 15.175 45.470 15.495 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 45.040 15.495 45.360 ;
      LAYER met4 ;
        RECT 15.175 45.040 15.495 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 44.610 15.495 44.930 ;
      LAYER met4 ;
        RECT 15.175 44.610 15.495 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 44.180 15.495 44.500 ;
      LAYER met4 ;
        RECT 15.175 44.180 15.495 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 43.750 15.495 44.070 ;
      LAYER met4 ;
        RECT 15.175 43.750 15.495 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 43.320 15.495 43.640 ;
      LAYER met4 ;
        RECT 15.175 43.320 15.495 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 42.890 15.495 43.210 ;
      LAYER met4 ;
        RECT 15.175 42.890 15.495 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 42.460 15.495 42.780 ;
      LAYER met4 ;
        RECT 15.175 42.460 15.495 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 42.030 15.495 42.350 ;
      LAYER met4 ;
        RECT 15.175 42.030 15.495 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.175 41.600 15.495 41.920 ;
      LAYER met4 ;
        RECT 15.175 41.600 15.495 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 45.900 15.090 46.220 ;
      LAYER met4 ;
        RECT 14.770 45.900 15.090 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 45.470 15.090 45.790 ;
      LAYER met4 ;
        RECT 14.770 45.470 15.090 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 45.040 15.090 45.360 ;
      LAYER met4 ;
        RECT 14.770 45.040 15.090 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 44.610 15.090 44.930 ;
      LAYER met4 ;
        RECT 14.770 44.610 15.090 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 44.180 15.090 44.500 ;
      LAYER met4 ;
        RECT 14.770 44.180 15.090 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 43.750 15.090 44.070 ;
      LAYER met4 ;
        RECT 14.770 43.750 15.090 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 43.320 15.090 43.640 ;
      LAYER met4 ;
        RECT 14.770 43.320 15.090 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 42.890 15.090 43.210 ;
      LAYER met4 ;
        RECT 14.770 42.890 15.090 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 42.460 15.090 42.780 ;
      LAYER met4 ;
        RECT 14.770 42.460 15.090 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 42.030 15.090 42.350 ;
      LAYER met4 ;
        RECT 14.770 42.030 15.090 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.770 41.600 15.090 41.920 ;
      LAYER met4 ;
        RECT 14.770 41.600 15.090 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 45.900 14.685 46.220 ;
      LAYER met4 ;
        RECT 14.365 45.900 14.685 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 45.470 14.685 45.790 ;
      LAYER met4 ;
        RECT 14.365 45.470 14.685 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 45.040 14.685 45.360 ;
      LAYER met4 ;
        RECT 14.365 45.040 14.685 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 44.610 14.685 44.930 ;
      LAYER met4 ;
        RECT 14.365 44.610 14.685 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 44.180 14.685 44.500 ;
      LAYER met4 ;
        RECT 14.365 44.180 14.685 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 43.750 14.685 44.070 ;
      LAYER met4 ;
        RECT 14.365 43.750 14.685 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 43.320 14.685 43.640 ;
      LAYER met4 ;
        RECT 14.365 43.320 14.685 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 42.890 14.685 43.210 ;
      LAYER met4 ;
        RECT 14.365 42.890 14.685 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 42.460 14.685 42.780 ;
      LAYER met4 ;
        RECT 14.365 42.460 14.685 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 42.030 14.685 42.350 ;
      LAYER met4 ;
        RECT 14.365 42.030 14.685 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.365 41.600 14.685 41.920 ;
      LAYER met4 ;
        RECT 14.365 41.600 14.685 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 45.900 14.280 46.220 ;
      LAYER met4 ;
        RECT 13.960 45.900 14.280 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 45.470 14.280 45.790 ;
      LAYER met4 ;
        RECT 13.960 45.470 14.280 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 45.040 14.280 45.360 ;
      LAYER met4 ;
        RECT 13.960 45.040 14.280 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 44.610 14.280 44.930 ;
      LAYER met4 ;
        RECT 13.960 44.610 14.280 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 44.180 14.280 44.500 ;
      LAYER met4 ;
        RECT 13.960 44.180 14.280 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 43.750 14.280 44.070 ;
      LAYER met4 ;
        RECT 13.960 43.750 14.280 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 43.320 14.280 43.640 ;
      LAYER met4 ;
        RECT 13.960 43.320 14.280 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 42.890 14.280 43.210 ;
      LAYER met4 ;
        RECT 13.960 42.890 14.280 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 42.460 14.280 42.780 ;
      LAYER met4 ;
        RECT 13.960 42.460 14.280 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 42.030 14.280 42.350 ;
      LAYER met4 ;
        RECT 13.960 42.030 14.280 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.960 41.600 14.280 41.920 ;
      LAYER met4 ;
        RECT 13.960 41.600 14.280 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 45.900 13.875 46.220 ;
      LAYER met4 ;
        RECT 13.555 45.900 13.875 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 45.470 13.875 45.790 ;
      LAYER met4 ;
        RECT 13.555 45.470 13.875 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 45.040 13.875 45.360 ;
      LAYER met4 ;
        RECT 13.555 45.040 13.875 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 44.610 13.875 44.930 ;
      LAYER met4 ;
        RECT 13.555 44.610 13.875 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 44.180 13.875 44.500 ;
      LAYER met4 ;
        RECT 13.555 44.180 13.875 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 43.750 13.875 44.070 ;
      LAYER met4 ;
        RECT 13.555 43.750 13.875 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 43.320 13.875 43.640 ;
      LAYER met4 ;
        RECT 13.555 43.320 13.875 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 42.890 13.875 43.210 ;
      LAYER met4 ;
        RECT 13.555 42.890 13.875 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 42.460 13.875 42.780 ;
      LAYER met4 ;
        RECT 13.555 42.460 13.875 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 42.030 13.875 42.350 ;
      LAYER met4 ;
        RECT 13.555 42.030 13.875 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.555 41.600 13.875 41.920 ;
      LAYER met4 ;
        RECT 13.555 41.600 13.875 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 45.900 13.470 46.220 ;
      LAYER met4 ;
        RECT 13.150 45.900 13.470 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 45.470 13.470 45.790 ;
      LAYER met4 ;
        RECT 13.150 45.470 13.470 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 45.040 13.470 45.360 ;
      LAYER met4 ;
        RECT 13.150 45.040 13.470 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 44.610 13.470 44.930 ;
      LAYER met4 ;
        RECT 13.150 44.610 13.470 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 44.180 13.470 44.500 ;
      LAYER met4 ;
        RECT 13.150 44.180 13.470 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 43.750 13.470 44.070 ;
      LAYER met4 ;
        RECT 13.150 43.750 13.470 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 43.320 13.470 43.640 ;
      LAYER met4 ;
        RECT 13.150 43.320 13.470 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 42.890 13.470 43.210 ;
      LAYER met4 ;
        RECT 13.150 42.890 13.470 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 42.460 13.470 42.780 ;
      LAYER met4 ;
        RECT 13.150 42.460 13.470 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 42.030 13.470 42.350 ;
      LAYER met4 ;
        RECT 13.150 42.030 13.470 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.150 41.600 13.470 41.920 ;
      LAYER met4 ;
        RECT 13.150 41.600 13.470 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 45.900 13.065 46.220 ;
      LAYER met4 ;
        RECT 12.745 45.900 13.065 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 45.470 13.065 45.790 ;
      LAYER met4 ;
        RECT 12.745 45.470 13.065 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 45.040 13.065 45.360 ;
      LAYER met4 ;
        RECT 12.745 45.040 13.065 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 44.610 13.065 44.930 ;
      LAYER met4 ;
        RECT 12.745 44.610 13.065 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 44.180 13.065 44.500 ;
      LAYER met4 ;
        RECT 12.745 44.180 13.065 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 43.750 13.065 44.070 ;
      LAYER met4 ;
        RECT 12.745 43.750 13.065 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 43.320 13.065 43.640 ;
      LAYER met4 ;
        RECT 12.745 43.320 13.065 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 42.890 13.065 43.210 ;
      LAYER met4 ;
        RECT 12.745 42.890 13.065 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 42.460 13.065 42.780 ;
      LAYER met4 ;
        RECT 12.745 42.460 13.065 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 42.030 13.065 42.350 ;
      LAYER met4 ;
        RECT 12.745 42.030 13.065 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.745 41.600 13.065 41.920 ;
      LAYER met4 ;
        RECT 12.745 41.600 13.065 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 45.900 12.660 46.220 ;
      LAYER met4 ;
        RECT 12.340 45.900 12.660 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 45.470 12.660 45.790 ;
      LAYER met4 ;
        RECT 12.340 45.470 12.660 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 45.040 12.660 45.360 ;
      LAYER met4 ;
        RECT 12.340 45.040 12.660 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 44.610 12.660 44.930 ;
      LAYER met4 ;
        RECT 12.340 44.610 12.660 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 44.180 12.660 44.500 ;
      LAYER met4 ;
        RECT 12.340 44.180 12.660 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 43.750 12.660 44.070 ;
      LAYER met4 ;
        RECT 12.340 43.750 12.660 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 43.320 12.660 43.640 ;
      LAYER met4 ;
        RECT 12.340 43.320 12.660 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 42.890 12.660 43.210 ;
      LAYER met4 ;
        RECT 12.340 42.890 12.660 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 42.460 12.660 42.780 ;
      LAYER met4 ;
        RECT 12.340 42.460 12.660 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 42.030 12.660 42.350 ;
      LAYER met4 ;
        RECT 12.340 42.030 12.660 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.340 41.600 12.660 41.920 ;
      LAYER met4 ;
        RECT 12.340 41.600 12.660 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 45.900 12.255 46.220 ;
      LAYER met4 ;
        RECT 11.935 45.900 12.255 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 45.470 12.255 45.790 ;
      LAYER met4 ;
        RECT 11.935 45.470 12.255 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 45.040 12.255 45.360 ;
      LAYER met4 ;
        RECT 11.935 45.040 12.255 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 44.610 12.255 44.930 ;
      LAYER met4 ;
        RECT 11.935 44.610 12.255 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 44.180 12.255 44.500 ;
      LAYER met4 ;
        RECT 11.935 44.180 12.255 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 43.750 12.255 44.070 ;
      LAYER met4 ;
        RECT 11.935 43.750 12.255 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 43.320 12.255 43.640 ;
      LAYER met4 ;
        RECT 11.935 43.320 12.255 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 42.890 12.255 43.210 ;
      LAYER met4 ;
        RECT 11.935 42.890 12.255 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 42.460 12.255 42.780 ;
      LAYER met4 ;
        RECT 11.935 42.460 12.255 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 42.030 12.255 42.350 ;
      LAYER met4 ;
        RECT 11.935 42.030 12.255 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.935 41.600 12.255 41.920 ;
      LAYER met4 ;
        RECT 11.935 41.600 12.255 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 45.900 11.850 46.220 ;
      LAYER met4 ;
        RECT 11.530 45.900 11.850 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 45.470 11.850 45.790 ;
      LAYER met4 ;
        RECT 11.530 45.470 11.850 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 45.040 11.850 45.360 ;
      LAYER met4 ;
        RECT 11.530 45.040 11.850 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 44.610 11.850 44.930 ;
      LAYER met4 ;
        RECT 11.530 44.610 11.850 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 44.180 11.850 44.500 ;
      LAYER met4 ;
        RECT 11.530 44.180 11.850 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 43.750 11.850 44.070 ;
      LAYER met4 ;
        RECT 11.530 43.750 11.850 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 43.320 11.850 43.640 ;
      LAYER met4 ;
        RECT 11.530 43.320 11.850 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 42.890 11.850 43.210 ;
      LAYER met4 ;
        RECT 11.530 42.890 11.850 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 42.460 11.850 42.780 ;
      LAYER met4 ;
        RECT 11.530 42.460 11.850 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 42.030 11.850 42.350 ;
      LAYER met4 ;
        RECT 11.530 42.030 11.850 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.530 41.600 11.850 41.920 ;
      LAYER met4 ;
        RECT 11.530 41.600 11.850 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 45.900 11.445 46.220 ;
      LAYER met4 ;
        RECT 11.125 45.900 11.445 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 45.470 11.445 45.790 ;
      LAYER met4 ;
        RECT 11.125 45.470 11.445 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 45.040 11.445 45.360 ;
      LAYER met4 ;
        RECT 11.125 45.040 11.445 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 44.610 11.445 44.930 ;
      LAYER met4 ;
        RECT 11.125 44.610 11.445 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 44.180 11.445 44.500 ;
      LAYER met4 ;
        RECT 11.125 44.180 11.445 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 43.750 11.445 44.070 ;
      LAYER met4 ;
        RECT 11.125 43.750 11.445 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 43.320 11.445 43.640 ;
      LAYER met4 ;
        RECT 11.125 43.320 11.445 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 42.890 11.445 43.210 ;
      LAYER met4 ;
        RECT 11.125 42.890 11.445 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 42.460 11.445 42.780 ;
      LAYER met4 ;
        RECT 11.125 42.460 11.445 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 42.030 11.445 42.350 ;
      LAYER met4 ;
        RECT 11.125 42.030 11.445 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.125 41.600 11.445 41.920 ;
      LAYER met4 ;
        RECT 11.125 41.600 11.445 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 45.900 11.040 46.220 ;
      LAYER met4 ;
        RECT 10.720 45.900 11.040 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 45.470 11.040 45.790 ;
      LAYER met4 ;
        RECT 10.720 45.470 11.040 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 45.040 11.040 45.360 ;
      LAYER met4 ;
        RECT 10.720 45.040 11.040 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 44.610 11.040 44.930 ;
      LAYER met4 ;
        RECT 10.720 44.610 11.040 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 44.180 11.040 44.500 ;
      LAYER met4 ;
        RECT 10.720 44.180 11.040 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 43.750 11.040 44.070 ;
      LAYER met4 ;
        RECT 10.720 43.750 11.040 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 43.320 11.040 43.640 ;
      LAYER met4 ;
        RECT 10.720 43.320 11.040 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 42.890 11.040 43.210 ;
      LAYER met4 ;
        RECT 10.720 42.890 11.040 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 42.460 11.040 42.780 ;
      LAYER met4 ;
        RECT 10.720 42.460 11.040 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 42.030 11.040 42.350 ;
      LAYER met4 ;
        RECT 10.720 42.030 11.040 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.720 41.600 11.040 41.920 ;
      LAYER met4 ;
        RECT 10.720 41.600 11.040 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 45.900 10.635 46.220 ;
      LAYER met4 ;
        RECT 10.315 45.900 10.635 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 45.470 10.635 45.790 ;
      LAYER met4 ;
        RECT 10.315 45.470 10.635 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 45.040 10.635 45.360 ;
      LAYER met4 ;
        RECT 10.315 45.040 10.635 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 44.610 10.635 44.930 ;
      LAYER met4 ;
        RECT 10.315 44.610 10.635 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 44.180 10.635 44.500 ;
      LAYER met4 ;
        RECT 10.315 44.180 10.635 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 43.750 10.635 44.070 ;
      LAYER met4 ;
        RECT 10.315 43.750 10.635 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 43.320 10.635 43.640 ;
      LAYER met4 ;
        RECT 10.315 43.320 10.635 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 42.890 10.635 43.210 ;
      LAYER met4 ;
        RECT 10.315 42.890 10.635 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 42.460 10.635 42.780 ;
      LAYER met4 ;
        RECT 10.315 42.460 10.635 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 42.030 10.635 42.350 ;
      LAYER met4 ;
        RECT 10.315 42.030 10.635 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.315 41.600 10.635 41.920 ;
      LAYER met4 ;
        RECT 10.315 41.600 10.635 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 45.900 10.230 46.220 ;
      LAYER met4 ;
        RECT 9.910 45.900 10.230 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 45.470 10.230 45.790 ;
      LAYER met4 ;
        RECT 9.910 45.470 10.230 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 45.040 10.230 45.360 ;
      LAYER met4 ;
        RECT 9.910 45.040 10.230 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 44.610 10.230 44.930 ;
      LAYER met4 ;
        RECT 9.910 44.610 10.230 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 44.180 10.230 44.500 ;
      LAYER met4 ;
        RECT 9.910 44.180 10.230 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 43.750 10.230 44.070 ;
      LAYER met4 ;
        RECT 9.910 43.750 10.230 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 43.320 10.230 43.640 ;
      LAYER met4 ;
        RECT 9.910 43.320 10.230 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 42.890 10.230 43.210 ;
      LAYER met4 ;
        RECT 9.910 42.890 10.230 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 42.460 10.230 42.780 ;
      LAYER met4 ;
        RECT 9.910 42.460 10.230 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 42.030 10.230 42.350 ;
      LAYER met4 ;
        RECT 9.910 42.030 10.230 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.910 41.600 10.230 41.920 ;
      LAYER met4 ;
        RECT 9.910 41.600 10.230 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 45.900 9.825 46.220 ;
      LAYER met4 ;
        RECT 9.505 45.900 9.825 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 45.470 9.825 45.790 ;
      LAYER met4 ;
        RECT 9.505 45.470 9.825 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 45.040 9.825 45.360 ;
      LAYER met4 ;
        RECT 9.505 45.040 9.825 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 44.610 9.825 44.930 ;
      LAYER met4 ;
        RECT 9.505 44.610 9.825 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 44.180 9.825 44.500 ;
      LAYER met4 ;
        RECT 9.505 44.180 9.825 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 43.750 9.825 44.070 ;
      LAYER met4 ;
        RECT 9.505 43.750 9.825 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 43.320 9.825 43.640 ;
      LAYER met4 ;
        RECT 9.505 43.320 9.825 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 42.890 9.825 43.210 ;
      LAYER met4 ;
        RECT 9.505 42.890 9.825 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 42.460 9.825 42.780 ;
      LAYER met4 ;
        RECT 9.505 42.460 9.825 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 42.030 9.825 42.350 ;
      LAYER met4 ;
        RECT 9.505 42.030 9.825 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.505 41.600 9.825 41.920 ;
      LAYER met4 ;
        RECT 9.505 41.600 9.825 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 45.900 9.420 46.220 ;
      LAYER met4 ;
        RECT 9.100 45.900 9.420 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 45.470 9.420 45.790 ;
      LAYER met4 ;
        RECT 9.100 45.470 9.420 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 45.040 9.420 45.360 ;
      LAYER met4 ;
        RECT 9.100 45.040 9.420 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 44.610 9.420 44.930 ;
      LAYER met4 ;
        RECT 9.100 44.610 9.420 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 44.180 9.420 44.500 ;
      LAYER met4 ;
        RECT 9.100 44.180 9.420 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 43.750 9.420 44.070 ;
      LAYER met4 ;
        RECT 9.100 43.750 9.420 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 43.320 9.420 43.640 ;
      LAYER met4 ;
        RECT 9.100 43.320 9.420 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 42.890 9.420 43.210 ;
      LAYER met4 ;
        RECT 9.100 42.890 9.420 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 42.460 9.420 42.780 ;
      LAYER met4 ;
        RECT 9.100 42.460 9.420 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 42.030 9.420 42.350 ;
      LAYER met4 ;
        RECT 9.100 42.030 9.420 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.100 41.600 9.420 41.920 ;
      LAYER met4 ;
        RECT 9.100 41.600 9.420 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 45.900 9.015 46.220 ;
      LAYER met4 ;
        RECT 8.695 45.900 9.015 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 45.470 9.015 45.790 ;
      LAYER met4 ;
        RECT 8.695 45.470 9.015 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 45.040 9.015 45.360 ;
      LAYER met4 ;
        RECT 8.695 45.040 9.015 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 44.610 9.015 44.930 ;
      LAYER met4 ;
        RECT 8.695 44.610 9.015 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 44.180 9.015 44.500 ;
      LAYER met4 ;
        RECT 8.695 44.180 9.015 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 43.750 9.015 44.070 ;
      LAYER met4 ;
        RECT 8.695 43.750 9.015 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 43.320 9.015 43.640 ;
      LAYER met4 ;
        RECT 8.695 43.320 9.015 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 42.890 9.015 43.210 ;
      LAYER met4 ;
        RECT 8.695 42.890 9.015 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 42.460 9.015 42.780 ;
      LAYER met4 ;
        RECT 8.695 42.460 9.015 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 42.030 9.015 42.350 ;
      LAYER met4 ;
        RECT 8.695 42.030 9.015 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.695 41.600 9.015 41.920 ;
      LAYER met4 ;
        RECT 8.695 41.600 9.015 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 45.900 8.610 46.220 ;
      LAYER met4 ;
        RECT 8.290 45.900 8.610 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 45.470 8.610 45.790 ;
      LAYER met4 ;
        RECT 8.290 45.470 8.610 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 45.040 8.610 45.360 ;
      LAYER met4 ;
        RECT 8.290 45.040 8.610 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 44.610 8.610 44.930 ;
      LAYER met4 ;
        RECT 8.290 44.610 8.610 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 44.180 8.610 44.500 ;
      LAYER met4 ;
        RECT 8.290 44.180 8.610 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 43.750 8.610 44.070 ;
      LAYER met4 ;
        RECT 8.290 43.750 8.610 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 43.320 8.610 43.640 ;
      LAYER met4 ;
        RECT 8.290 43.320 8.610 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 42.890 8.610 43.210 ;
      LAYER met4 ;
        RECT 8.290 42.890 8.610 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 42.460 8.610 42.780 ;
      LAYER met4 ;
        RECT 8.290 42.460 8.610 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 42.030 8.610 42.350 ;
      LAYER met4 ;
        RECT 8.290 42.030 8.610 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.290 41.600 8.610 41.920 ;
      LAYER met4 ;
        RECT 8.290 41.600 8.610 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 45.900 8.205 46.220 ;
      LAYER met4 ;
        RECT 7.885 45.900 8.205 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 45.470 8.205 45.790 ;
      LAYER met4 ;
        RECT 7.885 45.470 8.205 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 45.040 8.205 45.360 ;
      LAYER met4 ;
        RECT 7.885 45.040 8.205 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 44.610 8.205 44.930 ;
      LAYER met4 ;
        RECT 7.885 44.610 8.205 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 44.180 8.205 44.500 ;
      LAYER met4 ;
        RECT 7.885 44.180 8.205 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 43.750 8.205 44.070 ;
      LAYER met4 ;
        RECT 7.885 43.750 8.205 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 43.320 8.205 43.640 ;
      LAYER met4 ;
        RECT 7.885 43.320 8.205 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 42.890 8.205 43.210 ;
      LAYER met4 ;
        RECT 7.885 42.890 8.205 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 42.460 8.205 42.780 ;
      LAYER met4 ;
        RECT 7.885 42.460 8.205 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 42.030 8.205 42.350 ;
      LAYER met4 ;
        RECT 7.885 42.030 8.205 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.885 41.600 8.205 41.920 ;
      LAYER met4 ;
        RECT 7.885 41.600 8.205 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 45.900 7.800 46.220 ;
      LAYER met4 ;
        RECT 7.480 45.900 7.800 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 45.470 7.800 45.790 ;
      LAYER met4 ;
        RECT 7.480 45.470 7.800 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 45.040 7.800 45.360 ;
      LAYER met4 ;
        RECT 7.480 45.040 7.800 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 44.610 7.800 44.930 ;
      LAYER met4 ;
        RECT 7.480 44.610 7.800 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 44.180 7.800 44.500 ;
      LAYER met4 ;
        RECT 7.480 44.180 7.800 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 43.750 7.800 44.070 ;
      LAYER met4 ;
        RECT 7.480 43.750 7.800 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 43.320 7.800 43.640 ;
      LAYER met4 ;
        RECT 7.480 43.320 7.800 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 42.890 7.800 43.210 ;
      LAYER met4 ;
        RECT 7.480 42.890 7.800 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 42.460 7.800 42.780 ;
      LAYER met4 ;
        RECT 7.480 42.460 7.800 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 42.030 7.800 42.350 ;
      LAYER met4 ;
        RECT 7.480 42.030 7.800 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.480 41.600 7.800 41.920 ;
      LAYER met4 ;
        RECT 7.480 41.600 7.800 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 45.900 7.395 46.220 ;
      LAYER met4 ;
        RECT 7.075 45.900 7.395 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 45.470 7.395 45.790 ;
      LAYER met4 ;
        RECT 7.075 45.470 7.395 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 45.040 7.395 45.360 ;
      LAYER met4 ;
        RECT 7.075 45.040 7.395 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 44.610 7.395 44.930 ;
      LAYER met4 ;
        RECT 7.075 44.610 7.395 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 44.180 7.395 44.500 ;
      LAYER met4 ;
        RECT 7.075 44.180 7.395 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 43.750 7.395 44.070 ;
      LAYER met4 ;
        RECT 7.075 43.750 7.395 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 43.320 7.395 43.640 ;
      LAYER met4 ;
        RECT 7.075 43.320 7.395 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 42.890 7.395 43.210 ;
      LAYER met4 ;
        RECT 7.075 42.890 7.395 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 42.460 7.395 42.780 ;
      LAYER met4 ;
        RECT 7.075 42.460 7.395 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 42.030 7.395 42.350 ;
      LAYER met4 ;
        RECT 7.075 42.030 7.395 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.075 41.600 7.395 41.920 ;
      LAYER met4 ;
        RECT 7.075 41.600 7.395 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 45.900 6.990 46.220 ;
      LAYER met4 ;
        RECT 6.670 45.900 6.990 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 45.470 6.990 45.790 ;
      LAYER met4 ;
        RECT 6.670 45.470 6.990 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 45.040 6.990 45.360 ;
      LAYER met4 ;
        RECT 6.670 45.040 6.990 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 44.610 6.990 44.930 ;
      LAYER met4 ;
        RECT 6.670 44.610 6.990 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 44.180 6.990 44.500 ;
      LAYER met4 ;
        RECT 6.670 44.180 6.990 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 43.750 6.990 44.070 ;
      LAYER met4 ;
        RECT 6.670 43.750 6.990 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 43.320 6.990 43.640 ;
      LAYER met4 ;
        RECT 6.670 43.320 6.990 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 42.890 6.990 43.210 ;
      LAYER met4 ;
        RECT 6.670 42.890 6.990 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 42.460 6.990 42.780 ;
      LAYER met4 ;
        RECT 6.670 42.460 6.990 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 42.030 6.990 42.350 ;
      LAYER met4 ;
        RECT 6.670 42.030 6.990 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.670 41.600 6.990 41.920 ;
      LAYER met4 ;
        RECT 6.670 41.600 6.990 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 45.900 6.585 46.220 ;
      LAYER met4 ;
        RECT 6.265 45.900 6.585 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 45.470 6.585 45.790 ;
      LAYER met4 ;
        RECT 6.265 45.470 6.585 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 45.040 6.585 45.360 ;
      LAYER met4 ;
        RECT 6.265 45.040 6.585 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 44.610 6.585 44.930 ;
      LAYER met4 ;
        RECT 6.265 44.610 6.585 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 44.180 6.585 44.500 ;
      LAYER met4 ;
        RECT 6.265 44.180 6.585 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 43.750 6.585 44.070 ;
      LAYER met4 ;
        RECT 6.265 43.750 6.585 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 43.320 6.585 43.640 ;
      LAYER met4 ;
        RECT 6.265 43.320 6.585 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 42.890 6.585 43.210 ;
      LAYER met4 ;
        RECT 6.265 42.890 6.585 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 42.460 6.585 42.780 ;
      LAYER met4 ;
        RECT 6.265 42.460 6.585 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 42.030 6.585 42.350 ;
      LAYER met4 ;
        RECT 6.265 42.030 6.585 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.265 41.600 6.585 41.920 ;
      LAYER met4 ;
        RECT 6.265 41.600 6.585 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 45.900 6.180 46.220 ;
      LAYER met4 ;
        RECT 5.860 45.900 6.180 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 45.470 6.180 45.790 ;
      LAYER met4 ;
        RECT 5.860 45.470 6.180 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 45.040 6.180 45.360 ;
      LAYER met4 ;
        RECT 5.860 45.040 6.180 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 44.610 6.180 44.930 ;
      LAYER met4 ;
        RECT 5.860 44.610 6.180 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 44.180 6.180 44.500 ;
      LAYER met4 ;
        RECT 5.860 44.180 6.180 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 43.750 6.180 44.070 ;
      LAYER met4 ;
        RECT 5.860 43.750 6.180 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 43.320 6.180 43.640 ;
      LAYER met4 ;
        RECT 5.860 43.320 6.180 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 42.890 6.180 43.210 ;
      LAYER met4 ;
        RECT 5.860 42.890 6.180 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 42.460 6.180 42.780 ;
      LAYER met4 ;
        RECT 5.860 42.460 6.180 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 42.030 6.180 42.350 ;
      LAYER met4 ;
        RECT 5.860 42.030 6.180 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.860 41.600 6.180 41.920 ;
      LAYER met4 ;
        RECT 5.860 41.600 6.180 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 45.900 5.775 46.220 ;
      LAYER met4 ;
        RECT 5.455 45.900 5.775 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 45.470 5.775 45.790 ;
      LAYER met4 ;
        RECT 5.455 45.470 5.775 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 45.040 5.775 45.360 ;
      LAYER met4 ;
        RECT 5.455 45.040 5.775 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 44.610 5.775 44.930 ;
      LAYER met4 ;
        RECT 5.455 44.610 5.775 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 44.180 5.775 44.500 ;
      LAYER met4 ;
        RECT 5.455 44.180 5.775 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 43.750 5.775 44.070 ;
      LAYER met4 ;
        RECT 5.455 43.750 5.775 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 43.320 5.775 43.640 ;
      LAYER met4 ;
        RECT 5.455 43.320 5.775 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 42.890 5.775 43.210 ;
      LAYER met4 ;
        RECT 5.455 42.890 5.775 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 42.460 5.775 42.780 ;
      LAYER met4 ;
        RECT 5.455 42.460 5.775 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 42.030 5.775 42.350 ;
      LAYER met4 ;
        RECT 5.455 42.030 5.775 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.455 41.600 5.775 41.920 ;
      LAYER met4 ;
        RECT 5.455 41.600 5.775 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 45.900 5.370 46.220 ;
      LAYER met4 ;
        RECT 5.050 45.900 5.370 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 45.470 5.370 45.790 ;
      LAYER met4 ;
        RECT 5.050 45.470 5.370 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 45.040 5.370 45.360 ;
      LAYER met4 ;
        RECT 5.050 45.040 5.370 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 44.610 5.370 44.930 ;
      LAYER met4 ;
        RECT 5.050 44.610 5.370 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 44.180 5.370 44.500 ;
      LAYER met4 ;
        RECT 5.050 44.180 5.370 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 43.750 5.370 44.070 ;
      LAYER met4 ;
        RECT 5.050 43.750 5.370 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 43.320 5.370 43.640 ;
      LAYER met4 ;
        RECT 5.050 43.320 5.370 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 42.890 5.370 43.210 ;
      LAYER met4 ;
        RECT 5.050 42.890 5.370 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 42.460 5.370 42.780 ;
      LAYER met4 ;
        RECT 5.050 42.460 5.370 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 42.030 5.370 42.350 ;
      LAYER met4 ;
        RECT 5.050 42.030 5.370 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.050 41.600 5.370 41.920 ;
      LAYER met4 ;
        RECT 5.050 41.600 5.370 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 45.900 4.965 46.220 ;
      LAYER met4 ;
        RECT 4.645 45.900 4.965 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 45.470 4.965 45.790 ;
      LAYER met4 ;
        RECT 4.645 45.470 4.965 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 45.040 4.965 45.360 ;
      LAYER met4 ;
        RECT 4.645 45.040 4.965 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 44.610 4.965 44.930 ;
      LAYER met4 ;
        RECT 4.645 44.610 4.965 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 44.180 4.965 44.500 ;
      LAYER met4 ;
        RECT 4.645 44.180 4.965 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 43.750 4.965 44.070 ;
      LAYER met4 ;
        RECT 4.645 43.750 4.965 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 43.320 4.965 43.640 ;
      LAYER met4 ;
        RECT 4.645 43.320 4.965 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 42.890 4.965 43.210 ;
      LAYER met4 ;
        RECT 4.645 42.890 4.965 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 42.460 4.965 42.780 ;
      LAYER met4 ;
        RECT 4.645 42.460 4.965 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 42.030 4.965 42.350 ;
      LAYER met4 ;
        RECT 4.645 42.030 4.965 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.645 41.600 4.965 41.920 ;
      LAYER met4 ;
        RECT 4.645 41.600 4.965 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 45.900 4.560 46.220 ;
      LAYER met4 ;
        RECT 4.240 45.900 4.560 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 45.470 4.560 45.790 ;
      LAYER met4 ;
        RECT 4.240 45.470 4.560 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 45.040 4.560 45.360 ;
      LAYER met4 ;
        RECT 4.240 45.040 4.560 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 44.610 4.560 44.930 ;
      LAYER met4 ;
        RECT 4.240 44.610 4.560 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 44.180 4.560 44.500 ;
      LAYER met4 ;
        RECT 4.240 44.180 4.560 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 43.750 4.560 44.070 ;
      LAYER met4 ;
        RECT 4.240 43.750 4.560 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 43.320 4.560 43.640 ;
      LAYER met4 ;
        RECT 4.240 43.320 4.560 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 42.890 4.560 43.210 ;
      LAYER met4 ;
        RECT 4.240 42.890 4.560 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 42.460 4.560 42.780 ;
      LAYER met4 ;
        RECT 4.240 42.460 4.560 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 42.030 4.560 42.350 ;
      LAYER met4 ;
        RECT 4.240 42.030 4.560 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.240 41.600 4.560 41.920 ;
      LAYER met4 ;
        RECT 4.240 41.600 4.560 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 45.900 4.155 46.220 ;
      LAYER met4 ;
        RECT 3.835 45.900 4.155 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 45.470 4.155 45.790 ;
      LAYER met4 ;
        RECT 3.835 45.470 4.155 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 45.040 4.155 45.360 ;
      LAYER met4 ;
        RECT 3.835 45.040 4.155 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 44.610 4.155 44.930 ;
      LAYER met4 ;
        RECT 3.835 44.610 4.155 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 44.180 4.155 44.500 ;
      LAYER met4 ;
        RECT 3.835 44.180 4.155 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 43.750 4.155 44.070 ;
      LAYER met4 ;
        RECT 3.835 43.750 4.155 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 43.320 4.155 43.640 ;
      LAYER met4 ;
        RECT 3.835 43.320 4.155 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 42.890 4.155 43.210 ;
      LAYER met4 ;
        RECT 3.835 42.890 4.155 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 42.460 4.155 42.780 ;
      LAYER met4 ;
        RECT 3.835 42.460 4.155 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 42.030 4.155 42.350 ;
      LAYER met4 ;
        RECT 3.835 42.030 4.155 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.835 41.600 4.155 41.920 ;
      LAYER met4 ;
        RECT 3.835 41.600 4.155 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 45.900 3.750 46.220 ;
      LAYER met4 ;
        RECT 3.430 45.900 3.750 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 45.470 3.750 45.790 ;
      LAYER met4 ;
        RECT 3.430 45.470 3.750 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 45.040 3.750 45.360 ;
      LAYER met4 ;
        RECT 3.430 45.040 3.750 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 44.610 3.750 44.930 ;
      LAYER met4 ;
        RECT 3.430 44.610 3.750 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 44.180 3.750 44.500 ;
      LAYER met4 ;
        RECT 3.430 44.180 3.750 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 43.750 3.750 44.070 ;
      LAYER met4 ;
        RECT 3.430 43.750 3.750 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 43.320 3.750 43.640 ;
      LAYER met4 ;
        RECT 3.430 43.320 3.750 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 42.890 3.750 43.210 ;
      LAYER met4 ;
        RECT 3.430 42.890 3.750 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 42.460 3.750 42.780 ;
      LAYER met4 ;
        RECT 3.430 42.460 3.750 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 42.030 3.750 42.350 ;
      LAYER met4 ;
        RECT 3.430 42.030 3.750 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.430 41.600 3.750 41.920 ;
      LAYER met4 ;
        RECT 3.430 41.600 3.750 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 45.900 3.345 46.220 ;
      LAYER met4 ;
        RECT 3.025 45.900 3.345 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 45.470 3.345 45.790 ;
      LAYER met4 ;
        RECT 3.025 45.470 3.345 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 45.040 3.345 45.360 ;
      LAYER met4 ;
        RECT 3.025 45.040 3.345 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 44.610 3.345 44.930 ;
      LAYER met4 ;
        RECT 3.025 44.610 3.345 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 44.180 3.345 44.500 ;
      LAYER met4 ;
        RECT 3.025 44.180 3.345 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 43.750 3.345 44.070 ;
      LAYER met4 ;
        RECT 3.025 43.750 3.345 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 43.320 3.345 43.640 ;
      LAYER met4 ;
        RECT 3.025 43.320 3.345 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 42.890 3.345 43.210 ;
      LAYER met4 ;
        RECT 3.025 42.890 3.345 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 42.460 3.345 42.780 ;
      LAYER met4 ;
        RECT 3.025 42.460 3.345 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 42.030 3.345 42.350 ;
      LAYER met4 ;
        RECT 3.025 42.030 3.345 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 41.600 3.345 41.920 ;
      LAYER met4 ;
        RECT 3.025 41.600 3.345 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 45.900 2.940 46.220 ;
      LAYER met4 ;
        RECT 2.620 45.900 2.940 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 45.470 2.940 45.790 ;
      LAYER met4 ;
        RECT 2.620 45.470 2.940 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 45.040 2.940 45.360 ;
      LAYER met4 ;
        RECT 2.620 45.040 2.940 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 44.610 2.940 44.930 ;
      LAYER met4 ;
        RECT 2.620 44.610 2.940 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 44.180 2.940 44.500 ;
      LAYER met4 ;
        RECT 2.620 44.180 2.940 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 43.750 2.940 44.070 ;
      LAYER met4 ;
        RECT 2.620 43.750 2.940 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 43.320 2.940 43.640 ;
      LAYER met4 ;
        RECT 2.620 43.320 2.940 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 42.890 2.940 43.210 ;
      LAYER met4 ;
        RECT 2.620 42.890 2.940 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 42.460 2.940 42.780 ;
      LAYER met4 ;
        RECT 2.620 42.460 2.940 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 42.030 2.940 42.350 ;
      LAYER met4 ;
        RECT 2.620 42.030 2.940 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.620 41.600 2.940 41.920 ;
      LAYER met4 ;
        RECT 2.620 41.600 2.940 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 45.900 2.535 46.220 ;
      LAYER met4 ;
        RECT 2.215 45.900 2.535 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 45.470 2.535 45.790 ;
      LAYER met4 ;
        RECT 2.215 45.470 2.535 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 45.040 2.535 45.360 ;
      LAYER met4 ;
        RECT 2.215 45.040 2.535 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 44.610 2.535 44.930 ;
      LAYER met4 ;
        RECT 2.215 44.610 2.535 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 44.180 2.535 44.500 ;
      LAYER met4 ;
        RECT 2.215 44.180 2.535 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 43.750 2.535 44.070 ;
      LAYER met4 ;
        RECT 2.215 43.750 2.535 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 43.320 2.535 43.640 ;
      LAYER met4 ;
        RECT 2.215 43.320 2.535 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 42.890 2.535 43.210 ;
      LAYER met4 ;
        RECT 2.215 42.890 2.535 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 42.460 2.535 42.780 ;
      LAYER met4 ;
        RECT 2.215 42.460 2.535 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 42.030 2.535 42.350 ;
      LAYER met4 ;
        RECT 2.215 42.030 2.535 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.215 41.600 2.535 41.920 ;
      LAYER met4 ;
        RECT 2.215 41.600 2.535 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 45.900 2.130 46.220 ;
      LAYER met4 ;
        RECT 1.810 45.900 2.130 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 45.470 2.130 45.790 ;
      LAYER met4 ;
        RECT 1.810 45.470 2.130 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 45.040 2.130 45.360 ;
      LAYER met4 ;
        RECT 1.810 45.040 2.130 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 44.610 2.130 44.930 ;
      LAYER met4 ;
        RECT 1.810 44.610 2.130 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 44.180 2.130 44.500 ;
      LAYER met4 ;
        RECT 1.810 44.180 2.130 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 43.750 2.130 44.070 ;
      LAYER met4 ;
        RECT 1.810 43.750 2.130 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 43.320 2.130 43.640 ;
      LAYER met4 ;
        RECT 1.810 43.320 2.130 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 42.890 2.130 43.210 ;
      LAYER met4 ;
        RECT 1.810 42.890 2.130 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 42.460 2.130 42.780 ;
      LAYER met4 ;
        RECT 1.810 42.460 2.130 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 42.030 2.130 42.350 ;
      LAYER met4 ;
        RECT 1.810 42.030 2.130 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.810 41.600 2.130 41.920 ;
      LAYER met4 ;
        RECT 1.810 41.600 2.130 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 45.900 1.725 46.220 ;
      LAYER met4 ;
        RECT 1.405 45.900 1.725 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 45.470 1.725 45.790 ;
      LAYER met4 ;
        RECT 1.405 45.470 1.725 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 45.040 1.725 45.360 ;
      LAYER met4 ;
        RECT 1.405 45.040 1.725 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 44.610 1.725 44.930 ;
      LAYER met4 ;
        RECT 1.405 44.610 1.725 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 44.180 1.725 44.500 ;
      LAYER met4 ;
        RECT 1.405 44.180 1.725 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 43.750 1.725 44.070 ;
      LAYER met4 ;
        RECT 1.405 43.750 1.725 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 43.320 1.725 43.640 ;
      LAYER met4 ;
        RECT 1.405 43.320 1.725 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 42.890 1.725 43.210 ;
      LAYER met4 ;
        RECT 1.405 42.890 1.725 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 42.460 1.725 42.780 ;
      LAYER met4 ;
        RECT 1.405 42.460 1.725 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 42.030 1.725 42.350 ;
      LAYER met4 ;
        RECT 1.405 42.030 1.725 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 41.600 1.725 41.920 ;
      LAYER met4 ;
        RECT 1.405 41.600 1.725 41.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 45.900 1.320 46.220 ;
      LAYER met4 ;
        RECT 1.270 45.900 1.320 46.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 45.470 1.320 45.790 ;
      LAYER met4 ;
        RECT 1.270 45.470 1.320 45.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 45.040 1.320 45.360 ;
      LAYER met4 ;
        RECT 1.270 45.040 1.320 45.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 44.610 1.320 44.930 ;
      LAYER met4 ;
        RECT 1.270 44.610 1.320 44.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 44.180 1.320 44.500 ;
      LAYER met4 ;
        RECT 1.270 44.180 1.320 44.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 43.750 1.320 44.070 ;
      LAYER met4 ;
        RECT 1.270 43.750 1.320 44.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 43.320 1.320 43.640 ;
      LAYER met4 ;
        RECT 1.270 43.320 1.320 43.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 42.890 1.320 43.210 ;
      LAYER met4 ;
        RECT 1.270 42.890 1.320 43.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 42.460 1.320 42.780 ;
      LAYER met4 ;
        RECT 1.270 42.460 1.320 42.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 42.030 1.320 42.350 ;
      LAYER met4 ;
        RECT 1.270 42.030 1.320 42.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 41.600 1.320 41.920 ;
      LAYER met4 ;
        RECT 1.270 41.600 1.320 41.920 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
  END VSWITCH
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.970 41.590 24.395 46.230 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 96.585 75.000 174.185 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__overlay_vssd_hvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vssd_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vssd_lvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
  END VSSA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
  END VDDIO_Q
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 39.590 74.700 44.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 43.960 74.610 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 43.530 74.610 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 43.100 74.610 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 42.670 74.610 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 42.240 74.610 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 41.810 74.610 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 41.380 74.610 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 40.950 74.610 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 40.520 74.610 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 40.090 74.610 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.410 39.660 74.610 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 43.960 74.205 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 43.530 74.205 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 43.100 74.205 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 42.670 74.205 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 42.240 74.205 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 41.810 74.205 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 41.380 74.205 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 40.950 74.205 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 40.520 74.205 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 40.090 74.205 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.005 39.660 74.205 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 43.960 73.800 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 43.530 73.800 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 43.100 73.800 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 42.670 73.800 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 42.240 73.800 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 41.810 73.800 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 41.380 73.800 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 40.950 73.800 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 40.520 73.800 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 40.090 73.800 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.600 39.660 73.800 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 43.960 73.395 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 43.530 73.395 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 43.100 73.395 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 42.670 73.395 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 42.240 73.395 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 41.810 73.395 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 41.380 73.395 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 40.950 73.395 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 40.520 73.395 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 40.090 73.395 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.195 39.660 73.395 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 43.960 72.990 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 43.530 72.990 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 43.100 72.990 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 42.670 72.990 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 42.240 72.990 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 41.810 72.990 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 41.380 72.990 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 40.950 72.990 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 40.520 72.990 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 40.090 72.990 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.790 39.660 72.990 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 43.960 72.585 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 43.530 72.585 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 43.100 72.585 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 42.670 72.585 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 42.240 72.585 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 41.810 72.585 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 41.380 72.585 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 40.950 72.585 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 40.520 72.585 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 40.090 72.585 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.385 39.660 72.585 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 43.960 72.180 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 43.530 72.180 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 43.100 72.180 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 42.670 72.180 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 42.240 72.180 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 41.810 72.180 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 41.380 72.180 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 40.950 72.180 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 40.520 72.180 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 40.090 72.180 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 39.660 72.180 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 43.960 71.775 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 43.530 71.775 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 43.100 71.775 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 42.670 71.775 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 42.240 71.775 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 41.810 71.775 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 41.380 71.775 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 40.950 71.775 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 40.520 71.775 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 40.090 71.775 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.575 39.660 71.775 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 43.960 71.370 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 43.530 71.370 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 43.100 71.370 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 42.670 71.370 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 42.240 71.370 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 41.810 71.370 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 41.380 71.370 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 40.950 71.370 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 40.520 71.370 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 40.090 71.370 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.170 39.660 71.370 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 43.960 70.965 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 43.530 70.965 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 43.100 70.965 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 42.670 70.965 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 42.240 70.965 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 41.810 70.965 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 41.380 70.965 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 40.950 70.965 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 40.520 70.965 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 40.090 70.965 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.765 39.660 70.965 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 43.960 70.560 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 43.530 70.560 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 43.100 70.560 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 42.670 70.560 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 42.240 70.560 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 41.810 70.560 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 41.380 70.560 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 40.950 70.560 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 40.520 70.560 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 40.090 70.560 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.360 39.660 70.560 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 43.960 70.155 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 43.530 70.155 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 43.100 70.155 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 42.670 70.155 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 42.240 70.155 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 41.810 70.155 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 41.380 70.155 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 40.950 70.155 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 40.520 70.155 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 40.090 70.155 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.955 39.660 70.155 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 43.960 69.750 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 43.530 69.750 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 43.100 69.750 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 42.670 69.750 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 42.240 69.750 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 41.810 69.750 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 41.380 69.750 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 40.950 69.750 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 40.520 69.750 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 40.090 69.750 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.550 39.660 69.750 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 43.960 69.345 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 43.530 69.345 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 43.100 69.345 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 42.670 69.345 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 42.240 69.345 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 41.810 69.345 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 41.380 69.345 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 40.950 69.345 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 40.520 69.345 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 40.090 69.345 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.145 39.660 69.345 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 43.960 68.940 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 43.530 68.940 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 43.100 68.940 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 42.670 68.940 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 42.240 68.940 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 41.810 68.940 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 41.380 68.940 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 40.950 68.940 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 40.520 68.940 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 40.090 68.940 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.740 39.660 68.940 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 43.960 68.535 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 43.530 68.535 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 43.100 68.535 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 42.670 68.535 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 42.240 68.535 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 41.810 68.535 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 41.380 68.535 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 40.950 68.535 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 40.520 68.535 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 40.090 68.535 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.335 39.660 68.535 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 43.960 68.130 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 43.530 68.130 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 43.100 68.130 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 42.670 68.130 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 42.240 68.130 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 41.810 68.130 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 41.380 68.130 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 40.950 68.130 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 40.520 68.130 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 40.090 68.130 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 39.660 68.130 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 43.960 67.725 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 43.530 67.725 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 43.100 67.725 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 42.670 67.725 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 42.240 67.725 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 41.810 67.725 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 41.380 67.725 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 40.950 67.725 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 40.520 67.725 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 40.090 67.725 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.525 39.660 67.725 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 43.960 67.320 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 43.530 67.320 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 43.100 67.320 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 42.670 67.320 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 42.240 67.320 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 41.810 67.320 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 41.380 67.320 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 40.950 67.320 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 40.520 67.320 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 40.090 67.320 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.120 39.660 67.320 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 43.960 66.915 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 43.530 66.915 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 43.100 66.915 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 42.670 66.915 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 42.240 66.915 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 41.810 66.915 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 41.380 66.915 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 40.950 66.915 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 40.520 66.915 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 40.090 66.915 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.715 39.660 66.915 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 43.960 66.510 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 43.530 66.510 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 43.100 66.510 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 42.670 66.510 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 42.240 66.510 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 41.810 66.510 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 41.380 66.510 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 40.950 66.510 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 40.520 66.510 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 40.090 66.510 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.310 39.660 66.510 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 43.960 66.105 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 43.530 66.105 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 43.100 66.105 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 42.670 66.105 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 42.240 66.105 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 41.810 66.105 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 41.380 66.105 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 40.950 66.105 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 40.520 66.105 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 40.090 66.105 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.905 39.660 66.105 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 43.960 65.700 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 43.530 65.700 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 43.100 65.700 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 42.670 65.700 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 42.240 65.700 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 41.810 65.700 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 41.380 65.700 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 40.950 65.700 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 40.520 65.700 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 40.090 65.700 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.500 39.660 65.700 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 43.960 65.295 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 43.530 65.295 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 43.100 65.295 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 42.670 65.295 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 42.240 65.295 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 41.810 65.295 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 41.380 65.295 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 40.950 65.295 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 40.520 65.295 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 40.090 65.295 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.095 39.660 65.295 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 43.960 64.890 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 43.530 64.890 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 43.100 64.890 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 42.670 64.890 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 42.240 64.890 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 41.810 64.890 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 41.380 64.890 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 40.950 64.890 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 40.520 64.890 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 40.090 64.890 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.690 39.660 64.890 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 43.960 64.485 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 43.530 64.485 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 43.100 64.485 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 42.670 64.485 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 42.240 64.485 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 41.810 64.485 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 41.380 64.485 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 40.950 64.485 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 40.520 64.485 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 40.090 64.485 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.285 39.660 64.485 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 43.960 64.080 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 43.530 64.080 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 43.100 64.080 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 42.670 64.080 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 42.240 64.080 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 41.810 64.080 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 41.380 64.080 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 40.950 64.080 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 40.520 64.080 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 40.090 64.080 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.880 39.660 64.080 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 43.960 63.675 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 43.530 63.675 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 43.100 63.675 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 42.670 63.675 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 42.240 63.675 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 41.810 63.675 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 41.380 63.675 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 40.950 63.675 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 40.520 63.675 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 40.090 63.675 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.475 39.660 63.675 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 43.960 63.270 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 43.530 63.270 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 43.100 63.270 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 42.670 63.270 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 42.240 63.270 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 41.810 63.270 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 41.380 63.270 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 40.950 63.270 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 40.520 63.270 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 40.090 63.270 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.070 39.660 63.270 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 43.960 62.865 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 43.530 62.865 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 43.100 62.865 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 42.670 62.865 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 42.240 62.865 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 41.810 62.865 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 41.380 62.865 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 40.950 62.865 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 40.520 62.865 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 40.090 62.865 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.665 39.660 62.865 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 43.960 62.460 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 43.530 62.460 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 43.100 62.460 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 42.670 62.460 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 42.240 62.460 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 41.810 62.460 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 41.380 62.460 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 40.950 62.460 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 40.520 62.460 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 40.090 62.460 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.260 39.660 62.460 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 43.960 62.055 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 43.530 62.055 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 43.100 62.055 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 42.670 62.055 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 42.240 62.055 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 41.810 62.055 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 41.380 62.055 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 40.950 62.055 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 40.520 62.055 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 40.090 62.055 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.855 39.660 62.055 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 43.960 61.650 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 43.530 61.650 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 43.100 61.650 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 42.670 61.650 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 42.240 61.650 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 41.810 61.650 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 41.380 61.650 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 40.950 61.650 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 40.520 61.650 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 40.090 61.650 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.450 39.660 61.650 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 43.960 61.245 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 43.530 61.245 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 43.100 61.245 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 42.670 61.245 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 42.240 61.245 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 41.810 61.245 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 41.380 61.245 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 40.950 61.245 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 40.520 61.245 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 40.090 61.245 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.045 39.660 61.245 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 43.960 60.840 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 43.530 60.840 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 43.100 60.840 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 42.670 60.840 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 42.240 60.840 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 41.810 60.840 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 41.380 60.840 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 40.950 60.840 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 40.520 60.840 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 40.090 60.840 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.640 39.660 60.840 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 43.960 60.435 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 43.530 60.435 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 43.100 60.435 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 42.670 60.435 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 42.240 60.435 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 41.810 60.435 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 41.380 60.435 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 40.950 60.435 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 40.520 60.435 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 40.090 60.435 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.235 39.660 60.435 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 43.960 60.030 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 43.530 60.030 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 43.100 60.030 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 42.670 60.030 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 42.240 60.030 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 41.810 60.030 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 41.380 60.030 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 40.950 60.030 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 40.520 60.030 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 40.090 60.030 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.830 39.660 60.030 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 43.960 59.625 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 43.530 59.625 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 43.100 59.625 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 42.670 59.625 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 42.240 59.625 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 41.810 59.625 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 41.380 59.625 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 40.950 59.625 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 40.520 59.625 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 40.090 59.625 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 39.660 59.625 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 43.960 59.220 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 43.530 59.220 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 43.100 59.220 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 42.670 59.220 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 42.240 59.220 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 41.810 59.220 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 41.380 59.220 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 40.950 59.220 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 40.520 59.220 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 40.090 59.220 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.020 39.660 59.220 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 43.960 58.815 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 43.530 58.815 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 43.100 58.815 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 42.670 58.815 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 42.240 58.815 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 41.810 58.815 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 41.380 58.815 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 40.950 58.815 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 40.520 58.815 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 40.090 58.815 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.615 39.660 58.815 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 43.960 58.410 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 43.530 58.410 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 43.100 58.410 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 42.670 58.410 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 42.240 58.410 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 41.810 58.410 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 41.380 58.410 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 40.950 58.410 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 40.520 58.410 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 40.090 58.410 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.210 39.660 58.410 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 43.960 58.005 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 43.530 58.005 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 43.100 58.005 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 42.670 58.005 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 42.240 58.005 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 41.810 58.005 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 41.380 58.005 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 40.950 58.005 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 40.520 58.005 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 40.090 58.005 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.805 39.660 58.005 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 43.960 57.600 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 43.530 57.600 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 43.100 57.600 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 42.670 57.600 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 42.240 57.600 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 41.810 57.600 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 41.380 57.600 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 40.950 57.600 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 40.520 57.600 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 40.090 57.600 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.400 39.660 57.600 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 43.960 57.195 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 43.530 57.195 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 43.100 57.195 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 42.670 57.195 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 42.240 57.195 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 41.810 57.195 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 41.380 57.195 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 40.950 57.195 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 40.520 57.195 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 40.090 57.195 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.995 39.660 57.195 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 43.960 56.785 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 43.530 56.785 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 43.100 56.785 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 42.670 56.785 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 42.240 56.785 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 41.810 56.785 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 41.380 56.785 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 40.950 56.785 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 40.520 56.785 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 40.090 56.785 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 39.660 56.785 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 43.960 56.375 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 43.530 56.375 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 43.100 56.375 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 42.670 56.375 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 42.240 56.375 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 41.810 56.375 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 41.380 56.375 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 40.950 56.375 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 40.520 56.375 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 40.090 56.375 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 39.660 56.375 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 43.960 55.965 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 43.530 55.965 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 43.100 55.965 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 42.670 55.965 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 42.240 55.965 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 41.810 55.965 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 41.380 55.965 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 40.950 55.965 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 40.520 55.965 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 40.090 55.965 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 39.660 55.965 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 43.960 55.555 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 43.530 55.555 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 43.100 55.555 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 42.670 55.555 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 42.240 55.555 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 41.810 55.555 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 41.380 55.555 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 40.950 55.555 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 40.520 55.555 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 40.090 55.555 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 39.660 55.555 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 43.960 55.145 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 43.530 55.145 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 43.100 55.145 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 42.670 55.145 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 42.240 55.145 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 41.810 55.145 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 41.380 55.145 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 40.950 55.145 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 40.520 55.145 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 40.090 55.145 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 39.660 55.145 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 43.960 54.735 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 43.530 54.735 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 43.100 54.735 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 42.670 54.735 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 42.240 54.735 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 41.810 54.735 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 41.380 54.735 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 40.950 54.735 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 40.520 54.735 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 40.090 54.735 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 39.660 54.735 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 43.960 54.325 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 43.530 54.325 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 43.100 54.325 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 42.670 54.325 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 42.240 54.325 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 41.810 54.325 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 41.380 54.325 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 40.950 54.325 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 40.520 54.325 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 40.090 54.325 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 39.660 54.325 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 43.960 53.915 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 43.530 53.915 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 43.100 53.915 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 42.670 53.915 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 42.240 53.915 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 41.810 53.915 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 41.380 53.915 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 40.950 53.915 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 40.520 53.915 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 40.090 53.915 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 39.660 53.915 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 43.960 53.505 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 43.530 53.505 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 43.100 53.505 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 42.670 53.505 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 42.240 53.505 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 41.810 53.505 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 41.380 53.505 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 40.950 53.505 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 40.520 53.505 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 40.090 53.505 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 39.660 53.505 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 43.960 53.095 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 43.530 53.095 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 43.100 53.095 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 42.670 53.095 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 42.240 53.095 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 41.810 53.095 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 41.380 53.095 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 40.950 53.095 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 40.520 53.095 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 40.090 53.095 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 39.660 53.095 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 43.960 52.685 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 43.530 52.685 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 43.100 52.685 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 42.670 52.685 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 42.240 52.685 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 41.810 52.685 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 41.380 52.685 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 40.950 52.685 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 40.520 52.685 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 40.090 52.685 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 39.660 52.685 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 43.960 52.275 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 43.530 52.275 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 43.100 52.275 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 42.670 52.275 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 42.240 52.275 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 41.810 52.275 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 41.380 52.275 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 40.950 52.275 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 40.520 52.275 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 40.090 52.275 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 39.660 52.275 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 43.960 51.865 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 43.530 51.865 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 43.100 51.865 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 42.670 51.865 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 42.240 51.865 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 41.810 51.865 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 41.380 51.865 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 40.950 51.865 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 40.520 51.865 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 40.090 51.865 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 39.660 51.865 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 43.960 51.455 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 43.530 51.455 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 43.100 51.455 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 42.670 51.455 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 42.240 51.455 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 41.810 51.455 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 41.380 51.455 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 40.950 51.455 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 40.520 51.455 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 40.090 51.455 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 39.660 51.455 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 43.960 51.045 44.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 43.530 51.045 43.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 43.100 51.045 43.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 42.670 51.045 42.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 42.240 51.045 42.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 41.810 51.045 42.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 41.380 51.045 41.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 40.950 51.045 41.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 40.520 51.045 40.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 40.090 51.045 40.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 39.660 51.045 39.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 43.900 24.470 44.220 ;
      LAYER met4 ;
        RECT 24.150 43.900 24.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 43.470 24.470 43.790 ;
      LAYER met4 ;
        RECT 24.150 43.470 24.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 43.040 24.470 43.360 ;
      LAYER met4 ;
        RECT 24.150 43.040 24.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 42.610 24.470 42.930 ;
      LAYER met4 ;
        RECT 24.150 42.610 24.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 42.180 24.470 42.500 ;
      LAYER met4 ;
        RECT 24.150 42.180 24.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 41.750 24.470 42.070 ;
      LAYER met4 ;
        RECT 24.150 41.750 24.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 41.320 24.470 41.640 ;
      LAYER met4 ;
        RECT 24.150 41.320 24.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 40.890 24.470 41.210 ;
      LAYER met4 ;
        RECT 24.150 40.890 24.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 40.460 24.470 40.780 ;
      LAYER met4 ;
        RECT 24.150 40.460 24.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 40.030 24.470 40.350 ;
      LAYER met4 ;
        RECT 24.150 40.030 24.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.150 39.600 24.470 39.920 ;
      LAYER met4 ;
        RECT 24.150 39.600 24.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 43.900 24.070 44.220 ;
      LAYER met4 ;
        RECT 23.750 43.900 24.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 43.470 24.070 43.790 ;
      LAYER met4 ;
        RECT 23.750 43.470 24.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 43.040 24.070 43.360 ;
      LAYER met4 ;
        RECT 23.750 43.040 24.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 42.610 24.070 42.930 ;
      LAYER met4 ;
        RECT 23.750 42.610 24.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 42.180 24.070 42.500 ;
      LAYER met4 ;
        RECT 23.750 42.180 24.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 41.750 24.070 42.070 ;
      LAYER met4 ;
        RECT 23.750 41.750 24.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 41.320 24.070 41.640 ;
      LAYER met4 ;
        RECT 23.750 41.320 24.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 40.890 24.070 41.210 ;
      LAYER met4 ;
        RECT 23.750 40.890 24.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 40.460 24.070 40.780 ;
      LAYER met4 ;
        RECT 23.750 40.460 24.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 40.030 24.070 40.350 ;
      LAYER met4 ;
        RECT 23.750 40.030 24.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.750 39.600 24.070 39.920 ;
      LAYER met4 ;
        RECT 23.750 39.600 24.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 43.900 23.670 44.220 ;
      LAYER met4 ;
        RECT 23.350 43.900 23.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 43.470 23.670 43.790 ;
      LAYER met4 ;
        RECT 23.350 43.470 23.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 43.040 23.670 43.360 ;
      LAYER met4 ;
        RECT 23.350 43.040 23.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 42.610 23.670 42.930 ;
      LAYER met4 ;
        RECT 23.350 42.610 23.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 42.180 23.670 42.500 ;
      LAYER met4 ;
        RECT 23.350 42.180 23.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 41.750 23.670 42.070 ;
      LAYER met4 ;
        RECT 23.350 41.750 23.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 41.320 23.670 41.640 ;
      LAYER met4 ;
        RECT 23.350 41.320 23.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 40.890 23.670 41.210 ;
      LAYER met4 ;
        RECT 23.350 40.890 23.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 40.460 23.670 40.780 ;
      LAYER met4 ;
        RECT 23.350 40.460 23.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 40.030 23.670 40.350 ;
      LAYER met4 ;
        RECT 23.350 40.030 23.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.350 39.600 23.670 39.920 ;
      LAYER met4 ;
        RECT 23.350 39.600 23.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 43.900 23.270 44.220 ;
      LAYER met4 ;
        RECT 22.950 43.900 23.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 43.470 23.270 43.790 ;
      LAYER met4 ;
        RECT 22.950 43.470 23.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 43.040 23.270 43.360 ;
      LAYER met4 ;
        RECT 22.950 43.040 23.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 42.610 23.270 42.930 ;
      LAYER met4 ;
        RECT 22.950 42.610 23.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 42.180 23.270 42.500 ;
      LAYER met4 ;
        RECT 22.950 42.180 23.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 41.750 23.270 42.070 ;
      LAYER met4 ;
        RECT 22.950 41.750 23.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 41.320 23.270 41.640 ;
      LAYER met4 ;
        RECT 22.950 41.320 23.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 40.890 23.270 41.210 ;
      LAYER met4 ;
        RECT 22.950 40.890 23.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 40.460 23.270 40.780 ;
      LAYER met4 ;
        RECT 22.950 40.460 23.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 40.030 23.270 40.350 ;
      LAYER met4 ;
        RECT 22.950 40.030 23.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 39.600 23.270 39.920 ;
      LAYER met4 ;
        RECT 22.950 39.600 23.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 43.900 22.870 44.220 ;
      LAYER met4 ;
        RECT 22.550 43.900 22.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 43.470 22.870 43.790 ;
      LAYER met4 ;
        RECT 22.550 43.470 22.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 43.040 22.870 43.360 ;
      LAYER met4 ;
        RECT 22.550 43.040 22.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 42.610 22.870 42.930 ;
      LAYER met4 ;
        RECT 22.550 42.610 22.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 42.180 22.870 42.500 ;
      LAYER met4 ;
        RECT 22.550 42.180 22.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 41.750 22.870 42.070 ;
      LAYER met4 ;
        RECT 22.550 41.750 22.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 41.320 22.870 41.640 ;
      LAYER met4 ;
        RECT 22.550 41.320 22.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 40.890 22.870 41.210 ;
      LAYER met4 ;
        RECT 22.550 40.890 22.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 40.460 22.870 40.780 ;
      LAYER met4 ;
        RECT 22.550 40.460 22.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 40.030 22.870 40.350 ;
      LAYER met4 ;
        RECT 22.550 40.030 22.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.550 39.600 22.870 39.920 ;
      LAYER met4 ;
        RECT 22.550 39.600 22.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 43.900 22.470 44.220 ;
      LAYER met4 ;
        RECT 22.150 43.900 22.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 43.470 22.470 43.790 ;
      LAYER met4 ;
        RECT 22.150 43.470 22.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 43.040 22.470 43.360 ;
      LAYER met4 ;
        RECT 22.150 43.040 22.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 42.610 22.470 42.930 ;
      LAYER met4 ;
        RECT 22.150 42.610 22.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 42.180 22.470 42.500 ;
      LAYER met4 ;
        RECT 22.150 42.180 22.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 41.750 22.470 42.070 ;
      LAYER met4 ;
        RECT 22.150 41.750 22.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 41.320 22.470 41.640 ;
      LAYER met4 ;
        RECT 22.150 41.320 22.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 40.890 22.470 41.210 ;
      LAYER met4 ;
        RECT 22.150 40.890 22.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 40.460 22.470 40.780 ;
      LAYER met4 ;
        RECT 22.150 40.460 22.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 40.030 22.470 40.350 ;
      LAYER met4 ;
        RECT 22.150 40.030 22.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.150 39.600 22.470 39.920 ;
      LAYER met4 ;
        RECT 22.150 39.600 22.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 43.900 22.070 44.220 ;
      LAYER met4 ;
        RECT 21.750 43.900 22.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 43.470 22.070 43.790 ;
      LAYER met4 ;
        RECT 21.750 43.470 22.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 43.040 22.070 43.360 ;
      LAYER met4 ;
        RECT 21.750 43.040 22.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 42.610 22.070 42.930 ;
      LAYER met4 ;
        RECT 21.750 42.610 22.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 42.180 22.070 42.500 ;
      LAYER met4 ;
        RECT 21.750 42.180 22.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 41.750 22.070 42.070 ;
      LAYER met4 ;
        RECT 21.750 41.750 22.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 41.320 22.070 41.640 ;
      LAYER met4 ;
        RECT 21.750 41.320 22.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 40.890 22.070 41.210 ;
      LAYER met4 ;
        RECT 21.750 40.890 22.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 40.460 22.070 40.780 ;
      LAYER met4 ;
        RECT 21.750 40.460 22.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 40.030 22.070 40.350 ;
      LAYER met4 ;
        RECT 21.750 40.030 22.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.750 39.600 22.070 39.920 ;
      LAYER met4 ;
        RECT 21.750 39.600 22.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 43.900 21.670 44.220 ;
      LAYER met4 ;
        RECT 21.350 43.900 21.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 43.470 21.670 43.790 ;
      LAYER met4 ;
        RECT 21.350 43.470 21.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 43.040 21.670 43.360 ;
      LAYER met4 ;
        RECT 21.350 43.040 21.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 42.610 21.670 42.930 ;
      LAYER met4 ;
        RECT 21.350 42.610 21.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 42.180 21.670 42.500 ;
      LAYER met4 ;
        RECT 21.350 42.180 21.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 41.750 21.670 42.070 ;
      LAYER met4 ;
        RECT 21.350 41.750 21.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 41.320 21.670 41.640 ;
      LAYER met4 ;
        RECT 21.350 41.320 21.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 40.890 21.670 41.210 ;
      LAYER met4 ;
        RECT 21.350 40.890 21.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 40.460 21.670 40.780 ;
      LAYER met4 ;
        RECT 21.350 40.460 21.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 40.030 21.670 40.350 ;
      LAYER met4 ;
        RECT 21.350 40.030 21.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.350 39.600 21.670 39.920 ;
      LAYER met4 ;
        RECT 21.350 39.600 21.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 43.900 21.270 44.220 ;
      LAYER met4 ;
        RECT 20.950 43.900 21.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 43.470 21.270 43.790 ;
      LAYER met4 ;
        RECT 20.950 43.470 21.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 43.040 21.270 43.360 ;
      LAYER met4 ;
        RECT 20.950 43.040 21.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 42.610 21.270 42.930 ;
      LAYER met4 ;
        RECT 20.950 42.610 21.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 42.180 21.270 42.500 ;
      LAYER met4 ;
        RECT 20.950 42.180 21.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 41.750 21.270 42.070 ;
      LAYER met4 ;
        RECT 20.950 41.750 21.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 41.320 21.270 41.640 ;
      LAYER met4 ;
        RECT 20.950 41.320 21.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 40.890 21.270 41.210 ;
      LAYER met4 ;
        RECT 20.950 40.890 21.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 40.460 21.270 40.780 ;
      LAYER met4 ;
        RECT 20.950 40.460 21.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 40.030 21.270 40.350 ;
      LAYER met4 ;
        RECT 20.950 40.030 21.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.950 39.600 21.270 39.920 ;
      LAYER met4 ;
        RECT 20.950 39.600 21.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 43.900 20.870 44.220 ;
      LAYER met4 ;
        RECT 20.550 43.900 20.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 43.470 20.870 43.790 ;
      LAYER met4 ;
        RECT 20.550 43.470 20.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 43.040 20.870 43.360 ;
      LAYER met4 ;
        RECT 20.550 43.040 20.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 42.610 20.870 42.930 ;
      LAYER met4 ;
        RECT 20.550 42.610 20.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 42.180 20.870 42.500 ;
      LAYER met4 ;
        RECT 20.550 42.180 20.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 41.750 20.870 42.070 ;
      LAYER met4 ;
        RECT 20.550 41.750 20.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 41.320 20.870 41.640 ;
      LAYER met4 ;
        RECT 20.550 41.320 20.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 40.890 20.870 41.210 ;
      LAYER met4 ;
        RECT 20.550 40.890 20.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 40.460 20.870 40.780 ;
      LAYER met4 ;
        RECT 20.550 40.460 20.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 40.030 20.870 40.350 ;
      LAYER met4 ;
        RECT 20.550 40.030 20.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.550 39.600 20.870 39.920 ;
      LAYER met4 ;
        RECT 20.550 39.600 20.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 43.900 20.470 44.220 ;
      LAYER met4 ;
        RECT 20.150 43.900 20.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 43.470 20.470 43.790 ;
      LAYER met4 ;
        RECT 20.150 43.470 20.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 43.040 20.470 43.360 ;
      LAYER met4 ;
        RECT 20.150 43.040 20.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 42.610 20.470 42.930 ;
      LAYER met4 ;
        RECT 20.150 42.610 20.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 42.180 20.470 42.500 ;
      LAYER met4 ;
        RECT 20.150 42.180 20.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 41.750 20.470 42.070 ;
      LAYER met4 ;
        RECT 20.150 41.750 20.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 41.320 20.470 41.640 ;
      LAYER met4 ;
        RECT 20.150 41.320 20.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 40.890 20.470 41.210 ;
      LAYER met4 ;
        RECT 20.150 40.890 20.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 40.460 20.470 40.780 ;
      LAYER met4 ;
        RECT 20.150 40.460 20.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 40.030 20.470 40.350 ;
      LAYER met4 ;
        RECT 20.150 40.030 20.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.150 39.600 20.470 39.920 ;
      LAYER met4 ;
        RECT 20.150 39.600 20.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 43.900 20.070 44.220 ;
      LAYER met4 ;
        RECT 19.750 43.900 20.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 43.470 20.070 43.790 ;
      LAYER met4 ;
        RECT 19.750 43.470 20.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 43.040 20.070 43.360 ;
      LAYER met4 ;
        RECT 19.750 43.040 20.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 42.610 20.070 42.930 ;
      LAYER met4 ;
        RECT 19.750 42.610 20.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 42.180 20.070 42.500 ;
      LAYER met4 ;
        RECT 19.750 42.180 20.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 41.750 20.070 42.070 ;
      LAYER met4 ;
        RECT 19.750 41.750 20.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 41.320 20.070 41.640 ;
      LAYER met4 ;
        RECT 19.750 41.320 20.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 40.890 20.070 41.210 ;
      LAYER met4 ;
        RECT 19.750 40.890 20.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 40.460 20.070 40.780 ;
      LAYER met4 ;
        RECT 19.750 40.460 20.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 40.030 20.070 40.350 ;
      LAYER met4 ;
        RECT 19.750 40.030 20.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.750 39.600 20.070 39.920 ;
      LAYER met4 ;
        RECT 19.750 39.600 20.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 43.900 19.670 44.220 ;
      LAYER met4 ;
        RECT 19.350 43.900 19.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 43.470 19.670 43.790 ;
      LAYER met4 ;
        RECT 19.350 43.470 19.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 43.040 19.670 43.360 ;
      LAYER met4 ;
        RECT 19.350 43.040 19.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 42.610 19.670 42.930 ;
      LAYER met4 ;
        RECT 19.350 42.610 19.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 42.180 19.670 42.500 ;
      LAYER met4 ;
        RECT 19.350 42.180 19.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 41.750 19.670 42.070 ;
      LAYER met4 ;
        RECT 19.350 41.750 19.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 41.320 19.670 41.640 ;
      LAYER met4 ;
        RECT 19.350 41.320 19.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 40.890 19.670 41.210 ;
      LAYER met4 ;
        RECT 19.350 40.890 19.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 40.460 19.670 40.780 ;
      LAYER met4 ;
        RECT 19.350 40.460 19.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 40.030 19.670 40.350 ;
      LAYER met4 ;
        RECT 19.350 40.030 19.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.350 39.600 19.670 39.920 ;
      LAYER met4 ;
        RECT 19.350 39.600 19.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 43.900 19.270 44.220 ;
      LAYER met4 ;
        RECT 18.950 43.900 19.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 43.470 19.270 43.790 ;
      LAYER met4 ;
        RECT 18.950 43.470 19.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 43.040 19.270 43.360 ;
      LAYER met4 ;
        RECT 18.950 43.040 19.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 42.610 19.270 42.930 ;
      LAYER met4 ;
        RECT 18.950 42.610 19.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 42.180 19.270 42.500 ;
      LAYER met4 ;
        RECT 18.950 42.180 19.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 41.750 19.270 42.070 ;
      LAYER met4 ;
        RECT 18.950 41.750 19.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 41.320 19.270 41.640 ;
      LAYER met4 ;
        RECT 18.950 41.320 19.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 40.890 19.270 41.210 ;
      LAYER met4 ;
        RECT 18.950 40.890 19.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 40.460 19.270 40.780 ;
      LAYER met4 ;
        RECT 18.950 40.460 19.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 40.030 19.270 40.350 ;
      LAYER met4 ;
        RECT 18.950 40.030 19.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.950 39.600 19.270 39.920 ;
      LAYER met4 ;
        RECT 18.950 39.600 19.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 43.900 18.870 44.220 ;
      LAYER met4 ;
        RECT 18.550 43.900 18.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 43.470 18.870 43.790 ;
      LAYER met4 ;
        RECT 18.550 43.470 18.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 43.040 18.870 43.360 ;
      LAYER met4 ;
        RECT 18.550 43.040 18.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 42.610 18.870 42.930 ;
      LAYER met4 ;
        RECT 18.550 42.610 18.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 42.180 18.870 42.500 ;
      LAYER met4 ;
        RECT 18.550 42.180 18.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 41.750 18.870 42.070 ;
      LAYER met4 ;
        RECT 18.550 41.750 18.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 41.320 18.870 41.640 ;
      LAYER met4 ;
        RECT 18.550 41.320 18.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 40.890 18.870 41.210 ;
      LAYER met4 ;
        RECT 18.550 40.890 18.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 40.460 18.870 40.780 ;
      LAYER met4 ;
        RECT 18.550 40.460 18.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 40.030 18.870 40.350 ;
      LAYER met4 ;
        RECT 18.550 40.030 18.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.550 39.600 18.870 39.920 ;
      LAYER met4 ;
        RECT 18.550 39.600 18.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 43.900 18.470 44.220 ;
      LAYER met4 ;
        RECT 18.150 43.900 18.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 43.470 18.470 43.790 ;
      LAYER met4 ;
        RECT 18.150 43.470 18.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 43.040 18.470 43.360 ;
      LAYER met4 ;
        RECT 18.150 43.040 18.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 42.610 18.470 42.930 ;
      LAYER met4 ;
        RECT 18.150 42.610 18.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 42.180 18.470 42.500 ;
      LAYER met4 ;
        RECT 18.150 42.180 18.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 41.750 18.470 42.070 ;
      LAYER met4 ;
        RECT 18.150 41.750 18.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 41.320 18.470 41.640 ;
      LAYER met4 ;
        RECT 18.150 41.320 18.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 40.890 18.470 41.210 ;
      LAYER met4 ;
        RECT 18.150 40.890 18.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 40.460 18.470 40.780 ;
      LAYER met4 ;
        RECT 18.150 40.460 18.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 40.030 18.470 40.350 ;
      LAYER met4 ;
        RECT 18.150 40.030 18.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.150 39.600 18.470 39.920 ;
      LAYER met4 ;
        RECT 18.150 39.600 18.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 43.900 18.070 44.220 ;
      LAYER met4 ;
        RECT 17.750 43.900 18.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 43.470 18.070 43.790 ;
      LAYER met4 ;
        RECT 17.750 43.470 18.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 43.040 18.070 43.360 ;
      LAYER met4 ;
        RECT 17.750 43.040 18.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 42.610 18.070 42.930 ;
      LAYER met4 ;
        RECT 17.750 42.610 18.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 42.180 18.070 42.500 ;
      LAYER met4 ;
        RECT 17.750 42.180 18.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 41.750 18.070 42.070 ;
      LAYER met4 ;
        RECT 17.750 41.750 18.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 41.320 18.070 41.640 ;
      LAYER met4 ;
        RECT 17.750 41.320 18.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 40.890 18.070 41.210 ;
      LAYER met4 ;
        RECT 17.750 40.890 18.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 40.460 18.070 40.780 ;
      LAYER met4 ;
        RECT 17.750 40.460 18.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 40.030 18.070 40.350 ;
      LAYER met4 ;
        RECT 17.750 40.030 18.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.750 39.600 18.070 39.920 ;
      LAYER met4 ;
        RECT 17.750 39.600 18.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 43.900 17.670 44.220 ;
      LAYER met4 ;
        RECT 17.350 43.900 17.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 43.470 17.670 43.790 ;
      LAYER met4 ;
        RECT 17.350 43.470 17.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 43.040 17.670 43.360 ;
      LAYER met4 ;
        RECT 17.350 43.040 17.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 42.610 17.670 42.930 ;
      LAYER met4 ;
        RECT 17.350 42.610 17.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 42.180 17.670 42.500 ;
      LAYER met4 ;
        RECT 17.350 42.180 17.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 41.750 17.670 42.070 ;
      LAYER met4 ;
        RECT 17.350 41.750 17.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 41.320 17.670 41.640 ;
      LAYER met4 ;
        RECT 17.350 41.320 17.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 40.890 17.670 41.210 ;
      LAYER met4 ;
        RECT 17.350 40.890 17.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 40.460 17.670 40.780 ;
      LAYER met4 ;
        RECT 17.350 40.460 17.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 40.030 17.670 40.350 ;
      LAYER met4 ;
        RECT 17.350 40.030 17.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.350 39.600 17.670 39.920 ;
      LAYER met4 ;
        RECT 17.350 39.600 17.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 43.900 17.270 44.220 ;
      LAYER met4 ;
        RECT 16.950 43.900 17.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 43.470 17.270 43.790 ;
      LAYER met4 ;
        RECT 16.950 43.470 17.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 43.040 17.270 43.360 ;
      LAYER met4 ;
        RECT 16.950 43.040 17.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 42.610 17.270 42.930 ;
      LAYER met4 ;
        RECT 16.950 42.610 17.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 42.180 17.270 42.500 ;
      LAYER met4 ;
        RECT 16.950 42.180 17.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 41.750 17.270 42.070 ;
      LAYER met4 ;
        RECT 16.950 41.750 17.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 41.320 17.270 41.640 ;
      LAYER met4 ;
        RECT 16.950 41.320 17.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 40.890 17.270 41.210 ;
      LAYER met4 ;
        RECT 16.950 40.890 17.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 40.460 17.270 40.780 ;
      LAYER met4 ;
        RECT 16.950 40.460 17.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 40.030 17.270 40.350 ;
      LAYER met4 ;
        RECT 16.950 40.030 17.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.950 39.600 17.270 39.920 ;
      LAYER met4 ;
        RECT 16.950 39.600 17.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 43.900 16.870 44.220 ;
      LAYER met4 ;
        RECT 16.550 43.900 16.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 43.470 16.870 43.790 ;
      LAYER met4 ;
        RECT 16.550 43.470 16.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 43.040 16.870 43.360 ;
      LAYER met4 ;
        RECT 16.550 43.040 16.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 42.610 16.870 42.930 ;
      LAYER met4 ;
        RECT 16.550 42.610 16.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 42.180 16.870 42.500 ;
      LAYER met4 ;
        RECT 16.550 42.180 16.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 41.750 16.870 42.070 ;
      LAYER met4 ;
        RECT 16.550 41.750 16.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 41.320 16.870 41.640 ;
      LAYER met4 ;
        RECT 16.550 41.320 16.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 40.890 16.870 41.210 ;
      LAYER met4 ;
        RECT 16.550 40.890 16.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 40.460 16.870 40.780 ;
      LAYER met4 ;
        RECT 16.550 40.460 16.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 40.030 16.870 40.350 ;
      LAYER met4 ;
        RECT 16.550 40.030 16.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.550 39.600 16.870 39.920 ;
      LAYER met4 ;
        RECT 16.550 39.600 16.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 43.900 16.470 44.220 ;
      LAYER met4 ;
        RECT 16.150 43.900 16.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 43.470 16.470 43.790 ;
      LAYER met4 ;
        RECT 16.150 43.470 16.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 43.040 16.470 43.360 ;
      LAYER met4 ;
        RECT 16.150 43.040 16.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 42.610 16.470 42.930 ;
      LAYER met4 ;
        RECT 16.150 42.610 16.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 42.180 16.470 42.500 ;
      LAYER met4 ;
        RECT 16.150 42.180 16.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 41.750 16.470 42.070 ;
      LAYER met4 ;
        RECT 16.150 41.750 16.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 41.320 16.470 41.640 ;
      LAYER met4 ;
        RECT 16.150 41.320 16.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 40.890 16.470 41.210 ;
      LAYER met4 ;
        RECT 16.150 40.890 16.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 40.460 16.470 40.780 ;
      LAYER met4 ;
        RECT 16.150 40.460 16.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 40.030 16.470 40.350 ;
      LAYER met4 ;
        RECT 16.150 40.030 16.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.150 39.600 16.470 39.920 ;
      LAYER met4 ;
        RECT 16.150 39.600 16.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 43.900 16.070 44.220 ;
      LAYER met4 ;
        RECT 15.750 43.900 16.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 43.470 16.070 43.790 ;
      LAYER met4 ;
        RECT 15.750 43.470 16.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 43.040 16.070 43.360 ;
      LAYER met4 ;
        RECT 15.750 43.040 16.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 42.610 16.070 42.930 ;
      LAYER met4 ;
        RECT 15.750 42.610 16.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 42.180 16.070 42.500 ;
      LAYER met4 ;
        RECT 15.750 42.180 16.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 41.750 16.070 42.070 ;
      LAYER met4 ;
        RECT 15.750 41.750 16.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 41.320 16.070 41.640 ;
      LAYER met4 ;
        RECT 15.750 41.320 16.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 40.890 16.070 41.210 ;
      LAYER met4 ;
        RECT 15.750 40.890 16.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 40.460 16.070 40.780 ;
      LAYER met4 ;
        RECT 15.750 40.460 16.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 40.030 16.070 40.350 ;
      LAYER met4 ;
        RECT 15.750 40.030 16.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.750 39.600 16.070 39.920 ;
      LAYER met4 ;
        RECT 15.750 39.600 16.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 43.900 15.670 44.220 ;
      LAYER met4 ;
        RECT 15.350 43.900 15.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 43.470 15.670 43.790 ;
      LAYER met4 ;
        RECT 15.350 43.470 15.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 43.040 15.670 43.360 ;
      LAYER met4 ;
        RECT 15.350 43.040 15.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 42.610 15.670 42.930 ;
      LAYER met4 ;
        RECT 15.350 42.610 15.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 42.180 15.670 42.500 ;
      LAYER met4 ;
        RECT 15.350 42.180 15.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 41.750 15.670 42.070 ;
      LAYER met4 ;
        RECT 15.350 41.750 15.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 41.320 15.670 41.640 ;
      LAYER met4 ;
        RECT 15.350 41.320 15.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 40.890 15.670 41.210 ;
      LAYER met4 ;
        RECT 15.350 40.890 15.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 40.460 15.670 40.780 ;
      LAYER met4 ;
        RECT 15.350 40.460 15.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 40.030 15.670 40.350 ;
      LAYER met4 ;
        RECT 15.350 40.030 15.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.350 39.600 15.670 39.920 ;
      LAYER met4 ;
        RECT 15.350 39.600 15.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 43.900 15.270 44.220 ;
      LAYER met4 ;
        RECT 14.950 43.900 15.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 43.470 15.270 43.790 ;
      LAYER met4 ;
        RECT 14.950 43.470 15.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 43.040 15.270 43.360 ;
      LAYER met4 ;
        RECT 14.950 43.040 15.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 42.610 15.270 42.930 ;
      LAYER met4 ;
        RECT 14.950 42.610 15.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 42.180 15.270 42.500 ;
      LAYER met4 ;
        RECT 14.950 42.180 15.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 41.750 15.270 42.070 ;
      LAYER met4 ;
        RECT 14.950 41.750 15.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 41.320 15.270 41.640 ;
      LAYER met4 ;
        RECT 14.950 41.320 15.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 40.890 15.270 41.210 ;
      LAYER met4 ;
        RECT 14.950 40.890 15.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 40.460 15.270 40.780 ;
      LAYER met4 ;
        RECT 14.950 40.460 15.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 40.030 15.270 40.350 ;
      LAYER met4 ;
        RECT 14.950 40.030 15.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.950 39.600 15.270 39.920 ;
      LAYER met4 ;
        RECT 14.950 39.600 15.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 43.900 14.870 44.220 ;
      LAYER met4 ;
        RECT 14.550 43.900 14.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 43.470 14.870 43.790 ;
      LAYER met4 ;
        RECT 14.550 43.470 14.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 43.040 14.870 43.360 ;
      LAYER met4 ;
        RECT 14.550 43.040 14.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 42.610 14.870 42.930 ;
      LAYER met4 ;
        RECT 14.550 42.610 14.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 42.180 14.870 42.500 ;
      LAYER met4 ;
        RECT 14.550 42.180 14.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 41.750 14.870 42.070 ;
      LAYER met4 ;
        RECT 14.550 41.750 14.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 41.320 14.870 41.640 ;
      LAYER met4 ;
        RECT 14.550 41.320 14.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 40.890 14.870 41.210 ;
      LAYER met4 ;
        RECT 14.550 40.890 14.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 40.460 14.870 40.780 ;
      LAYER met4 ;
        RECT 14.550 40.460 14.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 40.030 14.870 40.350 ;
      LAYER met4 ;
        RECT 14.550 40.030 14.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.550 39.600 14.870 39.920 ;
      LAYER met4 ;
        RECT 14.550 39.600 14.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 43.900 14.470 44.220 ;
      LAYER met4 ;
        RECT 14.150 43.900 14.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 43.470 14.470 43.790 ;
      LAYER met4 ;
        RECT 14.150 43.470 14.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 43.040 14.470 43.360 ;
      LAYER met4 ;
        RECT 14.150 43.040 14.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 42.610 14.470 42.930 ;
      LAYER met4 ;
        RECT 14.150 42.610 14.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 42.180 14.470 42.500 ;
      LAYER met4 ;
        RECT 14.150 42.180 14.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 41.750 14.470 42.070 ;
      LAYER met4 ;
        RECT 14.150 41.750 14.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 41.320 14.470 41.640 ;
      LAYER met4 ;
        RECT 14.150 41.320 14.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 40.890 14.470 41.210 ;
      LAYER met4 ;
        RECT 14.150 40.890 14.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 40.460 14.470 40.780 ;
      LAYER met4 ;
        RECT 14.150 40.460 14.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 40.030 14.470 40.350 ;
      LAYER met4 ;
        RECT 14.150 40.030 14.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.150 39.600 14.470 39.920 ;
      LAYER met4 ;
        RECT 14.150 39.600 14.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 43.900 14.070 44.220 ;
      LAYER met4 ;
        RECT 13.750 43.900 14.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 43.470 14.070 43.790 ;
      LAYER met4 ;
        RECT 13.750 43.470 14.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 43.040 14.070 43.360 ;
      LAYER met4 ;
        RECT 13.750 43.040 14.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 42.610 14.070 42.930 ;
      LAYER met4 ;
        RECT 13.750 42.610 14.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 42.180 14.070 42.500 ;
      LAYER met4 ;
        RECT 13.750 42.180 14.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 41.750 14.070 42.070 ;
      LAYER met4 ;
        RECT 13.750 41.750 14.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 41.320 14.070 41.640 ;
      LAYER met4 ;
        RECT 13.750 41.320 14.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 40.890 14.070 41.210 ;
      LAYER met4 ;
        RECT 13.750 40.890 14.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 40.460 14.070 40.780 ;
      LAYER met4 ;
        RECT 13.750 40.460 14.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 40.030 14.070 40.350 ;
      LAYER met4 ;
        RECT 13.750 40.030 14.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.750 39.600 14.070 39.920 ;
      LAYER met4 ;
        RECT 13.750 39.600 14.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 43.900 13.670 44.220 ;
      LAYER met4 ;
        RECT 13.350 43.900 13.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 43.470 13.670 43.790 ;
      LAYER met4 ;
        RECT 13.350 43.470 13.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 43.040 13.670 43.360 ;
      LAYER met4 ;
        RECT 13.350 43.040 13.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 42.610 13.670 42.930 ;
      LAYER met4 ;
        RECT 13.350 42.610 13.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 42.180 13.670 42.500 ;
      LAYER met4 ;
        RECT 13.350 42.180 13.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 41.750 13.670 42.070 ;
      LAYER met4 ;
        RECT 13.350 41.750 13.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 41.320 13.670 41.640 ;
      LAYER met4 ;
        RECT 13.350 41.320 13.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 40.890 13.670 41.210 ;
      LAYER met4 ;
        RECT 13.350 40.890 13.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 40.460 13.670 40.780 ;
      LAYER met4 ;
        RECT 13.350 40.460 13.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 40.030 13.670 40.350 ;
      LAYER met4 ;
        RECT 13.350 40.030 13.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.350 39.600 13.670 39.920 ;
      LAYER met4 ;
        RECT 13.350 39.600 13.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 43.900 13.270 44.220 ;
      LAYER met4 ;
        RECT 12.950 43.900 13.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 43.470 13.270 43.790 ;
      LAYER met4 ;
        RECT 12.950 43.470 13.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 43.040 13.270 43.360 ;
      LAYER met4 ;
        RECT 12.950 43.040 13.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 42.610 13.270 42.930 ;
      LAYER met4 ;
        RECT 12.950 42.610 13.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 42.180 13.270 42.500 ;
      LAYER met4 ;
        RECT 12.950 42.180 13.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 41.750 13.270 42.070 ;
      LAYER met4 ;
        RECT 12.950 41.750 13.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 41.320 13.270 41.640 ;
      LAYER met4 ;
        RECT 12.950 41.320 13.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 40.890 13.270 41.210 ;
      LAYER met4 ;
        RECT 12.950 40.890 13.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 40.460 13.270 40.780 ;
      LAYER met4 ;
        RECT 12.950 40.460 13.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 40.030 13.270 40.350 ;
      LAYER met4 ;
        RECT 12.950 40.030 13.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.950 39.600 13.270 39.920 ;
      LAYER met4 ;
        RECT 12.950 39.600 13.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 43.900 12.870 44.220 ;
      LAYER met4 ;
        RECT 12.550 43.900 12.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 43.470 12.870 43.790 ;
      LAYER met4 ;
        RECT 12.550 43.470 12.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 43.040 12.870 43.360 ;
      LAYER met4 ;
        RECT 12.550 43.040 12.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 42.610 12.870 42.930 ;
      LAYER met4 ;
        RECT 12.550 42.610 12.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 42.180 12.870 42.500 ;
      LAYER met4 ;
        RECT 12.550 42.180 12.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 41.750 12.870 42.070 ;
      LAYER met4 ;
        RECT 12.550 41.750 12.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 41.320 12.870 41.640 ;
      LAYER met4 ;
        RECT 12.550 41.320 12.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 40.890 12.870 41.210 ;
      LAYER met4 ;
        RECT 12.550 40.890 12.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 40.460 12.870 40.780 ;
      LAYER met4 ;
        RECT 12.550 40.460 12.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 40.030 12.870 40.350 ;
      LAYER met4 ;
        RECT 12.550 40.030 12.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.550 39.600 12.870 39.920 ;
      LAYER met4 ;
        RECT 12.550 39.600 12.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 43.900 12.470 44.220 ;
      LAYER met4 ;
        RECT 12.150 43.900 12.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 43.470 12.470 43.790 ;
      LAYER met4 ;
        RECT 12.150 43.470 12.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 43.040 12.470 43.360 ;
      LAYER met4 ;
        RECT 12.150 43.040 12.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 42.610 12.470 42.930 ;
      LAYER met4 ;
        RECT 12.150 42.610 12.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 42.180 12.470 42.500 ;
      LAYER met4 ;
        RECT 12.150 42.180 12.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 41.750 12.470 42.070 ;
      LAYER met4 ;
        RECT 12.150 41.750 12.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 41.320 12.470 41.640 ;
      LAYER met4 ;
        RECT 12.150 41.320 12.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 40.890 12.470 41.210 ;
      LAYER met4 ;
        RECT 12.150 40.890 12.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 40.460 12.470 40.780 ;
      LAYER met4 ;
        RECT 12.150 40.460 12.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 40.030 12.470 40.350 ;
      LAYER met4 ;
        RECT 12.150 40.030 12.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.150 39.600 12.470 39.920 ;
      LAYER met4 ;
        RECT 12.150 39.600 12.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 43.900 12.070 44.220 ;
      LAYER met4 ;
        RECT 11.750 43.900 12.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 43.470 12.070 43.790 ;
      LAYER met4 ;
        RECT 11.750 43.470 12.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 43.040 12.070 43.360 ;
      LAYER met4 ;
        RECT 11.750 43.040 12.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 42.610 12.070 42.930 ;
      LAYER met4 ;
        RECT 11.750 42.610 12.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 42.180 12.070 42.500 ;
      LAYER met4 ;
        RECT 11.750 42.180 12.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 41.750 12.070 42.070 ;
      LAYER met4 ;
        RECT 11.750 41.750 12.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 41.320 12.070 41.640 ;
      LAYER met4 ;
        RECT 11.750 41.320 12.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 40.890 12.070 41.210 ;
      LAYER met4 ;
        RECT 11.750 40.890 12.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 40.460 12.070 40.780 ;
      LAYER met4 ;
        RECT 11.750 40.460 12.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 40.030 12.070 40.350 ;
      LAYER met4 ;
        RECT 11.750 40.030 12.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.750 39.600 12.070 39.920 ;
      LAYER met4 ;
        RECT 11.750 39.600 12.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 43.900 11.670 44.220 ;
      LAYER met4 ;
        RECT 11.350 43.900 11.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 43.470 11.670 43.790 ;
      LAYER met4 ;
        RECT 11.350 43.470 11.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 43.040 11.670 43.360 ;
      LAYER met4 ;
        RECT 11.350 43.040 11.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 42.610 11.670 42.930 ;
      LAYER met4 ;
        RECT 11.350 42.610 11.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 42.180 11.670 42.500 ;
      LAYER met4 ;
        RECT 11.350 42.180 11.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 41.750 11.670 42.070 ;
      LAYER met4 ;
        RECT 11.350 41.750 11.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 41.320 11.670 41.640 ;
      LAYER met4 ;
        RECT 11.350 41.320 11.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 40.890 11.670 41.210 ;
      LAYER met4 ;
        RECT 11.350 40.890 11.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 40.460 11.670 40.780 ;
      LAYER met4 ;
        RECT 11.350 40.460 11.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 40.030 11.670 40.350 ;
      LAYER met4 ;
        RECT 11.350 40.030 11.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.350 39.600 11.670 39.920 ;
      LAYER met4 ;
        RECT 11.350 39.600 11.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 43.900 11.270 44.220 ;
      LAYER met4 ;
        RECT 10.950 43.900 11.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 43.470 11.270 43.790 ;
      LAYER met4 ;
        RECT 10.950 43.470 11.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 43.040 11.270 43.360 ;
      LAYER met4 ;
        RECT 10.950 43.040 11.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 42.610 11.270 42.930 ;
      LAYER met4 ;
        RECT 10.950 42.610 11.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 42.180 11.270 42.500 ;
      LAYER met4 ;
        RECT 10.950 42.180 11.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 41.750 11.270 42.070 ;
      LAYER met4 ;
        RECT 10.950 41.750 11.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 41.320 11.270 41.640 ;
      LAYER met4 ;
        RECT 10.950 41.320 11.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 40.890 11.270 41.210 ;
      LAYER met4 ;
        RECT 10.950 40.890 11.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 40.460 11.270 40.780 ;
      LAYER met4 ;
        RECT 10.950 40.460 11.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 40.030 11.270 40.350 ;
      LAYER met4 ;
        RECT 10.950 40.030 11.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.950 39.600 11.270 39.920 ;
      LAYER met4 ;
        RECT 10.950 39.600 11.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 43.900 10.870 44.220 ;
      LAYER met4 ;
        RECT 10.550 43.900 10.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 43.470 10.870 43.790 ;
      LAYER met4 ;
        RECT 10.550 43.470 10.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 43.040 10.870 43.360 ;
      LAYER met4 ;
        RECT 10.550 43.040 10.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 42.610 10.870 42.930 ;
      LAYER met4 ;
        RECT 10.550 42.610 10.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 42.180 10.870 42.500 ;
      LAYER met4 ;
        RECT 10.550 42.180 10.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 41.750 10.870 42.070 ;
      LAYER met4 ;
        RECT 10.550 41.750 10.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 41.320 10.870 41.640 ;
      LAYER met4 ;
        RECT 10.550 41.320 10.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 40.890 10.870 41.210 ;
      LAYER met4 ;
        RECT 10.550 40.890 10.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 40.460 10.870 40.780 ;
      LAYER met4 ;
        RECT 10.550 40.460 10.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 40.030 10.870 40.350 ;
      LAYER met4 ;
        RECT 10.550 40.030 10.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 39.600 10.870 39.920 ;
      LAYER met4 ;
        RECT 10.550 39.600 10.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 43.900 10.470 44.220 ;
      LAYER met4 ;
        RECT 10.150 43.900 10.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 43.470 10.470 43.790 ;
      LAYER met4 ;
        RECT 10.150 43.470 10.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 43.040 10.470 43.360 ;
      LAYER met4 ;
        RECT 10.150 43.040 10.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 42.610 10.470 42.930 ;
      LAYER met4 ;
        RECT 10.150 42.610 10.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 42.180 10.470 42.500 ;
      LAYER met4 ;
        RECT 10.150 42.180 10.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 41.750 10.470 42.070 ;
      LAYER met4 ;
        RECT 10.150 41.750 10.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 41.320 10.470 41.640 ;
      LAYER met4 ;
        RECT 10.150 41.320 10.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 40.890 10.470 41.210 ;
      LAYER met4 ;
        RECT 10.150 40.890 10.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 40.460 10.470 40.780 ;
      LAYER met4 ;
        RECT 10.150 40.460 10.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 40.030 10.470 40.350 ;
      LAYER met4 ;
        RECT 10.150 40.030 10.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.150 39.600 10.470 39.920 ;
      LAYER met4 ;
        RECT 10.150 39.600 10.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 43.900 10.070 44.220 ;
      LAYER met4 ;
        RECT 9.750 43.900 10.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 43.470 10.070 43.790 ;
      LAYER met4 ;
        RECT 9.750 43.470 10.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 43.040 10.070 43.360 ;
      LAYER met4 ;
        RECT 9.750 43.040 10.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 42.610 10.070 42.930 ;
      LAYER met4 ;
        RECT 9.750 42.610 10.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 42.180 10.070 42.500 ;
      LAYER met4 ;
        RECT 9.750 42.180 10.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 41.750 10.070 42.070 ;
      LAYER met4 ;
        RECT 9.750 41.750 10.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 41.320 10.070 41.640 ;
      LAYER met4 ;
        RECT 9.750 41.320 10.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 40.890 10.070 41.210 ;
      LAYER met4 ;
        RECT 9.750 40.890 10.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 40.460 10.070 40.780 ;
      LAYER met4 ;
        RECT 9.750 40.460 10.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 40.030 10.070 40.350 ;
      LAYER met4 ;
        RECT 9.750 40.030 10.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.750 39.600 10.070 39.920 ;
      LAYER met4 ;
        RECT 9.750 39.600 10.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 43.900 9.670 44.220 ;
      LAYER met4 ;
        RECT 9.350 43.900 9.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 43.470 9.670 43.790 ;
      LAYER met4 ;
        RECT 9.350 43.470 9.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 43.040 9.670 43.360 ;
      LAYER met4 ;
        RECT 9.350 43.040 9.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 42.610 9.670 42.930 ;
      LAYER met4 ;
        RECT 9.350 42.610 9.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 42.180 9.670 42.500 ;
      LAYER met4 ;
        RECT 9.350 42.180 9.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 41.750 9.670 42.070 ;
      LAYER met4 ;
        RECT 9.350 41.750 9.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 41.320 9.670 41.640 ;
      LAYER met4 ;
        RECT 9.350 41.320 9.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 40.890 9.670 41.210 ;
      LAYER met4 ;
        RECT 9.350 40.890 9.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 40.460 9.670 40.780 ;
      LAYER met4 ;
        RECT 9.350 40.460 9.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 40.030 9.670 40.350 ;
      LAYER met4 ;
        RECT 9.350 40.030 9.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.350 39.600 9.670 39.920 ;
      LAYER met4 ;
        RECT 9.350 39.600 9.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 43.900 9.270 44.220 ;
      LAYER met4 ;
        RECT 8.950 43.900 9.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 43.470 9.270 43.790 ;
      LAYER met4 ;
        RECT 8.950 43.470 9.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 43.040 9.270 43.360 ;
      LAYER met4 ;
        RECT 8.950 43.040 9.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 42.610 9.270 42.930 ;
      LAYER met4 ;
        RECT 8.950 42.610 9.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 42.180 9.270 42.500 ;
      LAYER met4 ;
        RECT 8.950 42.180 9.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 41.750 9.270 42.070 ;
      LAYER met4 ;
        RECT 8.950 41.750 9.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 41.320 9.270 41.640 ;
      LAYER met4 ;
        RECT 8.950 41.320 9.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 40.890 9.270 41.210 ;
      LAYER met4 ;
        RECT 8.950 40.890 9.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 40.460 9.270 40.780 ;
      LAYER met4 ;
        RECT 8.950 40.460 9.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 40.030 9.270 40.350 ;
      LAYER met4 ;
        RECT 8.950 40.030 9.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.950 39.600 9.270 39.920 ;
      LAYER met4 ;
        RECT 8.950 39.600 9.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 43.900 8.870 44.220 ;
      LAYER met4 ;
        RECT 8.550 43.900 8.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 43.470 8.870 43.790 ;
      LAYER met4 ;
        RECT 8.550 43.470 8.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 43.040 8.870 43.360 ;
      LAYER met4 ;
        RECT 8.550 43.040 8.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 42.610 8.870 42.930 ;
      LAYER met4 ;
        RECT 8.550 42.610 8.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 42.180 8.870 42.500 ;
      LAYER met4 ;
        RECT 8.550 42.180 8.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 41.750 8.870 42.070 ;
      LAYER met4 ;
        RECT 8.550 41.750 8.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 41.320 8.870 41.640 ;
      LAYER met4 ;
        RECT 8.550 41.320 8.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 40.890 8.870 41.210 ;
      LAYER met4 ;
        RECT 8.550 40.890 8.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 40.460 8.870 40.780 ;
      LAYER met4 ;
        RECT 8.550 40.460 8.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 40.030 8.870 40.350 ;
      LAYER met4 ;
        RECT 8.550 40.030 8.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.550 39.600 8.870 39.920 ;
      LAYER met4 ;
        RECT 8.550 39.600 8.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 43.900 8.470 44.220 ;
      LAYER met4 ;
        RECT 8.150 43.900 8.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 43.470 8.470 43.790 ;
      LAYER met4 ;
        RECT 8.150 43.470 8.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 43.040 8.470 43.360 ;
      LAYER met4 ;
        RECT 8.150 43.040 8.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 42.610 8.470 42.930 ;
      LAYER met4 ;
        RECT 8.150 42.610 8.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 42.180 8.470 42.500 ;
      LAYER met4 ;
        RECT 8.150 42.180 8.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 41.750 8.470 42.070 ;
      LAYER met4 ;
        RECT 8.150 41.750 8.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 41.320 8.470 41.640 ;
      LAYER met4 ;
        RECT 8.150 41.320 8.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 40.890 8.470 41.210 ;
      LAYER met4 ;
        RECT 8.150 40.890 8.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 40.460 8.470 40.780 ;
      LAYER met4 ;
        RECT 8.150 40.460 8.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 40.030 8.470 40.350 ;
      LAYER met4 ;
        RECT 8.150 40.030 8.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 39.600 8.470 39.920 ;
      LAYER met4 ;
        RECT 8.150 39.600 8.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 43.900 8.070 44.220 ;
      LAYER met4 ;
        RECT 7.750 43.900 8.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 43.470 8.070 43.790 ;
      LAYER met4 ;
        RECT 7.750 43.470 8.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 43.040 8.070 43.360 ;
      LAYER met4 ;
        RECT 7.750 43.040 8.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 42.610 8.070 42.930 ;
      LAYER met4 ;
        RECT 7.750 42.610 8.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 42.180 8.070 42.500 ;
      LAYER met4 ;
        RECT 7.750 42.180 8.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 41.750 8.070 42.070 ;
      LAYER met4 ;
        RECT 7.750 41.750 8.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 41.320 8.070 41.640 ;
      LAYER met4 ;
        RECT 7.750 41.320 8.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 40.890 8.070 41.210 ;
      LAYER met4 ;
        RECT 7.750 40.890 8.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 40.460 8.070 40.780 ;
      LAYER met4 ;
        RECT 7.750 40.460 8.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 40.030 8.070 40.350 ;
      LAYER met4 ;
        RECT 7.750 40.030 8.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.750 39.600 8.070 39.920 ;
      LAYER met4 ;
        RECT 7.750 39.600 8.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 43.900 7.670 44.220 ;
      LAYER met4 ;
        RECT 7.350 43.900 7.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 43.470 7.670 43.790 ;
      LAYER met4 ;
        RECT 7.350 43.470 7.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 43.040 7.670 43.360 ;
      LAYER met4 ;
        RECT 7.350 43.040 7.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 42.610 7.670 42.930 ;
      LAYER met4 ;
        RECT 7.350 42.610 7.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 42.180 7.670 42.500 ;
      LAYER met4 ;
        RECT 7.350 42.180 7.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 41.750 7.670 42.070 ;
      LAYER met4 ;
        RECT 7.350 41.750 7.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 41.320 7.670 41.640 ;
      LAYER met4 ;
        RECT 7.350 41.320 7.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 40.890 7.670 41.210 ;
      LAYER met4 ;
        RECT 7.350 40.890 7.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 40.460 7.670 40.780 ;
      LAYER met4 ;
        RECT 7.350 40.460 7.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 40.030 7.670 40.350 ;
      LAYER met4 ;
        RECT 7.350 40.030 7.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.350 39.600 7.670 39.920 ;
      LAYER met4 ;
        RECT 7.350 39.600 7.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 43.900 7.270 44.220 ;
      LAYER met4 ;
        RECT 6.950 43.900 7.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 43.470 7.270 43.790 ;
      LAYER met4 ;
        RECT 6.950 43.470 7.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 43.040 7.270 43.360 ;
      LAYER met4 ;
        RECT 6.950 43.040 7.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 42.610 7.270 42.930 ;
      LAYER met4 ;
        RECT 6.950 42.610 7.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 42.180 7.270 42.500 ;
      LAYER met4 ;
        RECT 6.950 42.180 7.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 41.750 7.270 42.070 ;
      LAYER met4 ;
        RECT 6.950 41.750 7.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 41.320 7.270 41.640 ;
      LAYER met4 ;
        RECT 6.950 41.320 7.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 40.890 7.270 41.210 ;
      LAYER met4 ;
        RECT 6.950 40.890 7.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 40.460 7.270 40.780 ;
      LAYER met4 ;
        RECT 6.950 40.460 7.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 40.030 7.270 40.350 ;
      LAYER met4 ;
        RECT 6.950 40.030 7.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.950 39.600 7.270 39.920 ;
      LAYER met4 ;
        RECT 6.950 39.600 7.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 43.900 6.870 44.220 ;
      LAYER met4 ;
        RECT 6.550 43.900 6.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 43.470 6.870 43.790 ;
      LAYER met4 ;
        RECT 6.550 43.470 6.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 43.040 6.870 43.360 ;
      LAYER met4 ;
        RECT 6.550 43.040 6.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 42.610 6.870 42.930 ;
      LAYER met4 ;
        RECT 6.550 42.610 6.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 42.180 6.870 42.500 ;
      LAYER met4 ;
        RECT 6.550 42.180 6.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 41.750 6.870 42.070 ;
      LAYER met4 ;
        RECT 6.550 41.750 6.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 41.320 6.870 41.640 ;
      LAYER met4 ;
        RECT 6.550 41.320 6.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 40.890 6.870 41.210 ;
      LAYER met4 ;
        RECT 6.550 40.890 6.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 40.460 6.870 40.780 ;
      LAYER met4 ;
        RECT 6.550 40.460 6.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 40.030 6.870 40.350 ;
      LAYER met4 ;
        RECT 6.550 40.030 6.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.550 39.600 6.870 39.920 ;
      LAYER met4 ;
        RECT 6.550 39.600 6.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 43.900 6.470 44.220 ;
      LAYER met4 ;
        RECT 6.150 43.900 6.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 43.470 6.470 43.790 ;
      LAYER met4 ;
        RECT 6.150 43.470 6.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 43.040 6.470 43.360 ;
      LAYER met4 ;
        RECT 6.150 43.040 6.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 42.610 6.470 42.930 ;
      LAYER met4 ;
        RECT 6.150 42.610 6.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 42.180 6.470 42.500 ;
      LAYER met4 ;
        RECT 6.150 42.180 6.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 41.750 6.470 42.070 ;
      LAYER met4 ;
        RECT 6.150 41.750 6.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 41.320 6.470 41.640 ;
      LAYER met4 ;
        RECT 6.150 41.320 6.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 40.890 6.470 41.210 ;
      LAYER met4 ;
        RECT 6.150 40.890 6.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 40.460 6.470 40.780 ;
      LAYER met4 ;
        RECT 6.150 40.460 6.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 40.030 6.470 40.350 ;
      LAYER met4 ;
        RECT 6.150 40.030 6.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.150 39.600 6.470 39.920 ;
      LAYER met4 ;
        RECT 6.150 39.600 6.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 43.900 6.070 44.220 ;
      LAYER met4 ;
        RECT 5.750 43.900 6.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 43.470 6.070 43.790 ;
      LAYER met4 ;
        RECT 5.750 43.470 6.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 43.040 6.070 43.360 ;
      LAYER met4 ;
        RECT 5.750 43.040 6.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 42.610 6.070 42.930 ;
      LAYER met4 ;
        RECT 5.750 42.610 6.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 42.180 6.070 42.500 ;
      LAYER met4 ;
        RECT 5.750 42.180 6.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 41.750 6.070 42.070 ;
      LAYER met4 ;
        RECT 5.750 41.750 6.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 41.320 6.070 41.640 ;
      LAYER met4 ;
        RECT 5.750 41.320 6.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 40.890 6.070 41.210 ;
      LAYER met4 ;
        RECT 5.750 40.890 6.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 40.460 6.070 40.780 ;
      LAYER met4 ;
        RECT 5.750 40.460 6.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 40.030 6.070 40.350 ;
      LAYER met4 ;
        RECT 5.750 40.030 6.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.750 39.600 6.070 39.920 ;
      LAYER met4 ;
        RECT 5.750 39.600 6.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 43.900 5.670 44.220 ;
      LAYER met4 ;
        RECT 5.350 43.900 5.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 43.470 5.670 43.790 ;
      LAYER met4 ;
        RECT 5.350 43.470 5.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 43.040 5.670 43.360 ;
      LAYER met4 ;
        RECT 5.350 43.040 5.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 42.610 5.670 42.930 ;
      LAYER met4 ;
        RECT 5.350 42.610 5.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 42.180 5.670 42.500 ;
      LAYER met4 ;
        RECT 5.350 42.180 5.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 41.750 5.670 42.070 ;
      LAYER met4 ;
        RECT 5.350 41.750 5.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 41.320 5.670 41.640 ;
      LAYER met4 ;
        RECT 5.350 41.320 5.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 40.890 5.670 41.210 ;
      LAYER met4 ;
        RECT 5.350 40.890 5.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 40.460 5.670 40.780 ;
      LAYER met4 ;
        RECT 5.350 40.460 5.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 40.030 5.670 40.350 ;
      LAYER met4 ;
        RECT 5.350 40.030 5.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.350 39.600 5.670 39.920 ;
      LAYER met4 ;
        RECT 5.350 39.600 5.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 43.900 5.270 44.220 ;
      LAYER met4 ;
        RECT 4.950 43.900 5.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 43.470 5.270 43.790 ;
      LAYER met4 ;
        RECT 4.950 43.470 5.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 43.040 5.270 43.360 ;
      LAYER met4 ;
        RECT 4.950 43.040 5.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 42.610 5.270 42.930 ;
      LAYER met4 ;
        RECT 4.950 42.610 5.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 42.180 5.270 42.500 ;
      LAYER met4 ;
        RECT 4.950 42.180 5.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 41.750 5.270 42.070 ;
      LAYER met4 ;
        RECT 4.950 41.750 5.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 41.320 5.270 41.640 ;
      LAYER met4 ;
        RECT 4.950 41.320 5.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 40.890 5.270 41.210 ;
      LAYER met4 ;
        RECT 4.950 40.890 5.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 40.460 5.270 40.780 ;
      LAYER met4 ;
        RECT 4.950 40.460 5.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 40.030 5.270 40.350 ;
      LAYER met4 ;
        RECT 4.950 40.030 5.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.950 39.600 5.270 39.920 ;
      LAYER met4 ;
        RECT 4.950 39.600 5.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 43.900 4.870 44.220 ;
      LAYER met4 ;
        RECT 4.550 43.900 4.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 43.470 4.870 43.790 ;
      LAYER met4 ;
        RECT 4.550 43.470 4.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 43.040 4.870 43.360 ;
      LAYER met4 ;
        RECT 4.550 43.040 4.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 42.610 4.870 42.930 ;
      LAYER met4 ;
        RECT 4.550 42.610 4.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 42.180 4.870 42.500 ;
      LAYER met4 ;
        RECT 4.550 42.180 4.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 41.750 4.870 42.070 ;
      LAYER met4 ;
        RECT 4.550 41.750 4.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 41.320 4.870 41.640 ;
      LAYER met4 ;
        RECT 4.550 41.320 4.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 40.890 4.870 41.210 ;
      LAYER met4 ;
        RECT 4.550 40.890 4.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 40.460 4.870 40.780 ;
      LAYER met4 ;
        RECT 4.550 40.460 4.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 40.030 4.870 40.350 ;
      LAYER met4 ;
        RECT 4.550 40.030 4.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 39.600 4.870 39.920 ;
      LAYER met4 ;
        RECT 4.550 39.600 4.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 43.900 4.470 44.220 ;
      LAYER met4 ;
        RECT 4.150 43.900 4.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 43.470 4.470 43.790 ;
      LAYER met4 ;
        RECT 4.150 43.470 4.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 43.040 4.470 43.360 ;
      LAYER met4 ;
        RECT 4.150 43.040 4.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 42.610 4.470 42.930 ;
      LAYER met4 ;
        RECT 4.150 42.610 4.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 42.180 4.470 42.500 ;
      LAYER met4 ;
        RECT 4.150 42.180 4.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 41.750 4.470 42.070 ;
      LAYER met4 ;
        RECT 4.150 41.750 4.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 41.320 4.470 41.640 ;
      LAYER met4 ;
        RECT 4.150 41.320 4.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 40.890 4.470 41.210 ;
      LAYER met4 ;
        RECT 4.150 40.890 4.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 40.460 4.470 40.780 ;
      LAYER met4 ;
        RECT 4.150 40.460 4.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 40.030 4.470 40.350 ;
      LAYER met4 ;
        RECT 4.150 40.030 4.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.150 39.600 4.470 39.920 ;
      LAYER met4 ;
        RECT 4.150 39.600 4.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 43.900 4.070 44.220 ;
      LAYER met4 ;
        RECT 3.750 43.900 4.070 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 43.470 4.070 43.790 ;
      LAYER met4 ;
        RECT 3.750 43.470 4.070 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 43.040 4.070 43.360 ;
      LAYER met4 ;
        RECT 3.750 43.040 4.070 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 42.610 4.070 42.930 ;
      LAYER met4 ;
        RECT 3.750 42.610 4.070 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 42.180 4.070 42.500 ;
      LAYER met4 ;
        RECT 3.750 42.180 4.070 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 41.750 4.070 42.070 ;
      LAYER met4 ;
        RECT 3.750 41.750 4.070 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 41.320 4.070 41.640 ;
      LAYER met4 ;
        RECT 3.750 41.320 4.070 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 40.890 4.070 41.210 ;
      LAYER met4 ;
        RECT 3.750 40.890 4.070 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 40.460 4.070 40.780 ;
      LAYER met4 ;
        RECT 3.750 40.460 4.070 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 40.030 4.070 40.350 ;
      LAYER met4 ;
        RECT 3.750 40.030 4.070 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.750 39.600 4.070 39.920 ;
      LAYER met4 ;
        RECT 3.750 39.600 4.070 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 43.900 3.670 44.220 ;
      LAYER met4 ;
        RECT 3.350 43.900 3.670 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 43.470 3.670 43.790 ;
      LAYER met4 ;
        RECT 3.350 43.470 3.670 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 43.040 3.670 43.360 ;
      LAYER met4 ;
        RECT 3.350 43.040 3.670 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 42.610 3.670 42.930 ;
      LAYER met4 ;
        RECT 3.350 42.610 3.670 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 42.180 3.670 42.500 ;
      LAYER met4 ;
        RECT 3.350 42.180 3.670 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 41.750 3.670 42.070 ;
      LAYER met4 ;
        RECT 3.350 41.750 3.670 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 41.320 3.670 41.640 ;
      LAYER met4 ;
        RECT 3.350 41.320 3.670 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 40.890 3.670 41.210 ;
      LAYER met4 ;
        RECT 3.350 40.890 3.670 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 40.460 3.670 40.780 ;
      LAYER met4 ;
        RECT 3.350 40.460 3.670 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 40.030 3.670 40.350 ;
      LAYER met4 ;
        RECT 3.350 40.030 3.670 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.350 39.600 3.670 39.920 ;
      LAYER met4 ;
        RECT 3.350 39.600 3.670 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 43.900 3.270 44.220 ;
      LAYER met4 ;
        RECT 2.950 43.900 3.270 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 43.470 3.270 43.790 ;
      LAYER met4 ;
        RECT 2.950 43.470 3.270 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 43.040 3.270 43.360 ;
      LAYER met4 ;
        RECT 2.950 43.040 3.270 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 42.610 3.270 42.930 ;
      LAYER met4 ;
        RECT 2.950 42.610 3.270 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 42.180 3.270 42.500 ;
      LAYER met4 ;
        RECT 2.950 42.180 3.270 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 41.750 3.270 42.070 ;
      LAYER met4 ;
        RECT 2.950 41.750 3.270 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 41.320 3.270 41.640 ;
      LAYER met4 ;
        RECT 2.950 41.320 3.270 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 40.890 3.270 41.210 ;
      LAYER met4 ;
        RECT 2.950 40.890 3.270 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 40.460 3.270 40.780 ;
      LAYER met4 ;
        RECT 2.950 40.460 3.270 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 40.030 3.270 40.350 ;
      LAYER met4 ;
        RECT 2.950 40.030 3.270 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.950 39.600 3.270 39.920 ;
      LAYER met4 ;
        RECT 2.950 39.600 3.270 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 43.900 2.870 44.220 ;
      LAYER met4 ;
        RECT 2.550 43.900 2.870 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 43.470 2.870 43.790 ;
      LAYER met4 ;
        RECT 2.550 43.470 2.870 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 43.040 2.870 43.360 ;
      LAYER met4 ;
        RECT 2.550 43.040 2.870 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 42.610 2.870 42.930 ;
      LAYER met4 ;
        RECT 2.550 42.610 2.870 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 42.180 2.870 42.500 ;
      LAYER met4 ;
        RECT 2.550 42.180 2.870 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 41.750 2.870 42.070 ;
      LAYER met4 ;
        RECT 2.550 41.750 2.870 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 41.320 2.870 41.640 ;
      LAYER met4 ;
        RECT 2.550 41.320 2.870 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 40.890 2.870 41.210 ;
      LAYER met4 ;
        RECT 2.550 40.890 2.870 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 40.460 2.870 40.780 ;
      LAYER met4 ;
        RECT 2.550 40.460 2.870 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 40.030 2.870 40.350 ;
      LAYER met4 ;
        RECT 2.550 40.030 2.870 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.550 39.600 2.870 39.920 ;
      LAYER met4 ;
        RECT 2.550 39.600 2.870 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 43.900 2.470 44.220 ;
      LAYER met4 ;
        RECT 2.150 43.900 2.470 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 43.470 2.470 43.790 ;
      LAYER met4 ;
        RECT 2.150 43.470 2.470 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 43.040 2.470 43.360 ;
      LAYER met4 ;
        RECT 2.150 43.040 2.470 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 42.610 2.470 42.930 ;
      LAYER met4 ;
        RECT 2.150 42.610 2.470 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 42.180 2.470 42.500 ;
      LAYER met4 ;
        RECT 2.150 42.180 2.470 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 41.750 2.470 42.070 ;
      LAYER met4 ;
        RECT 2.150 41.750 2.470 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 41.320 2.470 41.640 ;
      LAYER met4 ;
        RECT 2.150 41.320 2.470 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 40.890 2.470 41.210 ;
      LAYER met4 ;
        RECT 2.150 40.890 2.470 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 40.460 2.470 40.780 ;
      LAYER met4 ;
        RECT 2.150 40.460 2.470 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 40.030 2.470 40.350 ;
      LAYER met4 ;
        RECT 2.150 40.030 2.470 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.150 39.600 2.470 39.920 ;
      LAYER met4 ;
        RECT 2.150 39.600 2.470 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 43.900 2.065 44.220 ;
      LAYER met4 ;
        RECT 1.745 43.900 2.065 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 43.470 2.065 43.790 ;
      LAYER met4 ;
        RECT 1.745 43.470 2.065 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 43.040 2.065 43.360 ;
      LAYER met4 ;
        RECT 1.745 43.040 2.065 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 42.610 2.065 42.930 ;
      LAYER met4 ;
        RECT 1.745 42.610 2.065 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 42.180 2.065 42.500 ;
      LAYER met4 ;
        RECT 1.745 42.180 2.065 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 41.750 2.065 42.070 ;
      LAYER met4 ;
        RECT 1.745 41.750 2.065 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 41.320 2.065 41.640 ;
      LAYER met4 ;
        RECT 1.745 41.320 2.065 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 40.890 2.065 41.210 ;
      LAYER met4 ;
        RECT 1.745 40.890 2.065 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 40.460 2.065 40.780 ;
      LAYER met4 ;
        RECT 1.745 40.460 2.065 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 40.030 2.065 40.350 ;
      LAYER met4 ;
        RECT 1.745 40.030 2.065 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.745 39.600 2.065 39.920 ;
      LAYER met4 ;
        RECT 1.745 39.600 2.065 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 43.900 1.660 44.220 ;
      LAYER met4 ;
        RECT 1.340 43.900 1.660 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 43.470 1.660 43.790 ;
      LAYER met4 ;
        RECT 1.340 43.470 1.660 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 43.040 1.660 43.360 ;
      LAYER met4 ;
        RECT 1.340 43.040 1.660 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 42.610 1.660 42.930 ;
      LAYER met4 ;
        RECT 1.340 42.610 1.660 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 42.180 1.660 42.500 ;
      LAYER met4 ;
        RECT 1.340 42.180 1.660 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 41.750 1.660 42.070 ;
      LAYER met4 ;
        RECT 1.340 41.750 1.660 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 41.320 1.660 41.640 ;
      LAYER met4 ;
        RECT 1.340 41.320 1.660 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 40.890 1.660 41.210 ;
      LAYER met4 ;
        RECT 1.340 40.890 1.660 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 40.460 1.660 40.780 ;
      LAYER met4 ;
        RECT 1.340 40.460 1.660 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 40.030 1.660 40.350 ;
      LAYER met4 ;
        RECT 1.340 40.030 1.660 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.340 39.600 1.660 39.920 ;
      LAYER met4 ;
        RECT 1.340 39.600 1.660 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 43.900 1.255 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 43.470 1.255 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 43.040 1.255 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 42.610 1.255 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 42.180 1.255 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 41.750 1.255 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 41.320 1.255 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 40.890 1.255 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 40.460 1.255 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 40.030 1.255 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 39.600 1.255 39.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 43.900 0.850 44.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 43.470 0.850 43.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 43.040 0.850 43.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 42.610 0.850 42.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 42.180 0.850 42.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 41.750 0.850 42.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 41.320 0.850 41.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 40.890 0.850 41.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 40.460 0.850 40.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 40.030 0.850 40.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 39.600 0.850 39.920 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
  END VSSIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
  END VSWITCH
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
  END VSSIO_Q
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
  END VCCHIB
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  OBS
      LAYER met3 ;
        RECT 0.500 39.590 24.500 44.230 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 94.585 75.000 172.185 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__overlay_vssd_lvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vssio_hvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vssio_hvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
  END VSSA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
  END VDDIO_Q
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.495 25.840 24.395 30.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 25.840 74.290 30.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.595 196.230 14.255 196.970 ;
    END
    PORT
      LAYER met4 ;
        RECT 13.630 197.170 61.325 199.930 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.680 196.230 61.340 196.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 30.210 74.200 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 29.780 74.200 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 29.350 74.200 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 28.920 74.200 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 28.490 74.200 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 28.060 74.200 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 27.630 74.200 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 27.200 74.200 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 26.770 74.200 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 26.340 74.200 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 25.910 74.200 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 199.595 74.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 199.190 74.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 198.785 74.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 198.380 74.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 197.975 74.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 197.570 74.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 197.165 74.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 196.760 74.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 196.355 74.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 195.950 74.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 195.545 74.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.930 195.140 74.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 175.935 74.250 195.055 ;
      LAYER met4 ;
        RECT 61.530 175.935 73.730 195.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 30.210 73.795 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 29.780 73.795 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 29.350 73.795 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 28.920 73.795 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 28.490 73.795 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 28.060 73.795 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 27.630 73.795 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 27.200 73.795 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 26.770 73.795 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 26.340 73.795 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 25.910 73.795 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 199.595 73.850 199.915 ;
      LAYER met4 ;
        RECT 73.530 199.595 73.730 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 199.190 73.850 199.510 ;
      LAYER met4 ;
        RECT 73.530 199.190 73.730 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 198.785 73.850 199.105 ;
      LAYER met4 ;
        RECT 73.530 198.785 73.730 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 198.380 73.850 198.700 ;
      LAYER met4 ;
        RECT 73.530 198.380 73.730 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 197.975 73.850 198.295 ;
      LAYER met4 ;
        RECT 73.530 197.975 73.730 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 197.570 73.850 197.890 ;
      LAYER met4 ;
        RECT 73.530 197.570 73.730 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 197.165 73.850 197.485 ;
      LAYER met4 ;
        RECT 73.530 197.165 73.730 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 196.760 73.850 197.080 ;
      LAYER met4 ;
        RECT 73.530 196.760 73.730 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 196.355 73.850 196.675 ;
      LAYER met4 ;
        RECT 73.530 196.355 73.730 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 195.950 73.850 196.270 ;
      LAYER met4 ;
        RECT 73.530 195.950 73.730 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 195.545 73.850 195.865 ;
      LAYER met4 ;
        RECT 73.530 195.545 73.730 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.530 195.140 73.850 195.460 ;
      LAYER met4 ;
        RECT 73.530 195.140 73.730 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 199.595 73.450 199.915 ;
      LAYER met4 ;
        RECT 73.130 199.595 73.450 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 199.190 73.450 199.510 ;
      LAYER met4 ;
        RECT 73.130 199.190 73.450 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 198.785 73.450 199.105 ;
      LAYER met4 ;
        RECT 73.130 198.785 73.450 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 198.380 73.450 198.700 ;
      LAYER met4 ;
        RECT 73.130 198.380 73.450 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 197.975 73.450 198.295 ;
      LAYER met4 ;
        RECT 73.130 197.975 73.450 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 197.570 73.450 197.890 ;
      LAYER met4 ;
        RECT 73.130 197.570 73.450 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 197.165 73.450 197.485 ;
      LAYER met4 ;
        RECT 73.130 197.165 73.450 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 196.760 73.450 197.080 ;
      LAYER met4 ;
        RECT 73.130 196.760 73.450 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 196.355 73.450 196.675 ;
      LAYER met4 ;
        RECT 73.130 196.355 73.450 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 195.950 73.450 196.270 ;
      LAYER met4 ;
        RECT 73.130 195.950 73.450 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 195.545 73.450 195.865 ;
      LAYER met4 ;
        RECT 73.130 195.545 73.450 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 195.140 73.450 195.460 ;
      LAYER met4 ;
        RECT 73.130 195.140 73.450 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 30.210 73.390 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 29.780 73.390 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 29.350 73.390 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 28.920 73.390 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 28.490 73.390 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 28.060 73.390 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 27.630 73.390 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 27.200 73.390 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 26.770 73.390 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 26.340 73.390 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 25.910 73.390 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 199.595 73.050 199.915 ;
      LAYER met4 ;
        RECT 72.730 199.595 73.050 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 199.190 73.050 199.510 ;
      LAYER met4 ;
        RECT 72.730 199.190 73.050 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 198.785 73.050 199.105 ;
      LAYER met4 ;
        RECT 72.730 198.785 73.050 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 198.380 73.050 198.700 ;
      LAYER met4 ;
        RECT 72.730 198.380 73.050 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 197.975 73.050 198.295 ;
      LAYER met4 ;
        RECT 72.730 197.975 73.050 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 197.570 73.050 197.890 ;
      LAYER met4 ;
        RECT 72.730 197.570 73.050 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 197.165 73.050 197.485 ;
      LAYER met4 ;
        RECT 72.730 197.165 73.050 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 196.760 73.050 197.080 ;
      LAYER met4 ;
        RECT 72.730 196.760 73.050 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 196.355 73.050 196.675 ;
      LAYER met4 ;
        RECT 72.730 196.355 73.050 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 195.950 73.050 196.270 ;
      LAYER met4 ;
        RECT 72.730 195.950 73.050 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 195.545 73.050 195.865 ;
      LAYER met4 ;
        RECT 72.730 195.545 73.050 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.730 195.140 73.050 195.460 ;
      LAYER met4 ;
        RECT 72.730 195.140 73.050 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 30.210 72.985 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 29.780 72.985 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 29.350 72.985 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 28.920 72.985 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 28.490 72.985 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 28.060 72.985 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 27.630 72.985 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 27.200 72.985 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 26.770 72.985 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 26.340 72.985 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 25.910 72.985 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 199.595 72.650 199.915 ;
      LAYER met4 ;
        RECT 72.330 199.595 72.650 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 199.190 72.650 199.510 ;
      LAYER met4 ;
        RECT 72.330 199.190 72.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 198.785 72.650 199.105 ;
      LAYER met4 ;
        RECT 72.330 198.785 72.650 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 198.380 72.650 198.700 ;
      LAYER met4 ;
        RECT 72.330 198.380 72.650 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 197.975 72.650 198.295 ;
      LAYER met4 ;
        RECT 72.330 197.975 72.650 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 197.570 72.650 197.890 ;
      LAYER met4 ;
        RECT 72.330 197.570 72.650 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 197.165 72.650 197.485 ;
      LAYER met4 ;
        RECT 72.330 197.165 72.650 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 196.760 72.650 197.080 ;
      LAYER met4 ;
        RECT 72.330 196.760 72.650 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 196.355 72.650 196.675 ;
      LAYER met4 ;
        RECT 72.330 196.355 72.650 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 195.950 72.650 196.270 ;
      LAYER met4 ;
        RECT 72.330 195.950 72.650 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 195.545 72.650 195.865 ;
      LAYER met4 ;
        RECT 72.330 195.545 72.650 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.330 195.140 72.650 195.460 ;
      LAYER met4 ;
        RECT 72.330 195.140 72.650 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 30.210 72.580 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 29.780 72.580 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 29.350 72.580 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 28.920 72.580 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 28.490 72.580 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 28.060 72.580 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 27.630 72.580 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 27.200 72.580 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 26.770 72.580 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 26.340 72.580 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 25.910 72.580 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 199.595 72.250 199.915 ;
      LAYER met4 ;
        RECT 71.930 199.595 72.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 199.190 72.250 199.510 ;
      LAYER met4 ;
        RECT 71.930 199.190 72.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 198.785 72.250 199.105 ;
      LAYER met4 ;
        RECT 71.930 198.785 72.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 198.380 72.250 198.700 ;
      LAYER met4 ;
        RECT 71.930 198.380 72.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 197.975 72.250 198.295 ;
      LAYER met4 ;
        RECT 71.930 197.975 72.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 197.570 72.250 197.890 ;
      LAYER met4 ;
        RECT 71.930 197.570 72.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 197.165 72.250 197.485 ;
      LAYER met4 ;
        RECT 71.930 197.165 72.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 196.760 72.250 197.080 ;
      LAYER met4 ;
        RECT 71.930 196.760 72.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 196.355 72.250 196.675 ;
      LAYER met4 ;
        RECT 71.930 196.355 72.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 195.950 72.250 196.270 ;
      LAYER met4 ;
        RECT 71.930 195.950 72.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 195.545 72.250 195.865 ;
      LAYER met4 ;
        RECT 71.930 195.545 72.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.930 195.140 72.250 195.460 ;
      LAYER met4 ;
        RECT 71.930 195.140 72.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 30.210 72.175 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 29.780 72.175 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 29.350 72.175 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 28.920 72.175 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 28.490 72.175 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 28.060 72.175 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 27.630 72.175 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 27.200 72.175 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 26.770 72.175 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 26.340 72.175 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 25.910 72.175 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 199.595 71.850 199.915 ;
      LAYER met4 ;
        RECT 71.530 199.595 71.850 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 199.190 71.850 199.510 ;
      LAYER met4 ;
        RECT 71.530 199.190 71.850 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 198.785 71.850 199.105 ;
      LAYER met4 ;
        RECT 71.530 198.785 71.850 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 198.380 71.850 198.700 ;
      LAYER met4 ;
        RECT 71.530 198.380 71.850 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 197.975 71.850 198.295 ;
      LAYER met4 ;
        RECT 71.530 197.975 71.850 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 197.570 71.850 197.890 ;
      LAYER met4 ;
        RECT 71.530 197.570 71.850 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 197.165 71.850 197.485 ;
      LAYER met4 ;
        RECT 71.530 197.165 71.850 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 196.760 71.850 197.080 ;
      LAYER met4 ;
        RECT 71.530 196.760 71.850 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 196.355 71.850 196.675 ;
      LAYER met4 ;
        RECT 71.530 196.355 71.850 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 195.950 71.850 196.270 ;
      LAYER met4 ;
        RECT 71.530 195.950 71.850 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 195.545 71.850 195.865 ;
      LAYER met4 ;
        RECT 71.530 195.545 71.850 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 195.140 71.850 195.460 ;
      LAYER met4 ;
        RECT 71.530 195.140 71.850 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 30.210 71.770 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 29.780 71.770 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 29.350 71.770 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 28.920 71.770 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 28.490 71.770 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 28.060 71.770 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 27.630 71.770 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 27.200 71.770 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 26.770 71.770 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 26.340 71.770 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 25.910 71.770 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 199.595 71.450 199.915 ;
      LAYER met4 ;
        RECT 71.130 199.595 71.450 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 199.190 71.450 199.510 ;
      LAYER met4 ;
        RECT 71.130 199.190 71.450 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 198.785 71.450 199.105 ;
      LAYER met4 ;
        RECT 71.130 198.785 71.450 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 198.380 71.450 198.700 ;
      LAYER met4 ;
        RECT 71.130 198.380 71.450 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 197.975 71.450 198.295 ;
      LAYER met4 ;
        RECT 71.130 197.975 71.450 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 197.570 71.450 197.890 ;
      LAYER met4 ;
        RECT 71.130 197.570 71.450 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 197.165 71.450 197.485 ;
      LAYER met4 ;
        RECT 71.130 197.165 71.450 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 196.760 71.450 197.080 ;
      LAYER met4 ;
        RECT 71.130 196.760 71.450 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 196.355 71.450 196.675 ;
      LAYER met4 ;
        RECT 71.130 196.355 71.450 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 195.950 71.450 196.270 ;
      LAYER met4 ;
        RECT 71.130 195.950 71.450 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 195.545 71.450 195.865 ;
      LAYER met4 ;
        RECT 71.130 195.545 71.450 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.130 195.140 71.450 195.460 ;
      LAYER met4 ;
        RECT 71.130 195.140 71.450 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 30.210 71.365 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 29.780 71.365 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 29.350 71.365 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 28.920 71.365 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 28.490 71.365 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 28.060 71.365 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 27.630 71.365 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 27.200 71.365 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 26.770 71.365 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 26.340 71.365 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 25.910 71.365 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 199.595 71.050 199.915 ;
      LAYER met4 ;
        RECT 70.730 199.595 71.050 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 199.190 71.050 199.510 ;
      LAYER met4 ;
        RECT 70.730 199.190 71.050 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 198.785 71.050 199.105 ;
      LAYER met4 ;
        RECT 70.730 198.785 71.050 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 198.380 71.050 198.700 ;
      LAYER met4 ;
        RECT 70.730 198.380 71.050 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 197.975 71.050 198.295 ;
      LAYER met4 ;
        RECT 70.730 197.975 71.050 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 197.570 71.050 197.890 ;
      LAYER met4 ;
        RECT 70.730 197.570 71.050 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 197.165 71.050 197.485 ;
      LAYER met4 ;
        RECT 70.730 197.165 71.050 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 196.760 71.050 197.080 ;
      LAYER met4 ;
        RECT 70.730 196.760 71.050 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 196.355 71.050 196.675 ;
      LAYER met4 ;
        RECT 70.730 196.355 71.050 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 195.950 71.050 196.270 ;
      LAYER met4 ;
        RECT 70.730 195.950 71.050 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 195.545 71.050 195.865 ;
      LAYER met4 ;
        RECT 70.730 195.545 71.050 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.730 195.140 71.050 195.460 ;
      LAYER met4 ;
        RECT 70.730 195.140 71.050 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 30.210 70.960 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 29.780 70.960 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 29.350 70.960 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 28.920 70.960 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 28.490 70.960 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 28.060 70.960 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 27.630 70.960 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 27.200 70.960 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 26.770 70.960 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 26.340 70.960 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 25.910 70.960 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 199.595 70.650 199.915 ;
      LAYER met4 ;
        RECT 70.330 199.595 70.650 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 199.190 70.650 199.510 ;
      LAYER met4 ;
        RECT 70.330 199.190 70.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 198.785 70.650 199.105 ;
      LAYER met4 ;
        RECT 70.330 198.785 70.650 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 198.380 70.650 198.700 ;
      LAYER met4 ;
        RECT 70.330 198.380 70.650 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 197.975 70.650 198.295 ;
      LAYER met4 ;
        RECT 70.330 197.975 70.650 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 197.570 70.650 197.890 ;
      LAYER met4 ;
        RECT 70.330 197.570 70.650 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 197.165 70.650 197.485 ;
      LAYER met4 ;
        RECT 70.330 197.165 70.650 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 196.760 70.650 197.080 ;
      LAYER met4 ;
        RECT 70.330 196.760 70.650 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 196.355 70.650 196.675 ;
      LAYER met4 ;
        RECT 70.330 196.355 70.650 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 195.950 70.650 196.270 ;
      LAYER met4 ;
        RECT 70.330 195.950 70.650 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 195.545 70.650 195.865 ;
      LAYER met4 ;
        RECT 70.330 195.545 70.650 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.330 195.140 70.650 195.460 ;
      LAYER met4 ;
        RECT 70.330 195.140 70.650 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 30.210 70.555 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 29.780 70.555 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 29.350 70.555 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 28.920 70.555 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 28.490 70.555 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 28.060 70.555 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 27.630 70.555 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 27.200 70.555 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 26.770 70.555 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 26.340 70.555 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 25.910 70.555 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 199.595 70.250 199.915 ;
      LAYER met4 ;
        RECT 69.930 199.595 70.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 199.190 70.250 199.510 ;
      LAYER met4 ;
        RECT 69.930 199.190 70.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 198.785 70.250 199.105 ;
      LAYER met4 ;
        RECT 69.930 198.785 70.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 198.380 70.250 198.700 ;
      LAYER met4 ;
        RECT 69.930 198.380 70.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 197.975 70.250 198.295 ;
      LAYER met4 ;
        RECT 69.930 197.975 70.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 197.570 70.250 197.890 ;
      LAYER met4 ;
        RECT 69.930 197.570 70.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 197.165 70.250 197.485 ;
      LAYER met4 ;
        RECT 69.930 197.165 70.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 196.760 70.250 197.080 ;
      LAYER met4 ;
        RECT 69.930 196.760 70.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 196.355 70.250 196.675 ;
      LAYER met4 ;
        RECT 69.930 196.355 70.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 195.950 70.250 196.270 ;
      LAYER met4 ;
        RECT 69.930 195.950 70.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 195.545 70.250 195.865 ;
      LAYER met4 ;
        RECT 69.930 195.545 70.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 195.140 70.250 195.460 ;
      LAYER met4 ;
        RECT 69.930 195.140 70.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 30.210 70.150 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 29.780 70.150 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 29.350 70.150 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 28.920 70.150 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 28.490 70.150 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 28.060 70.150 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 27.630 70.150 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 27.200 70.150 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 26.770 70.150 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 26.340 70.150 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 25.910 70.150 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 199.595 69.850 199.915 ;
      LAYER met4 ;
        RECT 69.530 199.595 69.850 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 199.190 69.850 199.510 ;
      LAYER met4 ;
        RECT 69.530 199.190 69.850 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 198.785 69.850 199.105 ;
      LAYER met4 ;
        RECT 69.530 198.785 69.850 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 198.380 69.850 198.700 ;
      LAYER met4 ;
        RECT 69.530 198.380 69.850 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 197.975 69.850 198.295 ;
      LAYER met4 ;
        RECT 69.530 197.975 69.850 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 197.570 69.850 197.890 ;
      LAYER met4 ;
        RECT 69.530 197.570 69.850 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 197.165 69.850 197.485 ;
      LAYER met4 ;
        RECT 69.530 197.165 69.850 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 196.760 69.850 197.080 ;
      LAYER met4 ;
        RECT 69.530 196.760 69.850 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 196.355 69.850 196.675 ;
      LAYER met4 ;
        RECT 69.530 196.355 69.850 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 195.950 69.850 196.270 ;
      LAYER met4 ;
        RECT 69.530 195.950 69.850 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 195.545 69.850 195.865 ;
      LAYER met4 ;
        RECT 69.530 195.545 69.850 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.530 195.140 69.850 195.460 ;
      LAYER met4 ;
        RECT 69.530 195.140 69.850 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 30.210 69.745 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 29.780 69.745 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 29.350 69.745 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 28.920 69.745 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 28.490 69.745 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 28.060 69.745 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 27.630 69.745 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 27.200 69.745 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 26.770 69.745 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 26.340 69.745 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 25.910 69.745 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 199.595 69.450 199.915 ;
      LAYER met4 ;
        RECT 69.130 199.595 69.450 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 199.190 69.450 199.510 ;
      LAYER met4 ;
        RECT 69.130 199.190 69.450 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 198.785 69.450 199.105 ;
      LAYER met4 ;
        RECT 69.130 198.785 69.450 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 198.380 69.450 198.700 ;
      LAYER met4 ;
        RECT 69.130 198.380 69.450 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 197.975 69.450 198.295 ;
      LAYER met4 ;
        RECT 69.130 197.975 69.450 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 197.570 69.450 197.890 ;
      LAYER met4 ;
        RECT 69.130 197.570 69.450 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 197.165 69.450 197.485 ;
      LAYER met4 ;
        RECT 69.130 197.165 69.450 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 196.760 69.450 197.080 ;
      LAYER met4 ;
        RECT 69.130 196.760 69.450 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 196.355 69.450 196.675 ;
      LAYER met4 ;
        RECT 69.130 196.355 69.450 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 195.950 69.450 196.270 ;
      LAYER met4 ;
        RECT 69.130 195.950 69.450 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 195.545 69.450 195.865 ;
      LAYER met4 ;
        RECT 69.130 195.545 69.450 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.130 195.140 69.450 195.460 ;
      LAYER met4 ;
        RECT 69.130 195.140 69.450 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 30.210 69.340 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 29.780 69.340 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 29.350 69.340 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 28.920 69.340 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 28.490 69.340 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 28.060 69.340 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 27.630 69.340 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 27.200 69.340 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 26.770 69.340 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 26.340 69.340 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 25.910 69.340 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 199.595 69.050 199.915 ;
      LAYER met4 ;
        RECT 68.730 199.595 69.050 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 199.190 69.050 199.510 ;
      LAYER met4 ;
        RECT 68.730 199.190 69.050 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 198.785 69.050 199.105 ;
      LAYER met4 ;
        RECT 68.730 198.785 69.050 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 198.380 69.050 198.700 ;
      LAYER met4 ;
        RECT 68.730 198.380 69.050 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 197.975 69.050 198.295 ;
      LAYER met4 ;
        RECT 68.730 197.975 69.050 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 197.570 69.050 197.890 ;
      LAYER met4 ;
        RECT 68.730 197.570 69.050 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 197.165 69.050 197.485 ;
      LAYER met4 ;
        RECT 68.730 197.165 69.050 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 196.760 69.050 197.080 ;
      LAYER met4 ;
        RECT 68.730 196.760 69.050 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 196.355 69.050 196.675 ;
      LAYER met4 ;
        RECT 68.730 196.355 69.050 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 195.950 69.050 196.270 ;
      LAYER met4 ;
        RECT 68.730 195.950 69.050 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 195.545 69.050 195.865 ;
      LAYER met4 ;
        RECT 68.730 195.545 69.050 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.730 195.140 69.050 195.460 ;
      LAYER met4 ;
        RECT 68.730 195.140 69.050 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 30.210 68.935 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 29.780 68.935 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 29.350 68.935 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 28.920 68.935 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 28.490 68.935 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 28.060 68.935 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 27.630 68.935 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 27.200 68.935 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 26.770 68.935 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 26.340 68.935 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 25.910 68.935 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 199.595 68.650 199.915 ;
      LAYER met4 ;
        RECT 68.330 199.595 68.650 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 199.190 68.650 199.510 ;
      LAYER met4 ;
        RECT 68.330 199.190 68.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 198.785 68.650 199.105 ;
      LAYER met4 ;
        RECT 68.330 198.785 68.650 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 198.380 68.650 198.700 ;
      LAYER met4 ;
        RECT 68.330 198.380 68.650 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 197.975 68.650 198.295 ;
      LAYER met4 ;
        RECT 68.330 197.975 68.650 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 197.570 68.650 197.890 ;
      LAYER met4 ;
        RECT 68.330 197.570 68.650 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 197.165 68.650 197.485 ;
      LAYER met4 ;
        RECT 68.330 197.165 68.650 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 196.760 68.650 197.080 ;
      LAYER met4 ;
        RECT 68.330 196.760 68.650 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 196.355 68.650 196.675 ;
      LAYER met4 ;
        RECT 68.330 196.355 68.650 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 195.950 68.650 196.270 ;
      LAYER met4 ;
        RECT 68.330 195.950 68.650 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 195.545 68.650 195.865 ;
      LAYER met4 ;
        RECT 68.330 195.545 68.650 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 195.140 68.650 195.460 ;
      LAYER met4 ;
        RECT 68.330 195.140 68.650 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 30.210 68.530 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 29.780 68.530 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 29.350 68.530 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 28.920 68.530 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 28.490 68.530 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 28.060 68.530 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 27.630 68.530 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 27.200 68.530 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 26.770 68.530 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 26.340 68.530 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 25.910 68.530 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 199.595 68.250 199.915 ;
      LAYER met4 ;
        RECT 67.930 199.595 68.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 199.190 68.250 199.510 ;
      LAYER met4 ;
        RECT 67.930 199.190 68.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 198.785 68.250 199.105 ;
      LAYER met4 ;
        RECT 67.930 198.785 68.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 198.380 68.250 198.700 ;
      LAYER met4 ;
        RECT 67.930 198.380 68.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 197.975 68.250 198.295 ;
      LAYER met4 ;
        RECT 67.930 197.975 68.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 197.570 68.250 197.890 ;
      LAYER met4 ;
        RECT 67.930 197.570 68.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 197.165 68.250 197.485 ;
      LAYER met4 ;
        RECT 67.930 197.165 68.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 196.760 68.250 197.080 ;
      LAYER met4 ;
        RECT 67.930 196.760 68.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 196.355 68.250 196.675 ;
      LAYER met4 ;
        RECT 67.930 196.355 68.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 195.950 68.250 196.270 ;
      LAYER met4 ;
        RECT 67.930 195.950 68.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 195.545 68.250 195.865 ;
      LAYER met4 ;
        RECT 67.930 195.545 68.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.930 195.140 68.250 195.460 ;
      LAYER met4 ;
        RECT 67.930 195.140 68.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 30.210 68.125 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 29.780 68.125 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 29.350 68.125 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 28.920 68.125 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 28.490 68.125 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 28.060 68.125 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 27.630 68.125 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 27.200 68.125 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 26.770 68.125 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 26.340 68.125 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 25.910 68.125 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 199.595 67.850 199.915 ;
      LAYER met4 ;
        RECT 67.530 199.595 67.850 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 199.190 67.850 199.510 ;
      LAYER met4 ;
        RECT 67.530 199.190 67.850 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 198.785 67.850 199.105 ;
      LAYER met4 ;
        RECT 67.530 198.785 67.850 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 198.380 67.850 198.700 ;
      LAYER met4 ;
        RECT 67.530 198.380 67.850 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 197.975 67.850 198.295 ;
      LAYER met4 ;
        RECT 67.530 197.975 67.850 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 197.570 67.850 197.890 ;
      LAYER met4 ;
        RECT 67.530 197.570 67.850 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 197.165 67.850 197.485 ;
      LAYER met4 ;
        RECT 67.530 197.165 67.850 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 196.760 67.850 197.080 ;
      LAYER met4 ;
        RECT 67.530 196.760 67.850 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 196.355 67.850 196.675 ;
      LAYER met4 ;
        RECT 67.530 196.355 67.850 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 195.950 67.850 196.270 ;
      LAYER met4 ;
        RECT 67.530 195.950 67.850 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 195.545 67.850 195.865 ;
      LAYER met4 ;
        RECT 67.530 195.545 67.850 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.530 195.140 67.850 195.460 ;
      LAYER met4 ;
        RECT 67.530 195.140 67.850 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 30.210 67.720 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 29.780 67.720 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 29.350 67.720 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 28.920 67.720 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 28.490 67.720 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 28.060 67.720 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 27.630 67.720 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 27.200 67.720 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 26.770 67.720 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 26.340 67.720 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 25.910 67.720 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 199.595 67.450 199.915 ;
      LAYER met4 ;
        RECT 67.130 199.595 67.450 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 199.190 67.450 199.510 ;
      LAYER met4 ;
        RECT 67.130 199.190 67.450 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 198.785 67.450 199.105 ;
      LAYER met4 ;
        RECT 67.130 198.785 67.450 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 198.380 67.450 198.700 ;
      LAYER met4 ;
        RECT 67.130 198.380 67.450 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 197.975 67.450 198.295 ;
      LAYER met4 ;
        RECT 67.130 197.975 67.450 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 197.570 67.450 197.890 ;
      LAYER met4 ;
        RECT 67.130 197.570 67.450 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 197.165 67.450 197.485 ;
      LAYER met4 ;
        RECT 67.130 197.165 67.450 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 196.760 67.450 197.080 ;
      LAYER met4 ;
        RECT 67.130 196.760 67.450 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 196.355 67.450 196.675 ;
      LAYER met4 ;
        RECT 67.130 196.355 67.450 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 195.950 67.450 196.270 ;
      LAYER met4 ;
        RECT 67.130 195.950 67.450 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 195.545 67.450 195.865 ;
      LAYER met4 ;
        RECT 67.130 195.545 67.450 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.130 195.140 67.450 195.460 ;
      LAYER met4 ;
        RECT 67.130 195.140 67.450 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 30.210 67.315 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 29.780 67.315 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 29.350 67.315 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 28.920 67.315 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 28.490 67.315 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 28.060 67.315 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 27.630 67.315 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 27.200 67.315 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 26.770 67.315 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 26.340 67.315 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 25.910 67.315 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 199.595 67.050 199.915 ;
      LAYER met4 ;
        RECT 66.730 199.595 67.050 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 199.190 67.050 199.510 ;
      LAYER met4 ;
        RECT 66.730 199.190 67.050 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 198.785 67.050 199.105 ;
      LAYER met4 ;
        RECT 66.730 198.785 67.050 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 198.380 67.050 198.700 ;
      LAYER met4 ;
        RECT 66.730 198.380 67.050 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 197.975 67.050 198.295 ;
      LAYER met4 ;
        RECT 66.730 197.975 67.050 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 197.570 67.050 197.890 ;
      LAYER met4 ;
        RECT 66.730 197.570 67.050 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 197.165 67.050 197.485 ;
      LAYER met4 ;
        RECT 66.730 197.165 67.050 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 196.760 67.050 197.080 ;
      LAYER met4 ;
        RECT 66.730 196.760 67.050 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 196.355 67.050 196.675 ;
      LAYER met4 ;
        RECT 66.730 196.355 67.050 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 195.950 67.050 196.270 ;
      LAYER met4 ;
        RECT 66.730 195.950 67.050 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 195.545 67.050 195.865 ;
      LAYER met4 ;
        RECT 66.730 195.545 67.050 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.730 195.140 67.050 195.460 ;
      LAYER met4 ;
        RECT 66.730 195.140 67.050 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 30.210 66.910 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 29.780 66.910 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 29.350 66.910 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 28.920 66.910 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 28.490 66.910 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 28.060 66.910 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 27.630 66.910 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 27.200 66.910 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 26.770 66.910 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 26.340 66.910 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 25.910 66.910 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 199.595 66.650 199.915 ;
      LAYER met4 ;
        RECT 66.330 199.595 66.650 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 199.190 66.650 199.510 ;
      LAYER met4 ;
        RECT 66.330 199.190 66.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 198.785 66.650 199.105 ;
      LAYER met4 ;
        RECT 66.330 198.785 66.650 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 198.380 66.650 198.700 ;
      LAYER met4 ;
        RECT 66.330 198.380 66.650 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 197.975 66.650 198.295 ;
      LAYER met4 ;
        RECT 66.330 197.975 66.650 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 197.570 66.650 197.890 ;
      LAYER met4 ;
        RECT 66.330 197.570 66.650 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 197.165 66.650 197.485 ;
      LAYER met4 ;
        RECT 66.330 197.165 66.650 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 196.760 66.650 197.080 ;
      LAYER met4 ;
        RECT 66.330 196.760 66.650 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 196.355 66.650 196.675 ;
      LAYER met4 ;
        RECT 66.330 196.355 66.650 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 195.950 66.650 196.270 ;
      LAYER met4 ;
        RECT 66.330 195.950 66.650 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 195.545 66.650 195.865 ;
      LAYER met4 ;
        RECT 66.330 195.545 66.650 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.330 195.140 66.650 195.460 ;
      LAYER met4 ;
        RECT 66.330 195.140 66.650 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 30.210 66.505 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 29.780 66.505 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 29.350 66.505 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 28.920 66.505 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 28.490 66.505 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 28.060 66.505 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 27.630 66.505 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 27.200 66.505 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 26.770 66.505 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 26.340 66.505 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 25.910 66.505 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 199.595 66.250 199.915 ;
      LAYER met4 ;
        RECT 65.930 199.595 66.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 199.190 66.250 199.510 ;
      LAYER met4 ;
        RECT 65.930 199.190 66.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 198.785 66.250 199.105 ;
      LAYER met4 ;
        RECT 65.930 198.785 66.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 198.380 66.250 198.700 ;
      LAYER met4 ;
        RECT 65.930 198.380 66.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 197.975 66.250 198.295 ;
      LAYER met4 ;
        RECT 65.930 197.975 66.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 197.570 66.250 197.890 ;
      LAYER met4 ;
        RECT 65.930 197.570 66.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 197.165 66.250 197.485 ;
      LAYER met4 ;
        RECT 65.930 197.165 66.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 196.760 66.250 197.080 ;
      LAYER met4 ;
        RECT 65.930 196.760 66.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 196.355 66.250 196.675 ;
      LAYER met4 ;
        RECT 65.930 196.355 66.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 195.950 66.250 196.270 ;
      LAYER met4 ;
        RECT 65.930 195.950 66.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 195.545 66.250 195.865 ;
      LAYER met4 ;
        RECT 65.930 195.545 66.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.930 195.140 66.250 195.460 ;
      LAYER met4 ;
        RECT 65.930 195.140 66.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 30.210 66.100 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 29.780 66.100 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 29.350 66.100 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 28.920 66.100 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 28.490 66.100 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 28.060 66.100 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 27.630 66.100 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 27.200 66.100 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 26.770 66.100 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 26.340 66.100 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 25.910 66.100 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 199.595 65.850 199.915 ;
      LAYER met4 ;
        RECT 65.530 199.595 65.850 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 199.190 65.850 199.510 ;
      LAYER met4 ;
        RECT 65.530 199.190 65.850 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 198.785 65.850 199.105 ;
      LAYER met4 ;
        RECT 65.530 198.785 65.850 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 198.380 65.850 198.700 ;
      LAYER met4 ;
        RECT 65.530 198.380 65.850 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 197.975 65.850 198.295 ;
      LAYER met4 ;
        RECT 65.530 197.975 65.850 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 197.570 65.850 197.890 ;
      LAYER met4 ;
        RECT 65.530 197.570 65.850 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 197.165 65.850 197.485 ;
      LAYER met4 ;
        RECT 65.530 197.165 65.850 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 196.760 65.850 197.080 ;
      LAYER met4 ;
        RECT 65.530 196.760 65.850 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 196.355 65.850 196.675 ;
      LAYER met4 ;
        RECT 65.530 196.355 65.850 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 195.950 65.850 196.270 ;
      LAYER met4 ;
        RECT 65.530 195.950 65.850 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 195.545 65.850 195.865 ;
      LAYER met4 ;
        RECT 65.530 195.545 65.850 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.530 195.140 65.850 195.460 ;
      LAYER met4 ;
        RECT 65.530 195.140 65.850 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 30.210 65.695 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 29.780 65.695 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 29.350 65.695 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 28.920 65.695 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 28.490 65.695 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 28.060 65.695 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 27.630 65.695 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 27.200 65.695 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 26.770 65.695 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 26.340 65.695 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 25.910 65.695 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 199.595 65.450 199.915 ;
      LAYER met4 ;
        RECT 65.130 199.595 65.450 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 199.190 65.450 199.510 ;
      LAYER met4 ;
        RECT 65.130 199.190 65.450 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 198.785 65.450 199.105 ;
      LAYER met4 ;
        RECT 65.130 198.785 65.450 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 198.380 65.450 198.700 ;
      LAYER met4 ;
        RECT 65.130 198.380 65.450 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 197.975 65.450 198.295 ;
      LAYER met4 ;
        RECT 65.130 197.975 65.450 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 197.570 65.450 197.890 ;
      LAYER met4 ;
        RECT 65.130 197.570 65.450 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 197.165 65.450 197.485 ;
      LAYER met4 ;
        RECT 65.130 197.165 65.450 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 196.760 65.450 197.080 ;
      LAYER met4 ;
        RECT 65.130 196.760 65.450 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 196.355 65.450 196.675 ;
      LAYER met4 ;
        RECT 65.130 196.355 65.450 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 195.950 65.450 196.270 ;
      LAYER met4 ;
        RECT 65.130 195.950 65.450 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 195.545 65.450 195.865 ;
      LAYER met4 ;
        RECT 65.130 195.545 65.450 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.130 195.140 65.450 195.460 ;
      LAYER met4 ;
        RECT 65.130 195.140 65.450 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 30.210 65.290 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 29.780 65.290 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 29.350 65.290 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 28.920 65.290 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 28.490 65.290 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 28.060 65.290 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 27.630 65.290 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 27.200 65.290 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 26.770 65.290 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 26.340 65.290 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 25.910 65.290 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 199.595 65.050 199.915 ;
      LAYER met4 ;
        RECT 64.730 199.595 65.050 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 199.190 65.050 199.510 ;
      LAYER met4 ;
        RECT 64.730 199.190 65.050 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 198.785 65.050 199.105 ;
      LAYER met4 ;
        RECT 64.730 198.785 65.050 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 198.380 65.050 198.700 ;
      LAYER met4 ;
        RECT 64.730 198.380 65.050 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 197.975 65.050 198.295 ;
      LAYER met4 ;
        RECT 64.730 197.975 65.050 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 197.570 65.050 197.890 ;
      LAYER met4 ;
        RECT 64.730 197.570 65.050 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 197.165 65.050 197.485 ;
      LAYER met4 ;
        RECT 64.730 197.165 65.050 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 196.760 65.050 197.080 ;
      LAYER met4 ;
        RECT 64.730 196.760 65.050 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 196.355 65.050 196.675 ;
      LAYER met4 ;
        RECT 64.730 196.355 65.050 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 195.950 65.050 196.270 ;
      LAYER met4 ;
        RECT 64.730 195.950 65.050 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 195.545 65.050 195.865 ;
      LAYER met4 ;
        RECT 64.730 195.545 65.050 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.730 195.140 65.050 195.460 ;
      LAYER met4 ;
        RECT 64.730 195.140 65.050 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 30.210 64.885 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 29.780 64.885 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 29.350 64.885 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 28.920 64.885 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 28.490 64.885 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 28.060 64.885 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 27.630 64.885 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 27.200 64.885 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 26.770 64.885 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 26.340 64.885 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 25.910 64.885 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 199.595 64.650 199.915 ;
      LAYER met4 ;
        RECT 64.330 199.595 64.650 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 199.190 64.650 199.510 ;
      LAYER met4 ;
        RECT 64.330 199.190 64.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 198.785 64.650 199.105 ;
      LAYER met4 ;
        RECT 64.330 198.785 64.650 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 198.380 64.650 198.700 ;
      LAYER met4 ;
        RECT 64.330 198.380 64.650 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 197.975 64.650 198.295 ;
      LAYER met4 ;
        RECT 64.330 197.975 64.650 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 197.570 64.650 197.890 ;
      LAYER met4 ;
        RECT 64.330 197.570 64.650 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 197.165 64.650 197.485 ;
      LAYER met4 ;
        RECT 64.330 197.165 64.650 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 196.760 64.650 197.080 ;
      LAYER met4 ;
        RECT 64.330 196.760 64.650 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 196.355 64.650 196.675 ;
      LAYER met4 ;
        RECT 64.330 196.355 64.650 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 195.950 64.650 196.270 ;
      LAYER met4 ;
        RECT 64.330 195.950 64.650 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 195.545 64.650 195.865 ;
      LAYER met4 ;
        RECT 64.330 195.545 64.650 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.330 195.140 64.650 195.460 ;
      LAYER met4 ;
        RECT 64.330 195.140 64.650 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 30.210 64.480 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 29.780 64.480 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 29.350 64.480 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 28.920 64.480 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 28.490 64.480 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 28.060 64.480 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 27.630 64.480 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 27.200 64.480 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 26.770 64.480 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 26.340 64.480 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 25.910 64.480 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 199.595 64.250 199.915 ;
      LAYER met4 ;
        RECT 63.930 199.595 64.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 199.190 64.250 199.510 ;
      LAYER met4 ;
        RECT 63.930 199.190 64.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 198.785 64.250 199.105 ;
      LAYER met4 ;
        RECT 63.930 198.785 64.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 198.380 64.250 198.700 ;
      LAYER met4 ;
        RECT 63.930 198.380 64.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 197.975 64.250 198.295 ;
      LAYER met4 ;
        RECT 63.930 197.975 64.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 197.570 64.250 197.890 ;
      LAYER met4 ;
        RECT 63.930 197.570 64.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 197.165 64.250 197.485 ;
      LAYER met4 ;
        RECT 63.930 197.165 64.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 196.760 64.250 197.080 ;
      LAYER met4 ;
        RECT 63.930 196.760 64.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 196.355 64.250 196.675 ;
      LAYER met4 ;
        RECT 63.930 196.355 64.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 195.950 64.250 196.270 ;
      LAYER met4 ;
        RECT 63.930 195.950 64.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 195.545 64.250 195.865 ;
      LAYER met4 ;
        RECT 63.930 195.545 64.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.930 195.140 64.250 195.460 ;
      LAYER met4 ;
        RECT 63.930 195.140 64.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 30.210 64.075 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 29.780 64.075 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 29.350 64.075 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 28.920 64.075 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 28.490 64.075 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 28.060 64.075 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 27.630 64.075 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 27.200 64.075 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 26.770 64.075 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 26.340 64.075 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 25.910 64.075 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 199.595 63.850 199.915 ;
      LAYER met4 ;
        RECT 63.530 199.595 63.850 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 199.190 63.850 199.510 ;
      LAYER met4 ;
        RECT 63.530 199.190 63.850 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 198.785 63.850 199.105 ;
      LAYER met4 ;
        RECT 63.530 198.785 63.850 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 198.380 63.850 198.700 ;
      LAYER met4 ;
        RECT 63.530 198.380 63.850 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 197.975 63.850 198.295 ;
      LAYER met4 ;
        RECT 63.530 197.975 63.850 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 197.570 63.850 197.890 ;
      LAYER met4 ;
        RECT 63.530 197.570 63.850 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 197.165 63.850 197.485 ;
      LAYER met4 ;
        RECT 63.530 197.165 63.850 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 196.760 63.850 197.080 ;
      LAYER met4 ;
        RECT 63.530 196.760 63.850 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 196.355 63.850 196.675 ;
      LAYER met4 ;
        RECT 63.530 196.355 63.850 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 195.950 63.850 196.270 ;
      LAYER met4 ;
        RECT 63.530 195.950 63.850 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 195.545 63.850 195.865 ;
      LAYER met4 ;
        RECT 63.530 195.545 63.850 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.530 195.140 63.850 195.460 ;
      LAYER met4 ;
        RECT 63.530 195.140 63.850 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 30.210 63.670 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 29.780 63.670 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 29.350 63.670 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 28.920 63.670 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 28.490 63.670 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 28.060 63.670 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 27.630 63.670 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 27.200 63.670 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 26.770 63.670 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 26.340 63.670 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 25.910 63.670 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 199.595 63.450 199.915 ;
      LAYER met4 ;
        RECT 63.130 199.595 63.450 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 199.190 63.450 199.510 ;
      LAYER met4 ;
        RECT 63.130 199.190 63.450 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 198.785 63.450 199.105 ;
      LAYER met4 ;
        RECT 63.130 198.785 63.450 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 198.380 63.450 198.700 ;
      LAYER met4 ;
        RECT 63.130 198.380 63.450 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 197.975 63.450 198.295 ;
      LAYER met4 ;
        RECT 63.130 197.975 63.450 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 197.570 63.450 197.890 ;
      LAYER met4 ;
        RECT 63.130 197.570 63.450 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 197.165 63.450 197.485 ;
      LAYER met4 ;
        RECT 63.130 197.165 63.450 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 196.760 63.450 197.080 ;
      LAYER met4 ;
        RECT 63.130 196.760 63.450 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 196.355 63.450 196.675 ;
      LAYER met4 ;
        RECT 63.130 196.355 63.450 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 195.950 63.450 196.270 ;
      LAYER met4 ;
        RECT 63.130 195.950 63.450 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 195.545 63.450 195.865 ;
      LAYER met4 ;
        RECT 63.130 195.545 63.450 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.130 195.140 63.450 195.460 ;
      LAYER met4 ;
        RECT 63.130 195.140 63.450 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 30.210 63.265 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 29.780 63.265 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 29.350 63.265 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 28.920 63.265 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 28.490 63.265 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 28.060 63.265 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 27.630 63.265 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 27.200 63.265 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 26.770 63.265 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 26.340 63.265 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 25.910 63.265 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 199.595 63.050 199.915 ;
      LAYER met4 ;
        RECT 62.730 199.595 63.050 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 199.190 63.050 199.510 ;
      LAYER met4 ;
        RECT 62.730 199.190 63.050 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 198.785 63.050 199.105 ;
      LAYER met4 ;
        RECT 62.730 198.785 63.050 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 198.380 63.050 198.700 ;
      LAYER met4 ;
        RECT 62.730 198.380 63.050 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 197.975 63.050 198.295 ;
      LAYER met4 ;
        RECT 62.730 197.975 63.050 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 197.570 63.050 197.890 ;
      LAYER met4 ;
        RECT 62.730 197.570 63.050 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 197.165 63.050 197.485 ;
      LAYER met4 ;
        RECT 62.730 197.165 63.050 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 196.760 63.050 197.080 ;
      LAYER met4 ;
        RECT 62.730 196.760 63.050 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 196.355 63.050 196.675 ;
      LAYER met4 ;
        RECT 62.730 196.355 63.050 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 195.950 63.050 196.270 ;
      LAYER met4 ;
        RECT 62.730 195.950 63.050 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 195.545 63.050 195.865 ;
      LAYER met4 ;
        RECT 62.730 195.545 63.050 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.730 195.140 63.050 195.460 ;
      LAYER met4 ;
        RECT 62.730 195.140 63.050 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 30.210 62.860 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 29.780 62.860 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 29.350 62.860 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 28.920 62.860 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 28.490 62.860 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 28.060 62.860 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 27.630 62.860 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 27.200 62.860 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 26.770 62.860 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 26.340 62.860 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 25.910 62.860 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 199.595 62.650 199.915 ;
      LAYER met4 ;
        RECT 62.330 199.595 62.650 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 199.190 62.650 199.510 ;
      LAYER met4 ;
        RECT 62.330 199.190 62.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 198.785 62.650 199.105 ;
      LAYER met4 ;
        RECT 62.330 198.785 62.650 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 198.380 62.650 198.700 ;
      LAYER met4 ;
        RECT 62.330 198.380 62.650 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 197.975 62.650 198.295 ;
      LAYER met4 ;
        RECT 62.330 197.975 62.650 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 197.570 62.650 197.890 ;
      LAYER met4 ;
        RECT 62.330 197.570 62.650 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 197.165 62.650 197.485 ;
      LAYER met4 ;
        RECT 62.330 197.165 62.650 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 196.760 62.650 197.080 ;
      LAYER met4 ;
        RECT 62.330 196.760 62.650 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 196.355 62.650 196.675 ;
      LAYER met4 ;
        RECT 62.330 196.355 62.650 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 195.950 62.650 196.270 ;
      LAYER met4 ;
        RECT 62.330 195.950 62.650 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 195.545 62.650 195.865 ;
      LAYER met4 ;
        RECT 62.330 195.545 62.650 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.330 195.140 62.650 195.460 ;
      LAYER met4 ;
        RECT 62.330 195.140 62.650 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 30.210 62.455 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 29.780 62.455 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 29.350 62.455 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 28.920 62.455 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 28.490 62.455 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 28.060 62.455 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 27.630 62.455 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 27.200 62.455 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 26.770 62.455 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 26.340 62.455 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 25.910 62.455 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 199.595 62.250 199.915 ;
      LAYER met4 ;
        RECT 61.930 199.595 62.250 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 199.190 62.250 199.510 ;
      LAYER met4 ;
        RECT 61.930 199.190 62.250 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 198.785 62.250 199.105 ;
      LAYER met4 ;
        RECT 61.930 198.785 62.250 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 198.380 62.250 198.700 ;
      LAYER met4 ;
        RECT 61.930 198.380 62.250 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 197.975 62.250 198.295 ;
      LAYER met4 ;
        RECT 61.930 197.975 62.250 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 197.570 62.250 197.890 ;
      LAYER met4 ;
        RECT 61.930 197.570 62.250 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 197.165 62.250 197.485 ;
      LAYER met4 ;
        RECT 61.930 197.165 62.250 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 196.760 62.250 197.080 ;
      LAYER met4 ;
        RECT 61.930 196.760 62.250 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 196.355 62.250 196.675 ;
      LAYER met4 ;
        RECT 61.930 196.355 62.250 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 195.950 62.250 196.270 ;
      LAYER met4 ;
        RECT 61.930 195.950 62.250 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 195.545 62.250 195.865 ;
      LAYER met4 ;
        RECT 61.930 195.545 62.250 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.930 195.140 62.250 195.460 ;
      LAYER met4 ;
        RECT 61.930 195.140 62.250 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 30.210 62.050 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 29.780 62.050 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 29.350 62.050 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 28.920 62.050 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 28.490 62.050 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 28.060 62.050 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 27.630 62.050 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 27.200 62.050 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 26.770 62.050 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 26.340 62.050 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 25.910 62.050 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 199.595 61.850 199.915 ;
      LAYER met4 ;
        RECT 61.530 199.595 61.850 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 199.190 61.850 199.510 ;
      LAYER met4 ;
        RECT 61.530 199.190 61.850 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 198.785 61.850 199.105 ;
      LAYER met4 ;
        RECT 61.530 198.785 61.850 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 198.380 61.850 198.700 ;
      LAYER met4 ;
        RECT 61.530 198.380 61.850 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 197.975 61.850 198.295 ;
      LAYER met4 ;
        RECT 61.530 197.975 61.850 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 197.570 61.850 197.890 ;
      LAYER met4 ;
        RECT 61.530 197.570 61.850 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 197.165 61.850 197.485 ;
      LAYER met4 ;
        RECT 61.530 197.165 61.850 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 196.760 61.850 197.080 ;
      LAYER met4 ;
        RECT 61.530 196.760 61.850 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 196.355 61.850 196.675 ;
      LAYER met4 ;
        RECT 61.530 196.355 61.850 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 195.950 61.850 196.270 ;
      LAYER met4 ;
        RECT 61.530 195.950 61.850 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 195.545 61.850 195.865 ;
      LAYER met4 ;
        RECT 61.530 195.545 61.850 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.530 195.140 61.850 195.460 ;
      LAYER met4 ;
        RECT 61.530 195.140 61.850 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 30.210 61.645 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 29.780 61.645 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 29.350 61.645 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 28.920 61.645 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 28.490 61.645 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 28.060 61.645 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 27.630 61.645 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 27.200 61.645 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 26.770 61.645 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 26.340 61.645 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 25.910 61.645 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.085 197.190 61.320 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 30.210 61.240 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 29.780 61.240 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 29.350 61.240 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 28.920 61.240 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 28.490 61.240 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 28.060 61.240 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 27.630 61.240 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 27.200 61.240 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 26.770 61.240 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 26.340 61.240 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 25.910 61.240 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.850 196.645 61.170 196.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.850 196.235 61.170 196.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 30.210 60.835 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 29.780 60.835 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 29.350 60.835 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 28.920 60.835 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 28.490 60.835 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 28.060 60.835 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 27.630 60.835 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 27.200 60.835 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 26.770 60.835 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 26.340 60.835 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 25.910 60.835 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 30.210 60.430 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 29.780 60.430 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 29.350 60.430 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 28.920 60.430 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 28.490 60.430 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 28.060 60.430 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 27.630 60.430 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 27.200 60.430 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 26.770 60.430 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 26.340 60.430 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 25.910 60.430 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 30.210 60.025 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 29.780 60.025 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 29.350 60.025 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 28.920 60.025 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 28.490 60.025 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 28.060 60.025 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 27.630 60.025 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 27.200 60.025 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 26.770 60.025 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 26.340 60.025 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 25.910 60.025 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 30.210 59.620 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 29.780 59.620 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 29.350 59.620 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 28.920 59.620 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 28.490 59.620 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 28.060 59.620 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 27.630 59.620 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 27.200 59.620 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 26.770 59.620 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 26.340 59.620 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 25.910 59.620 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 30.210 59.215 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 29.780 59.215 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 29.350 59.215 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 28.920 59.215 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 28.490 59.215 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 28.060 59.215 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 27.630 59.215 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 27.200 59.215 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 26.770 59.215 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 26.340 59.215 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 25.910 59.215 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 30.210 58.810 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 29.780 58.810 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 29.350 58.810 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 28.920 58.810 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 28.490 58.810 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 28.060 58.810 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 27.630 58.810 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 27.200 58.810 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 26.770 58.810 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 26.340 58.810 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 25.910 58.810 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 30.210 58.405 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 29.780 58.405 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 29.350 58.405 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 28.920 58.405 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 28.490 58.405 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 28.060 58.405 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 27.630 58.405 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 27.200 58.405 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 26.770 58.405 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 26.340 58.405 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 25.910 58.405 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 30.210 58.000 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 29.780 58.000 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 29.350 58.000 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 28.920 58.000 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 28.490 58.000 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 28.060 58.000 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 27.630 58.000 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 27.200 58.000 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 26.770 58.000 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 26.340 58.000 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 25.910 58.000 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 30.210 57.595 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 29.780 57.595 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 29.350 57.595 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 28.920 57.595 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 28.490 57.595 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 28.060 57.595 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 27.630 57.595 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 27.200 57.595 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 26.770 57.595 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 26.340 57.595 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 25.910 57.595 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 30.210 57.190 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 29.780 57.190 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 29.350 57.190 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 28.920 57.190 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 28.490 57.190 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 28.060 57.190 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 27.630 57.190 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 27.200 57.190 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 26.770 57.190 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 26.340 57.190 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 25.910 57.190 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 30.210 56.785 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 29.780 56.785 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 29.350 56.785 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 28.920 56.785 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 28.490 56.785 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 28.060 56.785 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 27.630 56.785 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 27.200 56.785 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 26.770 56.785 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 26.340 56.785 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 25.910 56.785 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 30.210 56.380 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 29.780 56.380 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 29.350 56.380 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 28.920 56.380 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 28.490 56.380 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 28.060 56.380 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 27.630 56.380 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 27.200 56.380 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 26.770 56.380 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 26.340 56.380 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.180 25.910 56.380 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 30.210 55.975 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 29.780 55.975 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 29.350 55.975 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 28.920 55.975 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 28.490 55.975 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 28.060 55.975 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 27.630 55.975 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 27.200 55.975 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 26.770 55.975 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 26.340 55.975 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.775 25.910 55.975 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 30.210 55.570 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 29.780 55.570 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 29.350 55.570 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 28.920 55.570 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 28.490 55.570 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 28.060 55.570 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 27.630 55.570 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 27.200 55.570 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 26.770 55.570 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 26.340 55.570 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.370 25.910 55.570 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 30.210 55.165 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 29.780 55.165 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 29.350 55.165 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 28.920 55.165 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 28.490 55.165 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 28.060 55.165 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 27.630 55.165 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 27.200 55.165 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 26.770 55.165 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 26.340 55.165 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.965 25.910 55.165 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 30.210 54.760 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 29.780 54.760 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 29.350 54.760 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 28.920 54.760 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 28.490 54.760 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 28.060 54.760 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 27.630 54.760 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 27.200 54.760 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 26.770 54.760 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 26.340 54.760 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.560 25.910 54.760 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 30.210 54.355 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 29.780 54.355 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 29.350 54.355 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 28.920 54.355 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 28.490 54.355 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 28.060 54.355 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 27.630 54.355 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 27.200 54.355 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 26.770 54.355 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 26.340 54.355 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.155 25.910 54.355 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 30.210 53.950 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 29.780 53.950 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 29.350 53.950 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 28.920 53.950 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 28.490 53.950 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 28.060 53.950 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 27.630 53.950 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 27.200 53.950 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 26.770 53.950 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 26.340 53.950 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.750 25.910 53.950 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 30.210 53.545 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 29.780 53.545 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 29.350 53.545 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 28.920 53.545 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 28.490 53.545 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 28.060 53.545 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 27.630 53.545 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 27.200 53.545 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 26.770 53.545 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 26.340 53.545 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.345 25.910 53.545 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 30.210 53.140 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 29.780 53.140 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 29.350 53.140 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 28.920 53.140 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 28.490 53.140 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 28.060 53.140 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 27.630 53.140 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 27.200 53.140 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 26.770 53.140 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 26.340 53.140 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.940 25.910 53.140 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 30.210 52.730 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 29.780 52.730 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 29.350 52.730 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 28.920 52.730 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 28.490 52.730 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 28.060 52.730 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 27.630 52.730 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 27.200 52.730 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 26.770 52.730 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 26.340 52.730 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.530 25.910 52.730 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 30.210 52.320 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 29.780 52.320 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 29.350 52.320 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 28.920 52.320 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 28.490 52.320 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 28.060 52.320 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 27.630 52.320 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 27.200 52.320 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 26.770 52.320 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 26.340 52.320 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.120 25.910 52.320 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 30.210 51.910 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 29.780 51.910 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 29.350 51.910 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 28.920 51.910 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 28.490 51.910 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 28.060 51.910 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 27.630 51.910 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 27.200 51.910 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 26.770 51.910 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 26.340 51.910 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.710 25.910 51.910 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 30.210 51.500 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 29.780 51.500 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 29.350 51.500 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 28.920 51.500 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 28.490 51.500 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 28.060 51.500 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 27.630 51.500 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 27.200 51.500 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 26.770 51.500 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 26.340 51.500 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.300 25.910 51.500 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 30.210 51.090 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 29.780 51.090 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 29.350 51.090 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 28.920 51.090 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 28.490 51.090 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 28.060 51.090 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 27.630 51.090 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 27.200 51.090 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 26.770 51.090 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 26.340 51.090 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.890 25.910 51.090 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 30.210 50.680 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 29.780 50.680 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 29.350 50.680 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 28.920 50.680 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 28.490 50.680 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 28.060 50.680 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 27.630 50.680 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 27.200 50.680 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 26.770 50.680 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 26.340 50.680 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.480 25.910 50.680 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.000 197.190 37.085 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 199.590 26.915 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 199.190 26.915 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 198.790 26.915 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 198.390 26.915 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 197.990 26.915 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 197.590 26.915 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.595 197.190 26.915 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 199.590 26.510 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 199.190 26.510 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 198.790 26.510 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 198.390 26.510 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 197.990 26.510 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 197.590 26.510 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.190 197.190 26.510 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 199.590 26.105 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 199.190 26.105 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 198.790 26.105 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 198.390 26.105 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 197.990 26.105 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 197.590 26.105 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.785 197.190 26.105 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 199.590 25.700 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 199.190 25.700 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 198.790 25.700 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 198.390 25.700 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 197.990 25.700 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 197.590 25.700 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.380 197.190 25.700 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 199.590 25.295 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 199.190 25.295 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 198.790 25.295 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 198.390 25.295 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 197.990 25.295 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 197.590 25.295 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.975 197.190 25.295 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 199.590 24.890 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 199.190 24.890 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 198.790 24.890 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 198.390 24.890 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 197.990 24.890 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 197.590 24.890 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.570 197.190 24.890 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 199.590 24.485 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 199.190 24.485 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 198.790 24.485 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 198.390 24.485 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 197.990 24.485 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 197.590 24.485 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.165 197.190 24.485 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 30.210 24.305 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 29.780 24.305 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 29.350 24.305 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 28.920 24.305 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 28.490 24.305 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 28.060 24.305 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 27.630 24.305 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 27.200 24.305 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 26.770 24.305 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 26.340 24.305 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.105 25.910 24.305 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 199.590 24.080 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 199.190 24.080 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 198.790 24.080 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 198.390 24.080 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 197.990 24.080 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 197.590 24.080 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.760 197.190 24.080 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 30.210 23.900 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 29.780 23.900 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 29.350 23.900 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 28.920 23.900 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 28.490 23.900 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 28.060 23.900 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 27.630 23.900 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 27.200 23.900 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 26.770 23.900 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 26.340 23.900 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.700 25.910 23.900 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 199.590 23.675 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 199.190 23.675 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 198.790 23.675 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 198.390 23.675 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 197.990 23.675 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 197.590 23.675 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.355 197.190 23.675 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 30.210 23.495 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 29.780 23.495 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 29.350 23.495 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 28.920 23.495 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 28.490 23.495 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 28.060 23.495 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 27.630 23.495 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 27.200 23.495 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 26.770 23.495 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 26.340 23.495 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.295 25.910 23.495 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 199.590 23.270 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 199.190 23.270 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 198.790 23.270 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 198.390 23.270 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 197.990 23.270 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 197.590 23.270 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.950 197.190 23.270 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 30.210 23.090 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 29.780 23.090 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 29.350 23.090 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 28.920 23.090 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 28.490 23.090 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 28.060 23.090 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 27.630 23.090 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 27.200 23.090 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 26.770 23.090 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 26.340 23.090 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.890 25.910 23.090 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 199.590 22.865 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 199.190 22.865 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 198.790 22.865 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 198.390 22.865 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 197.990 22.865 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 197.590 22.865 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.545 197.190 22.865 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 30.210 22.685 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 29.780 22.685 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 29.350 22.685 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 28.920 22.685 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 28.490 22.685 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 28.060 22.685 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 27.630 22.685 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 27.200 22.685 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 26.770 22.685 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 26.340 22.685 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.485 25.910 22.685 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 199.590 22.460 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 199.190 22.460 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 198.790 22.460 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 198.390 22.460 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 197.990 22.460 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 197.590 22.460 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.140 197.190 22.460 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 30.210 22.280 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 29.780 22.280 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 29.350 22.280 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 28.920 22.280 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 28.490 22.280 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 28.060 22.280 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 27.630 22.280 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 27.200 22.280 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 26.770 22.280 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 26.340 22.280 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.080 25.910 22.280 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 199.590 22.055 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 199.190 22.055 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 198.790 22.055 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 198.390 22.055 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 197.990 22.055 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 197.590 22.055 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.735 197.190 22.055 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 30.210 21.875 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 29.780 21.875 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 29.350 21.875 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 28.920 21.875 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 28.490 21.875 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 28.060 21.875 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 27.630 21.875 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 27.200 21.875 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 26.770 21.875 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 26.340 21.875 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.675 25.910 21.875 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 199.590 21.650 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 199.190 21.650 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 198.790 21.650 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 198.390 21.650 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 197.990 21.650 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 197.590 21.650 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.330 197.190 21.650 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 30.210 21.470 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 29.780 21.470 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 29.350 21.470 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 28.920 21.470 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 28.490 21.470 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 28.060 21.470 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 27.630 21.470 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 27.200 21.470 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 26.770 21.470 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 26.340 21.470 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.270 25.910 21.470 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 199.590 21.245 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 199.190 21.245 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 198.790 21.245 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 198.390 21.245 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 197.990 21.245 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 197.590 21.245 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.925 197.190 21.245 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 30.210 21.065 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 29.780 21.065 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 29.350 21.065 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 28.920 21.065 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 28.490 21.065 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 28.060 21.065 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 27.630 21.065 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 27.200 21.065 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 26.770 21.065 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 26.340 21.065 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.865 25.910 21.065 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 199.590 20.840 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 199.190 20.840 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 198.790 20.840 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 198.390 20.840 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 197.990 20.840 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 197.590 20.840 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.520 197.190 20.840 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 30.210 20.660 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 29.780 20.660 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 29.350 20.660 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 28.920 20.660 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 28.490 20.660 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 28.060 20.660 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 27.630 20.660 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 27.200 20.660 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 26.770 20.660 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 26.340 20.660 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.460 25.910 20.660 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 199.590 20.435 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 199.190 20.435 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 198.790 20.435 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 198.390 20.435 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 197.990 20.435 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 197.590 20.435 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.115 197.190 20.435 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 30.210 20.255 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 29.780 20.255 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 29.350 20.255 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 28.920 20.255 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 28.490 20.255 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 28.060 20.255 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 27.630 20.255 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 27.200 20.255 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 26.770 20.255 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 26.340 20.255 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.055 25.910 20.255 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 199.590 20.030 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 199.190 20.030 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 198.790 20.030 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 198.390 20.030 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 197.990 20.030 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 197.590 20.030 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.710 197.190 20.030 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 30.210 19.850 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 29.780 19.850 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 29.350 19.850 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 28.920 19.850 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 28.490 19.850 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 28.060 19.850 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 27.630 19.850 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 27.200 19.850 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 26.770 19.850 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 26.340 19.850 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.650 25.910 19.850 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 199.590 19.625 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 199.190 19.625 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 198.790 19.625 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 198.390 19.625 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 197.990 19.625 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 197.590 19.625 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.305 197.190 19.625 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 30.210 19.445 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 29.780 19.445 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 29.350 19.445 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 28.920 19.445 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 28.490 19.445 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 28.060 19.445 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 27.630 19.445 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 27.200 19.445 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 26.770 19.445 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 26.340 19.445 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 25.910 19.445 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 199.590 19.220 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 199.190 19.220 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 198.790 19.220 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 198.390 19.220 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 197.990 19.220 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 197.590 19.220 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.900 197.190 19.220 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 30.210 19.040 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 29.780 19.040 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 29.350 19.040 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 28.920 19.040 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 28.490 19.040 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 28.060 19.040 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 27.630 19.040 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 27.200 19.040 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 26.770 19.040 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 26.340 19.040 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.840 25.910 19.040 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 199.590 18.815 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 199.190 18.815 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 198.790 18.815 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 198.390 18.815 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 197.990 18.815 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 197.590 18.815 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 197.190 18.815 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 30.210 18.635 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 29.780 18.635 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 29.350 18.635 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 28.920 18.635 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 28.490 18.635 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 28.060 18.635 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 27.630 18.635 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 27.200 18.635 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 26.770 18.635 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 26.340 18.635 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.435 25.910 18.635 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 199.590 18.410 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 199.190 18.410 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 198.790 18.410 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 198.390 18.410 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 197.990 18.410 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 197.590 18.410 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.090 197.190 18.410 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 30.210 18.230 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 29.780 18.230 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 29.350 18.230 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 28.920 18.230 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 28.490 18.230 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 28.060 18.230 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 27.630 18.230 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 27.200 18.230 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 26.770 18.230 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 26.340 18.230 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.030 25.910 18.230 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 199.590 18.005 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 199.190 18.005 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 198.790 18.005 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 198.390 18.005 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 197.990 18.005 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 197.590 18.005 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.685 197.190 18.005 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 30.210 17.825 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 29.780 17.825 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 29.350 17.825 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 28.920 17.825 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 28.490 17.825 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 28.060 17.825 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 27.630 17.825 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 27.200 17.825 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 26.770 17.825 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 26.340 17.825 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.625 25.910 17.825 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 199.590 17.600 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 199.190 17.600 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 198.790 17.600 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 198.390 17.600 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 197.990 17.600 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 197.590 17.600 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.280 197.190 17.600 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 30.210 17.420 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 29.780 17.420 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 29.350 17.420 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 28.920 17.420 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 28.490 17.420 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 28.060 17.420 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 27.630 17.420 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 27.200 17.420 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 26.770 17.420 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 26.340 17.420 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.220 25.910 17.420 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 199.590 17.195 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 199.190 17.195 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 198.790 17.195 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 198.390 17.195 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 197.990 17.195 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 197.590 17.195 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.875 197.190 17.195 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 30.210 17.015 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 29.780 17.015 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 29.350 17.015 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 28.920 17.015 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 28.490 17.015 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 28.060 17.015 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 27.630 17.015 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 27.200 17.015 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 26.770 17.015 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 26.340 17.015 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.815 25.910 17.015 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 199.590 16.790 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 199.190 16.790 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 198.790 16.790 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 198.390 16.790 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 197.990 16.790 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 197.590 16.790 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.470 197.190 16.790 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 30.210 16.610 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 29.780 16.610 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 29.350 16.610 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 28.920 16.610 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 28.490 16.610 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 28.060 16.610 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 27.630 16.610 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 27.200 16.610 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 26.770 16.610 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 26.340 16.610 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.410 25.910 16.610 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 199.590 16.385 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 199.190 16.385 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 198.790 16.385 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 198.390 16.385 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 197.990 16.385 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 197.590 16.385 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.065 197.190 16.385 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 30.210 16.205 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 29.780 16.205 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 29.350 16.205 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 28.920 16.205 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 28.490 16.205 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 28.060 16.205 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 27.630 16.205 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 27.200 16.205 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 26.770 16.205 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 26.340 16.205 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.005 25.910 16.205 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 199.590 15.980 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 199.190 15.980 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 198.790 15.980 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 198.390 15.980 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 197.990 15.980 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 197.590 15.980 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.660 197.190 15.980 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 30.210 15.800 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 29.780 15.800 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 29.350 15.800 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 28.920 15.800 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 28.490 15.800 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 28.060 15.800 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 27.630 15.800 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 27.200 15.800 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 26.770 15.800 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 26.340 15.800 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.600 25.910 15.800 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 199.590 15.575 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 199.190 15.575 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 198.790 15.575 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 198.390 15.575 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 197.990 15.575 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 197.590 15.575 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.255 197.190 15.575 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 30.210 15.395 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 29.780 15.395 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 29.350 15.395 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 28.920 15.395 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 28.490 15.395 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 28.060 15.395 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 27.630 15.395 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 27.200 15.395 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 26.770 15.395 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 26.340 15.395 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.195 25.910 15.395 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 199.590 15.170 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 199.190 15.170 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 198.790 15.170 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 198.390 15.170 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 197.990 15.170 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 197.590 15.170 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.850 197.190 15.170 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 30.210 14.990 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 29.780 14.990 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 29.350 14.990 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 28.920 14.990 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 28.490 14.990 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 28.060 14.990 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 27.630 14.990 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 27.200 14.990 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 26.770 14.990 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 26.340 14.990 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.790 25.910 14.990 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 199.590 14.765 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 199.190 14.765 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 198.790 14.765 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 198.390 14.765 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 197.990 14.765 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 197.590 14.765 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.445 197.190 14.765 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 30.210 14.585 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 29.780 14.585 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 29.350 14.585 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 28.920 14.585 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 28.490 14.585 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 28.060 14.585 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 27.630 14.585 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 27.200 14.585 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 26.770 14.585 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 26.340 14.585 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.385 25.910 14.585 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 199.590 14.360 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 199.190 14.360 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 198.790 14.360 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 198.390 14.360 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 197.990 14.360 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 197.590 14.360 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.040 197.190 14.360 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 30.210 14.180 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 29.780 14.180 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 29.350 14.180 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 28.920 14.180 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 28.490 14.180 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 28.060 14.180 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 27.630 14.180 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 27.200 14.180 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 26.770 14.180 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 26.340 14.180 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.980 25.910 14.180 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.765 196.645 14.085 196.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.765 196.235 14.085 196.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 199.590 13.955 199.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 199.190 13.955 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 198.790 13.955 199.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 198.390 13.955 198.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 197.990 13.955 198.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 197.590 13.955 197.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.635 197.190 13.955 197.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 30.210 13.775 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 29.780 13.775 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 29.350 13.775 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 28.920 13.775 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 28.490 13.775 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 28.060 13.775 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 27.630 13.775 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 27.200 13.775 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 26.770 13.775 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 26.340 13.775 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.575 25.910 13.775 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 30.210 13.370 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 29.780 13.370 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 29.350 13.370 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 28.920 13.370 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 28.490 13.370 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 28.060 13.370 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 27.630 13.370 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 27.200 13.370 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 26.770 13.370 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 26.340 13.370 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.170 25.910 13.370 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 199.595 13.345 199.915 ;
      LAYER met4 ;
        RECT 13.025 199.595 13.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 199.190 13.345 199.510 ;
      LAYER met4 ;
        RECT 13.025 199.190 13.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 198.785 13.345 199.105 ;
      LAYER met4 ;
        RECT 13.025 198.785 13.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 198.380 13.345 198.700 ;
      LAYER met4 ;
        RECT 13.025 198.380 13.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 197.975 13.345 198.295 ;
      LAYER met4 ;
        RECT 13.025 197.975 13.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 197.570 13.345 197.890 ;
      LAYER met4 ;
        RECT 13.025 197.570 13.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 197.165 13.345 197.485 ;
      LAYER met4 ;
        RECT 13.025 197.165 13.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 196.760 13.345 197.080 ;
      LAYER met4 ;
        RECT 13.025 196.760 13.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 196.355 13.345 196.675 ;
      LAYER met4 ;
        RECT 13.025 196.355 13.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 195.950 13.345 196.270 ;
      LAYER met4 ;
        RECT 13.025 195.950 13.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 195.545 13.345 195.865 ;
      LAYER met4 ;
        RECT 13.025 195.545 13.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.025 195.140 13.345 195.460 ;
      LAYER met4 ;
        RECT 13.025 195.140 13.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 175.935 13.345 195.055 ;
      LAYER met4 ;
        RECT 1.270 175.935 13.345 195.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 30.210 12.965 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 29.780 12.965 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 29.350 12.965 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 28.920 12.965 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 28.490 12.965 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 28.060 12.965 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 27.630 12.965 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 27.200 12.965 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 26.770 12.965 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 26.340 12.965 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.765 25.910 12.965 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 199.595 12.945 199.915 ;
      LAYER met4 ;
        RECT 12.625 199.595 12.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 199.190 12.945 199.510 ;
      LAYER met4 ;
        RECT 12.625 199.190 12.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 198.785 12.945 199.105 ;
      LAYER met4 ;
        RECT 12.625 198.785 12.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 198.380 12.945 198.700 ;
      LAYER met4 ;
        RECT 12.625 198.380 12.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 197.975 12.945 198.295 ;
      LAYER met4 ;
        RECT 12.625 197.975 12.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 197.570 12.945 197.890 ;
      LAYER met4 ;
        RECT 12.625 197.570 12.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 197.165 12.945 197.485 ;
      LAYER met4 ;
        RECT 12.625 197.165 12.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 196.760 12.945 197.080 ;
      LAYER met4 ;
        RECT 12.625 196.760 12.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 196.355 12.945 196.675 ;
      LAYER met4 ;
        RECT 12.625 196.355 12.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 195.950 12.945 196.270 ;
      LAYER met4 ;
        RECT 12.625 195.950 12.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 195.545 12.945 195.865 ;
      LAYER met4 ;
        RECT 12.625 195.545 12.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.625 195.140 12.945 195.460 ;
      LAYER met4 ;
        RECT 12.625 195.140 12.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 30.210 12.560 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 29.780 12.560 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 29.350 12.560 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 28.920 12.560 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 28.490 12.560 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 28.060 12.560 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 27.630 12.560 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 27.200 12.560 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 26.770 12.560 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 26.340 12.560 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.360 25.910 12.560 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 199.595 12.545 199.915 ;
      LAYER met4 ;
        RECT 12.225 199.595 12.545 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 199.190 12.545 199.510 ;
      LAYER met4 ;
        RECT 12.225 199.190 12.545 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 198.785 12.545 199.105 ;
      LAYER met4 ;
        RECT 12.225 198.785 12.545 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 198.380 12.545 198.700 ;
      LAYER met4 ;
        RECT 12.225 198.380 12.545 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 197.975 12.545 198.295 ;
      LAYER met4 ;
        RECT 12.225 197.975 12.545 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 197.570 12.545 197.890 ;
      LAYER met4 ;
        RECT 12.225 197.570 12.545 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 197.165 12.545 197.485 ;
      LAYER met4 ;
        RECT 12.225 197.165 12.545 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 196.760 12.545 197.080 ;
      LAYER met4 ;
        RECT 12.225 196.760 12.545 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 196.355 12.545 196.675 ;
      LAYER met4 ;
        RECT 12.225 196.355 12.545 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 195.950 12.545 196.270 ;
      LAYER met4 ;
        RECT 12.225 195.950 12.545 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 195.545 12.545 195.865 ;
      LAYER met4 ;
        RECT 12.225 195.545 12.545 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.225 195.140 12.545 195.460 ;
      LAYER met4 ;
        RECT 12.225 195.140 12.545 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 30.210 12.155 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 29.780 12.155 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 29.350 12.155 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 28.920 12.155 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 28.490 12.155 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 28.060 12.155 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 27.630 12.155 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 27.200 12.155 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 26.770 12.155 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 26.340 12.155 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.955 25.910 12.155 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 199.595 12.145 199.915 ;
      LAYER met4 ;
        RECT 11.825 199.595 12.145 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 199.190 12.145 199.510 ;
      LAYER met4 ;
        RECT 11.825 199.190 12.145 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 198.785 12.145 199.105 ;
      LAYER met4 ;
        RECT 11.825 198.785 12.145 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 198.380 12.145 198.700 ;
      LAYER met4 ;
        RECT 11.825 198.380 12.145 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 197.975 12.145 198.295 ;
      LAYER met4 ;
        RECT 11.825 197.975 12.145 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 197.570 12.145 197.890 ;
      LAYER met4 ;
        RECT 11.825 197.570 12.145 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 197.165 12.145 197.485 ;
      LAYER met4 ;
        RECT 11.825 197.165 12.145 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 196.760 12.145 197.080 ;
      LAYER met4 ;
        RECT 11.825 196.760 12.145 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 196.355 12.145 196.675 ;
      LAYER met4 ;
        RECT 11.825 196.355 12.145 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 195.950 12.145 196.270 ;
      LAYER met4 ;
        RECT 11.825 195.950 12.145 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 195.545 12.145 195.865 ;
      LAYER met4 ;
        RECT 11.825 195.545 12.145 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.825 195.140 12.145 195.460 ;
      LAYER met4 ;
        RECT 11.825 195.140 12.145 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 30.210 11.750 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 29.780 11.750 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 29.350 11.750 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 28.920 11.750 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 28.490 11.750 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 28.060 11.750 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 27.630 11.750 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 27.200 11.750 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 26.770 11.750 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 26.340 11.750 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.550 25.910 11.750 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 199.595 11.745 199.915 ;
      LAYER met4 ;
        RECT 11.425 199.595 11.745 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 199.190 11.745 199.510 ;
      LAYER met4 ;
        RECT 11.425 199.190 11.745 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 198.785 11.745 199.105 ;
      LAYER met4 ;
        RECT 11.425 198.785 11.745 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 198.380 11.745 198.700 ;
      LAYER met4 ;
        RECT 11.425 198.380 11.745 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 197.975 11.745 198.295 ;
      LAYER met4 ;
        RECT 11.425 197.975 11.745 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 197.570 11.745 197.890 ;
      LAYER met4 ;
        RECT 11.425 197.570 11.745 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 197.165 11.745 197.485 ;
      LAYER met4 ;
        RECT 11.425 197.165 11.745 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 196.760 11.745 197.080 ;
      LAYER met4 ;
        RECT 11.425 196.760 11.745 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 196.355 11.745 196.675 ;
      LAYER met4 ;
        RECT 11.425 196.355 11.745 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 195.950 11.745 196.270 ;
      LAYER met4 ;
        RECT 11.425 195.950 11.745 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 195.545 11.745 195.865 ;
      LAYER met4 ;
        RECT 11.425 195.545 11.745 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.425 195.140 11.745 195.460 ;
      LAYER met4 ;
        RECT 11.425 195.140 11.745 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 30.210 11.345 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 29.780 11.345 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 29.350 11.345 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 28.920 11.345 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 28.490 11.345 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 28.060 11.345 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 27.630 11.345 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 27.200 11.345 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 26.770 11.345 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 26.340 11.345 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.145 25.910 11.345 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 199.595 11.345 199.915 ;
      LAYER met4 ;
        RECT 11.025 199.595 11.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 199.190 11.345 199.510 ;
      LAYER met4 ;
        RECT 11.025 199.190 11.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 198.785 11.345 199.105 ;
      LAYER met4 ;
        RECT 11.025 198.785 11.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 198.380 11.345 198.700 ;
      LAYER met4 ;
        RECT 11.025 198.380 11.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 197.975 11.345 198.295 ;
      LAYER met4 ;
        RECT 11.025 197.975 11.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 197.570 11.345 197.890 ;
      LAYER met4 ;
        RECT 11.025 197.570 11.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 197.165 11.345 197.485 ;
      LAYER met4 ;
        RECT 11.025 197.165 11.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 196.760 11.345 197.080 ;
      LAYER met4 ;
        RECT 11.025 196.760 11.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 196.355 11.345 196.675 ;
      LAYER met4 ;
        RECT 11.025 196.355 11.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 195.950 11.345 196.270 ;
      LAYER met4 ;
        RECT 11.025 195.950 11.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 195.545 11.345 195.865 ;
      LAYER met4 ;
        RECT 11.025 195.545 11.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.025 195.140 11.345 195.460 ;
      LAYER met4 ;
        RECT 11.025 195.140 11.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 30.210 10.940 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 29.780 10.940 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 29.350 10.940 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 28.920 10.940 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 28.490 10.940 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 28.060 10.940 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 27.630 10.940 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 27.200 10.940 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 26.770 10.940 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 26.340 10.940 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.740 25.910 10.940 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 199.595 10.945 199.915 ;
      LAYER met4 ;
        RECT 10.625 199.595 10.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 199.190 10.945 199.510 ;
      LAYER met4 ;
        RECT 10.625 199.190 10.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 198.785 10.945 199.105 ;
      LAYER met4 ;
        RECT 10.625 198.785 10.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 198.380 10.945 198.700 ;
      LAYER met4 ;
        RECT 10.625 198.380 10.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 197.975 10.945 198.295 ;
      LAYER met4 ;
        RECT 10.625 197.975 10.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 197.570 10.945 197.890 ;
      LAYER met4 ;
        RECT 10.625 197.570 10.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 197.165 10.945 197.485 ;
      LAYER met4 ;
        RECT 10.625 197.165 10.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 196.760 10.945 197.080 ;
      LAYER met4 ;
        RECT 10.625 196.760 10.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 196.355 10.945 196.675 ;
      LAYER met4 ;
        RECT 10.625 196.355 10.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 195.950 10.945 196.270 ;
      LAYER met4 ;
        RECT 10.625 195.950 10.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 195.545 10.945 195.865 ;
      LAYER met4 ;
        RECT 10.625 195.545 10.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.625 195.140 10.945 195.460 ;
      LAYER met4 ;
        RECT 10.625 195.140 10.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 30.210 10.535 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 29.780 10.535 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 29.350 10.535 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 28.920 10.535 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 28.490 10.535 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 28.060 10.535 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 27.630 10.535 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 27.200 10.535 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 26.770 10.535 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 26.340 10.535 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.335 25.910 10.535 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 199.595 10.545 199.915 ;
      LAYER met4 ;
        RECT 10.225 199.595 10.545 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 199.190 10.545 199.510 ;
      LAYER met4 ;
        RECT 10.225 199.190 10.545 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 198.785 10.545 199.105 ;
      LAYER met4 ;
        RECT 10.225 198.785 10.545 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 198.380 10.545 198.700 ;
      LAYER met4 ;
        RECT 10.225 198.380 10.545 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 197.975 10.545 198.295 ;
      LAYER met4 ;
        RECT 10.225 197.975 10.545 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 197.570 10.545 197.890 ;
      LAYER met4 ;
        RECT 10.225 197.570 10.545 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 197.165 10.545 197.485 ;
      LAYER met4 ;
        RECT 10.225 197.165 10.545 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 196.760 10.545 197.080 ;
      LAYER met4 ;
        RECT 10.225 196.760 10.545 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 196.355 10.545 196.675 ;
      LAYER met4 ;
        RECT 10.225 196.355 10.545 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 195.950 10.545 196.270 ;
      LAYER met4 ;
        RECT 10.225 195.950 10.545 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 195.545 10.545 195.865 ;
      LAYER met4 ;
        RECT 10.225 195.545 10.545 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.225 195.140 10.545 195.460 ;
      LAYER met4 ;
        RECT 10.225 195.140 10.545 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 30.210 10.130 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 29.780 10.130 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 29.350 10.130 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 28.920 10.130 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 28.490 10.130 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 28.060 10.130 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 27.630 10.130 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 27.200 10.130 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 26.770 10.130 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 26.340 10.130 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.930 25.910 10.130 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 199.595 10.145 199.915 ;
      LAYER met4 ;
        RECT 9.825 199.595 10.145 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 199.190 10.145 199.510 ;
      LAYER met4 ;
        RECT 9.825 199.190 10.145 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 198.785 10.145 199.105 ;
      LAYER met4 ;
        RECT 9.825 198.785 10.145 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 198.380 10.145 198.700 ;
      LAYER met4 ;
        RECT 9.825 198.380 10.145 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 197.975 10.145 198.295 ;
      LAYER met4 ;
        RECT 9.825 197.975 10.145 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 197.570 10.145 197.890 ;
      LAYER met4 ;
        RECT 9.825 197.570 10.145 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 197.165 10.145 197.485 ;
      LAYER met4 ;
        RECT 9.825 197.165 10.145 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 196.760 10.145 197.080 ;
      LAYER met4 ;
        RECT 9.825 196.760 10.145 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 196.355 10.145 196.675 ;
      LAYER met4 ;
        RECT 9.825 196.355 10.145 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 195.950 10.145 196.270 ;
      LAYER met4 ;
        RECT 9.825 195.950 10.145 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 195.545 10.145 195.865 ;
      LAYER met4 ;
        RECT 9.825 195.545 10.145 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.825 195.140 10.145 195.460 ;
      LAYER met4 ;
        RECT 9.825 195.140 10.145 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 30.210 9.725 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 29.780 9.725 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 29.350 9.725 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 28.920 9.725 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 28.490 9.725 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 28.060 9.725 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 27.630 9.725 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 27.200 9.725 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 26.770 9.725 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 26.340 9.725 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.525 25.910 9.725 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 199.595 9.745 199.915 ;
      LAYER met4 ;
        RECT 9.425 199.595 9.745 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 199.190 9.745 199.510 ;
      LAYER met4 ;
        RECT 9.425 199.190 9.745 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 198.785 9.745 199.105 ;
      LAYER met4 ;
        RECT 9.425 198.785 9.745 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 198.380 9.745 198.700 ;
      LAYER met4 ;
        RECT 9.425 198.380 9.745 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 197.975 9.745 198.295 ;
      LAYER met4 ;
        RECT 9.425 197.975 9.745 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 197.570 9.745 197.890 ;
      LAYER met4 ;
        RECT 9.425 197.570 9.745 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 197.165 9.745 197.485 ;
      LAYER met4 ;
        RECT 9.425 197.165 9.745 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 196.760 9.745 197.080 ;
      LAYER met4 ;
        RECT 9.425 196.760 9.745 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 196.355 9.745 196.675 ;
      LAYER met4 ;
        RECT 9.425 196.355 9.745 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 195.950 9.745 196.270 ;
      LAYER met4 ;
        RECT 9.425 195.950 9.745 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 195.545 9.745 195.865 ;
      LAYER met4 ;
        RECT 9.425 195.545 9.745 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.425 195.140 9.745 195.460 ;
      LAYER met4 ;
        RECT 9.425 195.140 9.745 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 30.210 9.320 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 29.780 9.320 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 29.350 9.320 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 28.920 9.320 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 28.490 9.320 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 28.060 9.320 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 27.630 9.320 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 27.200 9.320 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 26.770 9.320 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 26.340 9.320 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.120 25.910 9.320 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 199.595 9.345 199.915 ;
      LAYER met4 ;
        RECT 9.025 199.595 9.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 199.190 9.345 199.510 ;
      LAYER met4 ;
        RECT 9.025 199.190 9.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 198.785 9.345 199.105 ;
      LAYER met4 ;
        RECT 9.025 198.785 9.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 198.380 9.345 198.700 ;
      LAYER met4 ;
        RECT 9.025 198.380 9.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 197.975 9.345 198.295 ;
      LAYER met4 ;
        RECT 9.025 197.975 9.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 197.570 9.345 197.890 ;
      LAYER met4 ;
        RECT 9.025 197.570 9.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 197.165 9.345 197.485 ;
      LAYER met4 ;
        RECT 9.025 197.165 9.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 196.760 9.345 197.080 ;
      LAYER met4 ;
        RECT 9.025 196.760 9.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 196.355 9.345 196.675 ;
      LAYER met4 ;
        RECT 9.025 196.355 9.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 195.950 9.345 196.270 ;
      LAYER met4 ;
        RECT 9.025 195.950 9.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 195.545 9.345 195.865 ;
      LAYER met4 ;
        RECT 9.025 195.545 9.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.025 195.140 9.345 195.460 ;
      LAYER met4 ;
        RECT 9.025 195.140 9.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 30.210 8.915 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 29.780 8.915 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 29.350 8.915 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 28.920 8.915 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 28.490 8.915 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 28.060 8.915 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 27.630 8.915 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 27.200 8.915 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 26.770 8.915 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 26.340 8.915 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.715 25.910 8.915 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 199.595 8.945 199.915 ;
      LAYER met4 ;
        RECT 8.625 199.595 8.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 199.190 8.945 199.510 ;
      LAYER met4 ;
        RECT 8.625 199.190 8.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 198.785 8.945 199.105 ;
      LAYER met4 ;
        RECT 8.625 198.785 8.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 198.380 8.945 198.700 ;
      LAYER met4 ;
        RECT 8.625 198.380 8.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 197.975 8.945 198.295 ;
      LAYER met4 ;
        RECT 8.625 197.975 8.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 197.570 8.945 197.890 ;
      LAYER met4 ;
        RECT 8.625 197.570 8.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 197.165 8.945 197.485 ;
      LAYER met4 ;
        RECT 8.625 197.165 8.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 196.760 8.945 197.080 ;
      LAYER met4 ;
        RECT 8.625 196.760 8.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 196.355 8.945 196.675 ;
      LAYER met4 ;
        RECT 8.625 196.355 8.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 195.950 8.945 196.270 ;
      LAYER met4 ;
        RECT 8.625 195.950 8.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 195.545 8.945 195.865 ;
      LAYER met4 ;
        RECT 8.625 195.545 8.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.625 195.140 8.945 195.460 ;
      LAYER met4 ;
        RECT 8.625 195.140 8.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 30.210 8.510 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 29.780 8.510 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 29.350 8.510 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 28.920 8.510 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 28.490 8.510 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 28.060 8.510 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 27.630 8.510 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 27.200 8.510 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 26.770 8.510 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 26.340 8.510 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.310 25.910 8.510 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 199.595 8.545 199.915 ;
      LAYER met4 ;
        RECT 8.225 199.595 8.545 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 199.190 8.545 199.510 ;
      LAYER met4 ;
        RECT 8.225 199.190 8.545 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 198.785 8.545 199.105 ;
      LAYER met4 ;
        RECT 8.225 198.785 8.545 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 198.380 8.545 198.700 ;
      LAYER met4 ;
        RECT 8.225 198.380 8.545 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 197.975 8.545 198.295 ;
      LAYER met4 ;
        RECT 8.225 197.975 8.545 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 197.570 8.545 197.890 ;
      LAYER met4 ;
        RECT 8.225 197.570 8.545 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 197.165 8.545 197.485 ;
      LAYER met4 ;
        RECT 8.225 197.165 8.545 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 196.760 8.545 197.080 ;
      LAYER met4 ;
        RECT 8.225 196.760 8.545 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 196.355 8.545 196.675 ;
      LAYER met4 ;
        RECT 8.225 196.355 8.545 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 195.950 8.545 196.270 ;
      LAYER met4 ;
        RECT 8.225 195.950 8.545 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 195.545 8.545 195.865 ;
      LAYER met4 ;
        RECT 8.225 195.545 8.545 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.225 195.140 8.545 195.460 ;
      LAYER met4 ;
        RECT 8.225 195.140 8.545 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 30.210 8.105 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 29.780 8.105 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 29.350 8.105 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 28.920 8.105 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 28.490 8.105 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 28.060 8.105 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 27.630 8.105 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 27.200 8.105 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 26.770 8.105 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 26.340 8.105 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.905 25.910 8.105 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 199.595 8.145 199.915 ;
      LAYER met4 ;
        RECT 7.825 199.595 8.145 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 199.190 8.145 199.510 ;
      LAYER met4 ;
        RECT 7.825 199.190 8.145 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 198.785 8.145 199.105 ;
      LAYER met4 ;
        RECT 7.825 198.785 8.145 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 198.380 8.145 198.700 ;
      LAYER met4 ;
        RECT 7.825 198.380 8.145 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 197.975 8.145 198.295 ;
      LAYER met4 ;
        RECT 7.825 197.975 8.145 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 197.570 8.145 197.890 ;
      LAYER met4 ;
        RECT 7.825 197.570 8.145 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 197.165 8.145 197.485 ;
      LAYER met4 ;
        RECT 7.825 197.165 8.145 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 196.760 8.145 197.080 ;
      LAYER met4 ;
        RECT 7.825 196.760 8.145 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 196.355 8.145 196.675 ;
      LAYER met4 ;
        RECT 7.825 196.355 8.145 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 195.950 8.145 196.270 ;
      LAYER met4 ;
        RECT 7.825 195.950 8.145 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 195.545 8.145 195.865 ;
      LAYER met4 ;
        RECT 7.825 195.545 8.145 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.825 195.140 8.145 195.460 ;
      LAYER met4 ;
        RECT 7.825 195.140 8.145 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 30.210 7.700 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 29.780 7.700 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 29.350 7.700 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 28.920 7.700 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 28.490 7.700 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 28.060 7.700 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 27.630 7.700 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 27.200 7.700 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 26.770 7.700 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 26.340 7.700 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.500 25.910 7.700 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 199.595 7.745 199.915 ;
      LAYER met4 ;
        RECT 7.425 199.595 7.745 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 199.190 7.745 199.510 ;
      LAYER met4 ;
        RECT 7.425 199.190 7.745 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 198.785 7.745 199.105 ;
      LAYER met4 ;
        RECT 7.425 198.785 7.745 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 198.380 7.745 198.700 ;
      LAYER met4 ;
        RECT 7.425 198.380 7.745 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 197.975 7.745 198.295 ;
      LAYER met4 ;
        RECT 7.425 197.975 7.745 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 197.570 7.745 197.890 ;
      LAYER met4 ;
        RECT 7.425 197.570 7.745 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 197.165 7.745 197.485 ;
      LAYER met4 ;
        RECT 7.425 197.165 7.745 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 196.760 7.745 197.080 ;
      LAYER met4 ;
        RECT 7.425 196.760 7.745 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 196.355 7.745 196.675 ;
      LAYER met4 ;
        RECT 7.425 196.355 7.745 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 195.950 7.745 196.270 ;
      LAYER met4 ;
        RECT 7.425 195.950 7.745 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 195.545 7.745 195.865 ;
      LAYER met4 ;
        RECT 7.425 195.545 7.745 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.425 195.140 7.745 195.460 ;
      LAYER met4 ;
        RECT 7.425 195.140 7.745 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 30.210 7.295 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 29.780 7.295 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 29.350 7.295 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 28.920 7.295 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 28.490 7.295 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 28.060 7.295 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 27.630 7.295 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 27.200 7.295 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 26.770 7.295 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 26.340 7.295 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.095 25.910 7.295 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 199.595 7.345 199.915 ;
      LAYER met4 ;
        RECT 7.025 199.595 7.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 199.190 7.345 199.510 ;
      LAYER met4 ;
        RECT 7.025 199.190 7.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 198.785 7.345 199.105 ;
      LAYER met4 ;
        RECT 7.025 198.785 7.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 198.380 7.345 198.700 ;
      LAYER met4 ;
        RECT 7.025 198.380 7.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 197.975 7.345 198.295 ;
      LAYER met4 ;
        RECT 7.025 197.975 7.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 197.570 7.345 197.890 ;
      LAYER met4 ;
        RECT 7.025 197.570 7.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 197.165 7.345 197.485 ;
      LAYER met4 ;
        RECT 7.025 197.165 7.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 196.760 7.345 197.080 ;
      LAYER met4 ;
        RECT 7.025 196.760 7.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 196.355 7.345 196.675 ;
      LAYER met4 ;
        RECT 7.025 196.355 7.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 195.950 7.345 196.270 ;
      LAYER met4 ;
        RECT 7.025 195.950 7.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 195.545 7.345 195.865 ;
      LAYER met4 ;
        RECT 7.025 195.545 7.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.025 195.140 7.345 195.460 ;
      LAYER met4 ;
        RECT 7.025 195.140 7.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 30.210 6.890 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 29.780 6.890 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 29.350 6.890 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 28.920 6.890 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 28.490 6.890 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 28.060 6.890 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 27.630 6.890 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 27.200 6.890 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 26.770 6.890 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 26.340 6.890 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.690 25.910 6.890 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 199.595 6.945 199.915 ;
      LAYER met4 ;
        RECT 6.625 199.595 6.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 199.190 6.945 199.510 ;
      LAYER met4 ;
        RECT 6.625 199.190 6.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 198.785 6.945 199.105 ;
      LAYER met4 ;
        RECT 6.625 198.785 6.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 198.380 6.945 198.700 ;
      LAYER met4 ;
        RECT 6.625 198.380 6.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 197.975 6.945 198.295 ;
      LAYER met4 ;
        RECT 6.625 197.975 6.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 197.570 6.945 197.890 ;
      LAYER met4 ;
        RECT 6.625 197.570 6.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 197.165 6.945 197.485 ;
      LAYER met4 ;
        RECT 6.625 197.165 6.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 196.760 6.945 197.080 ;
      LAYER met4 ;
        RECT 6.625 196.760 6.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 196.355 6.945 196.675 ;
      LAYER met4 ;
        RECT 6.625 196.355 6.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 195.950 6.945 196.270 ;
      LAYER met4 ;
        RECT 6.625 195.950 6.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 195.545 6.945 195.865 ;
      LAYER met4 ;
        RECT 6.625 195.545 6.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.625 195.140 6.945 195.460 ;
      LAYER met4 ;
        RECT 6.625 195.140 6.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 199.595 6.545 199.915 ;
      LAYER met4 ;
        RECT 6.225 199.595 6.545 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 199.190 6.545 199.510 ;
      LAYER met4 ;
        RECT 6.225 199.190 6.545 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 198.785 6.545 199.105 ;
      LAYER met4 ;
        RECT 6.225 198.785 6.545 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 198.380 6.545 198.700 ;
      LAYER met4 ;
        RECT 6.225 198.380 6.545 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 197.975 6.545 198.295 ;
      LAYER met4 ;
        RECT 6.225 197.975 6.545 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 197.570 6.545 197.890 ;
      LAYER met4 ;
        RECT 6.225 197.570 6.545 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 197.165 6.545 197.485 ;
      LAYER met4 ;
        RECT 6.225 197.165 6.545 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 196.760 6.545 197.080 ;
      LAYER met4 ;
        RECT 6.225 196.760 6.545 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 196.355 6.545 196.675 ;
      LAYER met4 ;
        RECT 6.225 196.355 6.545 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 195.950 6.545 196.270 ;
      LAYER met4 ;
        RECT 6.225 195.950 6.545 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 195.545 6.545 195.865 ;
      LAYER met4 ;
        RECT 6.225 195.545 6.545 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 195.140 6.545 195.460 ;
      LAYER met4 ;
        RECT 6.225 195.140 6.545 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 30.210 6.485 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 29.780 6.485 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 29.350 6.485 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 28.920 6.485 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 28.490 6.485 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 28.060 6.485 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 27.630 6.485 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 27.200 6.485 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 26.770 6.485 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 26.340 6.485 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.285 25.910 6.485 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 199.595 6.145 199.915 ;
      LAYER met4 ;
        RECT 5.825 199.595 6.145 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 199.190 6.145 199.510 ;
      LAYER met4 ;
        RECT 5.825 199.190 6.145 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 198.785 6.145 199.105 ;
      LAYER met4 ;
        RECT 5.825 198.785 6.145 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 198.380 6.145 198.700 ;
      LAYER met4 ;
        RECT 5.825 198.380 6.145 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 197.975 6.145 198.295 ;
      LAYER met4 ;
        RECT 5.825 197.975 6.145 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 197.570 6.145 197.890 ;
      LAYER met4 ;
        RECT 5.825 197.570 6.145 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 197.165 6.145 197.485 ;
      LAYER met4 ;
        RECT 5.825 197.165 6.145 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 196.760 6.145 197.080 ;
      LAYER met4 ;
        RECT 5.825 196.760 6.145 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 196.355 6.145 196.675 ;
      LAYER met4 ;
        RECT 5.825 196.355 6.145 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 195.950 6.145 196.270 ;
      LAYER met4 ;
        RECT 5.825 195.950 6.145 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 195.545 6.145 195.865 ;
      LAYER met4 ;
        RECT 5.825 195.545 6.145 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 195.140 6.145 195.460 ;
      LAYER met4 ;
        RECT 5.825 195.140 6.145 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 30.210 6.080 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 29.780 6.080 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 29.350 6.080 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 28.920 6.080 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 28.490 6.080 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 28.060 6.080 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 27.630 6.080 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 27.200 6.080 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 26.770 6.080 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 26.340 6.080 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.880 25.910 6.080 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 199.595 5.745 199.915 ;
      LAYER met4 ;
        RECT 5.425 199.595 5.745 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 199.190 5.745 199.510 ;
      LAYER met4 ;
        RECT 5.425 199.190 5.745 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 198.785 5.745 199.105 ;
      LAYER met4 ;
        RECT 5.425 198.785 5.745 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 198.380 5.745 198.700 ;
      LAYER met4 ;
        RECT 5.425 198.380 5.745 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 197.975 5.745 198.295 ;
      LAYER met4 ;
        RECT 5.425 197.975 5.745 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 197.570 5.745 197.890 ;
      LAYER met4 ;
        RECT 5.425 197.570 5.745 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 197.165 5.745 197.485 ;
      LAYER met4 ;
        RECT 5.425 197.165 5.745 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 196.760 5.745 197.080 ;
      LAYER met4 ;
        RECT 5.425 196.760 5.745 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 196.355 5.745 196.675 ;
      LAYER met4 ;
        RECT 5.425 196.355 5.745 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 195.950 5.745 196.270 ;
      LAYER met4 ;
        RECT 5.425 195.950 5.745 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 195.545 5.745 195.865 ;
      LAYER met4 ;
        RECT 5.425 195.545 5.745 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.425 195.140 5.745 195.460 ;
      LAYER met4 ;
        RECT 5.425 195.140 5.745 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 30.210 5.675 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 29.780 5.675 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 29.350 5.675 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 28.920 5.675 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 28.490 5.675 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 28.060 5.675 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 27.630 5.675 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 27.200 5.675 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 26.770 5.675 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 26.340 5.675 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.475 25.910 5.675 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 199.595 5.345 199.915 ;
      LAYER met4 ;
        RECT 5.025 199.595 5.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 199.190 5.345 199.510 ;
      LAYER met4 ;
        RECT 5.025 199.190 5.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 198.785 5.345 199.105 ;
      LAYER met4 ;
        RECT 5.025 198.785 5.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 198.380 5.345 198.700 ;
      LAYER met4 ;
        RECT 5.025 198.380 5.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 197.975 5.345 198.295 ;
      LAYER met4 ;
        RECT 5.025 197.975 5.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 197.570 5.345 197.890 ;
      LAYER met4 ;
        RECT 5.025 197.570 5.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 197.165 5.345 197.485 ;
      LAYER met4 ;
        RECT 5.025 197.165 5.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 196.760 5.345 197.080 ;
      LAYER met4 ;
        RECT 5.025 196.760 5.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 196.355 5.345 196.675 ;
      LAYER met4 ;
        RECT 5.025 196.355 5.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 195.950 5.345 196.270 ;
      LAYER met4 ;
        RECT 5.025 195.950 5.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 195.545 5.345 195.865 ;
      LAYER met4 ;
        RECT 5.025 195.545 5.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.025 195.140 5.345 195.460 ;
      LAYER met4 ;
        RECT 5.025 195.140 5.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 30.210 5.270 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 29.780 5.270 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 29.350 5.270 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 28.920 5.270 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 28.490 5.270 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 28.060 5.270 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 27.630 5.270 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 27.200 5.270 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 26.770 5.270 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 26.340 5.270 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.070 25.910 5.270 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 199.595 4.945 199.915 ;
      LAYER met4 ;
        RECT 4.625 199.595 4.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 199.190 4.945 199.510 ;
      LAYER met4 ;
        RECT 4.625 199.190 4.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 198.785 4.945 199.105 ;
      LAYER met4 ;
        RECT 4.625 198.785 4.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 198.380 4.945 198.700 ;
      LAYER met4 ;
        RECT 4.625 198.380 4.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 197.975 4.945 198.295 ;
      LAYER met4 ;
        RECT 4.625 197.975 4.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 197.570 4.945 197.890 ;
      LAYER met4 ;
        RECT 4.625 197.570 4.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 197.165 4.945 197.485 ;
      LAYER met4 ;
        RECT 4.625 197.165 4.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 196.760 4.945 197.080 ;
      LAYER met4 ;
        RECT 4.625 196.760 4.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 196.355 4.945 196.675 ;
      LAYER met4 ;
        RECT 4.625 196.355 4.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 195.950 4.945 196.270 ;
      LAYER met4 ;
        RECT 4.625 195.950 4.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 195.545 4.945 195.865 ;
      LAYER met4 ;
        RECT 4.625 195.545 4.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.625 195.140 4.945 195.460 ;
      LAYER met4 ;
        RECT 4.625 195.140 4.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 30.210 4.865 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 29.780 4.865 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 29.350 4.865 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 28.920 4.865 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 28.490 4.865 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 28.060 4.865 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 27.630 4.865 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 27.200 4.865 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 26.770 4.865 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 26.340 4.865 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.665 25.910 4.865 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 199.595 4.545 199.915 ;
      LAYER met4 ;
        RECT 4.225 199.595 4.545 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 199.190 4.545 199.510 ;
      LAYER met4 ;
        RECT 4.225 199.190 4.545 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 198.785 4.545 199.105 ;
      LAYER met4 ;
        RECT 4.225 198.785 4.545 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 198.380 4.545 198.700 ;
      LAYER met4 ;
        RECT 4.225 198.380 4.545 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 197.975 4.545 198.295 ;
      LAYER met4 ;
        RECT 4.225 197.975 4.545 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 197.570 4.545 197.890 ;
      LAYER met4 ;
        RECT 4.225 197.570 4.545 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 197.165 4.545 197.485 ;
      LAYER met4 ;
        RECT 4.225 197.165 4.545 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 196.760 4.545 197.080 ;
      LAYER met4 ;
        RECT 4.225 196.760 4.545 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 196.355 4.545 196.675 ;
      LAYER met4 ;
        RECT 4.225 196.355 4.545 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 195.950 4.545 196.270 ;
      LAYER met4 ;
        RECT 4.225 195.950 4.545 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 195.545 4.545 195.865 ;
      LAYER met4 ;
        RECT 4.225 195.545 4.545 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.225 195.140 4.545 195.460 ;
      LAYER met4 ;
        RECT 4.225 195.140 4.545 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 30.210 4.460 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 29.780 4.460 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 29.350 4.460 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 28.920 4.460 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 28.490 4.460 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 28.060 4.460 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 27.630 4.460 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 27.200 4.460 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 26.770 4.460 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 26.340 4.460 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.260 25.910 4.460 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 199.595 4.145 199.915 ;
      LAYER met4 ;
        RECT 3.825 199.595 4.145 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 199.190 4.145 199.510 ;
      LAYER met4 ;
        RECT 3.825 199.190 4.145 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 198.785 4.145 199.105 ;
      LAYER met4 ;
        RECT 3.825 198.785 4.145 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 198.380 4.145 198.700 ;
      LAYER met4 ;
        RECT 3.825 198.380 4.145 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 197.975 4.145 198.295 ;
      LAYER met4 ;
        RECT 3.825 197.975 4.145 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 197.570 4.145 197.890 ;
      LAYER met4 ;
        RECT 3.825 197.570 4.145 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 197.165 4.145 197.485 ;
      LAYER met4 ;
        RECT 3.825 197.165 4.145 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 196.760 4.145 197.080 ;
      LAYER met4 ;
        RECT 3.825 196.760 4.145 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 196.355 4.145 196.675 ;
      LAYER met4 ;
        RECT 3.825 196.355 4.145 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 195.950 4.145 196.270 ;
      LAYER met4 ;
        RECT 3.825 195.950 4.145 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 195.545 4.145 195.865 ;
      LAYER met4 ;
        RECT 3.825 195.545 4.145 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.825 195.140 4.145 195.460 ;
      LAYER met4 ;
        RECT 3.825 195.140 4.145 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 30.210 4.055 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 29.780 4.055 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 29.350 4.055 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 28.920 4.055 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 28.490 4.055 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 28.060 4.055 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 27.630 4.055 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 27.200 4.055 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 26.770 4.055 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 26.340 4.055 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.855 25.910 4.055 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 199.595 3.745 199.915 ;
      LAYER met4 ;
        RECT 3.425 199.595 3.745 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 199.190 3.745 199.510 ;
      LAYER met4 ;
        RECT 3.425 199.190 3.745 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 198.785 3.745 199.105 ;
      LAYER met4 ;
        RECT 3.425 198.785 3.745 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 198.380 3.745 198.700 ;
      LAYER met4 ;
        RECT 3.425 198.380 3.745 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 197.975 3.745 198.295 ;
      LAYER met4 ;
        RECT 3.425 197.975 3.745 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 197.570 3.745 197.890 ;
      LAYER met4 ;
        RECT 3.425 197.570 3.745 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 197.165 3.745 197.485 ;
      LAYER met4 ;
        RECT 3.425 197.165 3.745 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 196.760 3.745 197.080 ;
      LAYER met4 ;
        RECT 3.425 196.760 3.745 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 196.355 3.745 196.675 ;
      LAYER met4 ;
        RECT 3.425 196.355 3.745 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 195.950 3.745 196.270 ;
      LAYER met4 ;
        RECT 3.425 195.950 3.745 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 195.545 3.745 195.865 ;
      LAYER met4 ;
        RECT 3.425 195.545 3.745 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.425 195.140 3.745 195.460 ;
      LAYER met4 ;
        RECT 3.425 195.140 3.745 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 30.210 3.650 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 29.780 3.650 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 29.350 3.650 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 28.920 3.650 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 28.490 3.650 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 28.060 3.650 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 27.630 3.650 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 27.200 3.650 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 26.770 3.650 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 26.340 3.650 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.450 25.910 3.650 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 199.595 3.345 199.915 ;
      LAYER met4 ;
        RECT 3.025 199.595 3.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 199.190 3.345 199.510 ;
      LAYER met4 ;
        RECT 3.025 199.190 3.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 198.785 3.345 199.105 ;
      LAYER met4 ;
        RECT 3.025 198.785 3.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 198.380 3.345 198.700 ;
      LAYER met4 ;
        RECT 3.025 198.380 3.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 197.975 3.345 198.295 ;
      LAYER met4 ;
        RECT 3.025 197.975 3.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 197.570 3.345 197.890 ;
      LAYER met4 ;
        RECT 3.025 197.570 3.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 197.165 3.345 197.485 ;
      LAYER met4 ;
        RECT 3.025 197.165 3.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 196.760 3.345 197.080 ;
      LAYER met4 ;
        RECT 3.025 196.760 3.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 196.355 3.345 196.675 ;
      LAYER met4 ;
        RECT 3.025 196.355 3.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 195.950 3.345 196.270 ;
      LAYER met4 ;
        RECT 3.025 195.950 3.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 195.545 3.345 195.865 ;
      LAYER met4 ;
        RECT 3.025 195.545 3.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.025 195.140 3.345 195.460 ;
      LAYER met4 ;
        RECT 3.025 195.140 3.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 30.210 3.245 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 29.780 3.245 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 29.350 3.245 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 28.920 3.245 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 28.490 3.245 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 28.060 3.245 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 27.630 3.245 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 27.200 3.245 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 26.770 3.245 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 26.340 3.245 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.045 25.910 3.245 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 199.595 2.945 199.915 ;
      LAYER met4 ;
        RECT 2.625 199.595 2.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 199.190 2.945 199.510 ;
      LAYER met4 ;
        RECT 2.625 199.190 2.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 198.785 2.945 199.105 ;
      LAYER met4 ;
        RECT 2.625 198.785 2.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 198.380 2.945 198.700 ;
      LAYER met4 ;
        RECT 2.625 198.380 2.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 197.975 2.945 198.295 ;
      LAYER met4 ;
        RECT 2.625 197.975 2.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 197.570 2.945 197.890 ;
      LAYER met4 ;
        RECT 2.625 197.570 2.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 197.165 2.945 197.485 ;
      LAYER met4 ;
        RECT 2.625 197.165 2.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 196.760 2.945 197.080 ;
      LAYER met4 ;
        RECT 2.625 196.760 2.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 196.355 2.945 196.675 ;
      LAYER met4 ;
        RECT 2.625 196.355 2.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 195.950 2.945 196.270 ;
      LAYER met4 ;
        RECT 2.625 195.950 2.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 195.545 2.945 195.865 ;
      LAYER met4 ;
        RECT 2.625 195.545 2.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.625 195.140 2.945 195.460 ;
      LAYER met4 ;
        RECT 2.625 195.140 2.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 30.210 2.835 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 29.780 2.835 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 29.350 2.835 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 28.920 2.835 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 28.490 2.835 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 28.060 2.835 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 27.630 2.835 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 27.200 2.835 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 26.770 2.835 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 26.340 2.835 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.635 25.910 2.835 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 199.595 2.545 199.915 ;
      LAYER met4 ;
        RECT 2.225 199.595 2.545 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 199.190 2.545 199.510 ;
      LAYER met4 ;
        RECT 2.225 199.190 2.545 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 198.785 2.545 199.105 ;
      LAYER met4 ;
        RECT 2.225 198.785 2.545 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 198.380 2.545 198.700 ;
      LAYER met4 ;
        RECT 2.225 198.380 2.545 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 197.975 2.545 198.295 ;
      LAYER met4 ;
        RECT 2.225 197.975 2.545 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 197.570 2.545 197.890 ;
      LAYER met4 ;
        RECT 2.225 197.570 2.545 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 197.165 2.545 197.485 ;
      LAYER met4 ;
        RECT 2.225 197.165 2.545 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 196.760 2.545 197.080 ;
      LAYER met4 ;
        RECT 2.225 196.760 2.545 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 196.355 2.545 196.675 ;
      LAYER met4 ;
        RECT 2.225 196.355 2.545 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 195.950 2.545 196.270 ;
      LAYER met4 ;
        RECT 2.225 195.950 2.545 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 195.545 2.545 195.865 ;
      LAYER met4 ;
        RECT 2.225 195.545 2.545 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 195.140 2.545 195.460 ;
      LAYER met4 ;
        RECT 2.225 195.140 2.545 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 30.210 2.425 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 29.780 2.425 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 29.350 2.425 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 28.920 2.425 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 28.490 2.425 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 28.060 2.425 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 27.630 2.425 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 27.200 2.425 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 26.770 2.425 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 26.340 2.425 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.225 25.910 2.425 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 199.595 2.145 199.915 ;
      LAYER met4 ;
        RECT 1.825 199.595 2.145 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 199.190 2.145 199.510 ;
      LAYER met4 ;
        RECT 1.825 199.190 2.145 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 198.785 2.145 199.105 ;
      LAYER met4 ;
        RECT 1.825 198.785 2.145 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 198.380 2.145 198.700 ;
      LAYER met4 ;
        RECT 1.825 198.380 2.145 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 197.975 2.145 198.295 ;
      LAYER met4 ;
        RECT 1.825 197.975 2.145 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 197.570 2.145 197.890 ;
      LAYER met4 ;
        RECT 1.825 197.570 2.145 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 197.165 2.145 197.485 ;
      LAYER met4 ;
        RECT 1.825 197.165 2.145 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 196.760 2.145 197.080 ;
      LAYER met4 ;
        RECT 1.825 196.760 2.145 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 196.355 2.145 196.675 ;
      LAYER met4 ;
        RECT 1.825 196.355 2.145 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 195.950 2.145 196.270 ;
      LAYER met4 ;
        RECT 1.825 195.950 2.145 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 195.545 2.145 195.865 ;
      LAYER met4 ;
        RECT 1.825 195.545 2.145 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.825 195.140 2.145 195.460 ;
      LAYER met4 ;
        RECT 1.825 195.140 2.145 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 30.210 2.015 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 29.780 2.015 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 29.350 2.015 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 28.920 2.015 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 28.490 2.015 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 28.060 2.015 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 27.630 2.015 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 27.200 2.015 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 26.770 2.015 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 26.340 2.015 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.815 25.910 2.015 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 199.595 1.745 199.915 ;
      LAYER met4 ;
        RECT 1.425 199.595 1.745 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 199.190 1.745 199.510 ;
      LAYER met4 ;
        RECT 1.425 199.190 1.745 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 198.785 1.745 199.105 ;
      LAYER met4 ;
        RECT 1.425 198.785 1.745 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 198.380 1.745 198.700 ;
      LAYER met4 ;
        RECT 1.425 198.380 1.745 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 197.975 1.745 198.295 ;
      LAYER met4 ;
        RECT 1.425 197.975 1.745 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 197.570 1.745 197.890 ;
      LAYER met4 ;
        RECT 1.425 197.570 1.745 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 197.165 1.745 197.485 ;
      LAYER met4 ;
        RECT 1.425 197.165 1.745 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 196.760 1.745 197.080 ;
      LAYER met4 ;
        RECT 1.425 196.760 1.745 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 196.355 1.745 196.675 ;
      LAYER met4 ;
        RECT 1.425 196.355 1.745 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 195.950 1.745 196.270 ;
      LAYER met4 ;
        RECT 1.425 195.950 1.745 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 195.545 1.745 195.865 ;
      LAYER met4 ;
        RECT 1.425 195.545 1.745 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.425 195.140 1.745 195.460 ;
      LAYER met4 ;
        RECT 1.425 195.140 1.745 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 30.210 1.605 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 29.780 1.605 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 29.350 1.605 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 28.920 1.605 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 28.490 1.605 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 28.060 1.605 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 27.630 1.605 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 27.200 1.605 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 26.770 1.605 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 26.340 1.605 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.405 25.910 1.605 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 199.595 1.345 199.915 ;
      LAYER met4 ;
        RECT 1.270 199.595 1.345 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 199.190 1.345 199.510 ;
      LAYER met4 ;
        RECT 1.270 199.190 1.345 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 198.785 1.345 199.105 ;
      LAYER met4 ;
        RECT 1.270 198.785 1.345 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 198.380 1.345 198.700 ;
      LAYER met4 ;
        RECT 1.270 198.380 1.345 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 197.975 1.345 198.295 ;
      LAYER met4 ;
        RECT 1.270 197.975 1.345 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 197.570 1.345 197.890 ;
      LAYER met4 ;
        RECT 1.270 197.570 1.345 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 197.165 1.345 197.485 ;
      LAYER met4 ;
        RECT 1.270 197.165 1.345 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 196.760 1.345 197.080 ;
      LAYER met4 ;
        RECT 1.270 196.760 1.345 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 196.355 1.345 196.675 ;
      LAYER met4 ;
        RECT 1.270 196.355 1.345 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 195.950 1.345 196.270 ;
      LAYER met4 ;
        RECT 1.270 195.950 1.345 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 195.545 1.345 195.865 ;
      LAYER met4 ;
        RECT 1.270 195.545 1.345 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.025 195.140 1.345 195.460 ;
      LAYER met4 ;
        RECT 1.270 195.140 1.345 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 30.210 1.195 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 29.780 1.195 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 29.350 1.195 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 28.920 1.195 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 28.490 1.195 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 28.060 1.195 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 27.630 1.195 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 27.200 1.195 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 26.770 1.195 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 26.340 1.195 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.995 25.910 1.195 26.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 199.595 0.945 199.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 199.190 0.945 199.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 198.785 0.945 199.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 198.380 0.945 198.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 197.975 0.945 198.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 197.570 0.945 197.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 197.165 0.945 197.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 196.760 0.945 197.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 196.355 0.945 196.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 195.950 0.945 196.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 195.545 0.945 195.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.625 195.140 0.945 195.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 30.210 0.785 30.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 29.780 0.785 29.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 29.350 0.785 29.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 28.920 0.785 29.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 28.490 0.785 28.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 28.060 0.785 28.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 27.630 0.785 27.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 27.200 0.785 27.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 26.770 0.785 26.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 26.340 0.785 26.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.585 25.910 0.785 26.110 ;
    END
  END VSSIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
  END VSWITCH
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 62.350 74.260 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 61.940 74.260 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 61.530 74.260 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 61.120 74.260 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 60.710 74.260 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 60.300 74.260 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 59.890 74.260 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 59.480 74.260 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 59.070 74.260 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 58.660 74.260 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.940 58.250 74.260 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 62.350 73.855 62.670 ;
      LAYER met4 ;
        RECT 73.535 62.350 73.730 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 61.940 73.855 62.260 ;
      LAYER met4 ;
        RECT 73.535 61.940 73.730 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 61.530 73.855 61.850 ;
      LAYER met4 ;
        RECT 73.535 61.530 73.730 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 61.120 73.855 61.440 ;
      LAYER met4 ;
        RECT 73.535 61.120 73.730 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 60.710 73.855 61.030 ;
      LAYER met4 ;
        RECT 73.535 60.710 73.730 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 60.300 73.855 60.620 ;
      LAYER met4 ;
        RECT 73.535 60.300 73.730 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 59.890 73.855 60.210 ;
      LAYER met4 ;
        RECT 73.535 59.890 73.730 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 59.480 73.855 59.800 ;
      LAYER met4 ;
        RECT 73.535 59.480 73.730 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 59.070 73.855 59.390 ;
      LAYER met4 ;
        RECT 73.535 59.070 73.730 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 58.660 73.855 58.980 ;
      LAYER met4 ;
        RECT 73.535 58.660 73.730 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.535 58.250 73.855 58.570 ;
      LAYER met4 ;
        RECT 73.535 58.250 73.730 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 62.350 73.450 62.670 ;
      LAYER met4 ;
        RECT 73.130 62.350 73.450 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 61.940 73.450 62.260 ;
      LAYER met4 ;
        RECT 73.130 61.940 73.450 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 61.530 73.450 61.850 ;
      LAYER met4 ;
        RECT 73.130 61.530 73.450 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 61.120 73.450 61.440 ;
      LAYER met4 ;
        RECT 73.130 61.120 73.450 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 60.710 73.450 61.030 ;
      LAYER met4 ;
        RECT 73.130 60.710 73.450 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 60.300 73.450 60.620 ;
      LAYER met4 ;
        RECT 73.130 60.300 73.450 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 59.890 73.450 60.210 ;
      LAYER met4 ;
        RECT 73.130 59.890 73.450 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 59.480 73.450 59.800 ;
      LAYER met4 ;
        RECT 73.130 59.480 73.450 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 59.070 73.450 59.390 ;
      LAYER met4 ;
        RECT 73.130 59.070 73.450 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 58.660 73.450 58.980 ;
      LAYER met4 ;
        RECT 73.130 58.660 73.450 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.130 58.250 73.450 58.570 ;
      LAYER met4 ;
        RECT 73.130 58.250 73.450 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 62.350 73.045 62.670 ;
      LAYER met4 ;
        RECT 72.725 62.350 73.045 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 61.940 73.045 62.260 ;
      LAYER met4 ;
        RECT 72.725 61.940 73.045 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 61.530 73.045 61.850 ;
      LAYER met4 ;
        RECT 72.725 61.530 73.045 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 61.120 73.045 61.440 ;
      LAYER met4 ;
        RECT 72.725 61.120 73.045 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 60.710 73.045 61.030 ;
      LAYER met4 ;
        RECT 72.725 60.710 73.045 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 60.300 73.045 60.620 ;
      LAYER met4 ;
        RECT 72.725 60.300 73.045 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 59.890 73.045 60.210 ;
      LAYER met4 ;
        RECT 72.725 59.890 73.045 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 59.480 73.045 59.800 ;
      LAYER met4 ;
        RECT 72.725 59.480 73.045 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 59.070 73.045 59.390 ;
      LAYER met4 ;
        RECT 72.725 59.070 73.045 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 58.660 73.045 58.980 ;
      LAYER met4 ;
        RECT 72.725 58.660 73.045 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.725 58.250 73.045 58.570 ;
      LAYER met4 ;
        RECT 72.725 58.250 73.045 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 62.350 72.640 62.670 ;
      LAYER met4 ;
        RECT 72.320 62.350 72.640 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 61.940 72.640 62.260 ;
      LAYER met4 ;
        RECT 72.320 61.940 72.640 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 61.530 72.640 61.850 ;
      LAYER met4 ;
        RECT 72.320 61.530 72.640 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 61.120 72.640 61.440 ;
      LAYER met4 ;
        RECT 72.320 61.120 72.640 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 60.710 72.640 61.030 ;
      LAYER met4 ;
        RECT 72.320 60.710 72.640 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 60.300 72.640 60.620 ;
      LAYER met4 ;
        RECT 72.320 60.300 72.640 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 59.890 72.640 60.210 ;
      LAYER met4 ;
        RECT 72.320 59.890 72.640 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 59.480 72.640 59.800 ;
      LAYER met4 ;
        RECT 72.320 59.480 72.640 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 59.070 72.640 59.390 ;
      LAYER met4 ;
        RECT 72.320 59.070 72.640 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 58.660 72.640 58.980 ;
      LAYER met4 ;
        RECT 72.320 58.660 72.640 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.320 58.250 72.640 58.570 ;
      LAYER met4 ;
        RECT 72.320 58.250 72.640 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 62.350 72.235 62.670 ;
      LAYER met4 ;
        RECT 71.915 62.350 72.235 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 61.940 72.235 62.260 ;
      LAYER met4 ;
        RECT 71.915 61.940 72.235 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 61.530 72.235 61.850 ;
      LAYER met4 ;
        RECT 71.915 61.530 72.235 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 61.120 72.235 61.440 ;
      LAYER met4 ;
        RECT 71.915 61.120 72.235 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 60.710 72.235 61.030 ;
      LAYER met4 ;
        RECT 71.915 60.710 72.235 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 60.300 72.235 60.620 ;
      LAYER met4 ;
        RECT 71.915 60.300 72.235 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 59.890 72.235 60.210 ;
      LAYER met4 ;
        RECT 71.915 59.890 72.235 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 59.480 72.235 59.800 ;
      LAYER met4 ;
        RECT 71.915 59.480 72.235 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 59.070 72.235 59.390 ;
      LAYER met4 ;
        RECT 71.915 59.070 72.235 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 58.660 72.235 58.980 ;
      LAYER met4 ;
        RECT 71.915 58.660 72.235 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 58.250 72.235 58.570 ;
      LAYER met4 ;
        RECT 71.915 58.250 72.235 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 62.350 71.830 62.670 ;
      LAYER met4 ;
        RECT 71.510 62.350 71.830 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 61.940 71.830 62.260 ;
      LAYER met4 ;
        RECT 71.510 61.940 71.830 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 61.530 71.830 61.850 ;
      LAYER met4 ;
        RECT 71.510 61.530 71.830 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 61.120 71.830 61.440 ;
      LAYER met4 ;
        RECT 71.510 61.120 71.830 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 60.710 71.830 61.030 ;
      LAYER met4 ;
        RECT 71.510 60.710 71.830 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 60.300 71.830 60.620 ;
      LAYER met4 ;
        RECT 71.510 60.300 71.830 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 59.890 71.830 60.210 ;
      LAYER met4 ;
        RECT 71.510 59.890 71.830 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 59.480 71.830 59.800 ;
      LAYER met4 ;
        RECT 71.510 59.480 71.830 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 59.070 71.830 59.390 ;
      LAYER met4 ;
        RECT 71.510 59.070 71.830 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 58.660 71.830 58.980 ;
      LAYER met4 ;
        RECT 71.510 58.660 71.830 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.510 58.250 71.830 58.570 ;
      LAYER met4 ;
        RECT 71.510 58.250 71.830 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 62.350 71.425 62.670 ;
      LAYER met4 ;
        RECT 71.105 62.350 71.425 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 61.940 71.425 62.260 ;
      LAYER met4 ;
        RECT 71.105 61.940 71.425 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 61.530 71.425 61.850 ;
      LAYER met4 ;
        RECT 71.105 61.530 71.425 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 61.120 71.425 61.440 ;
      LAYER met4 ;
        RECT 71.105 61.120 71.425 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 60.710 71.425 61.030 ;
      LAYER met4 ;
        RECT 71.105 60.710 71.425 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 60.300 71.425 60.620 ;
      LAYER met4 ;
        RECT 71.105 60.300 71.425 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 59.890 71.425 60.210 ;
      LAYER met4 ;
        RECT 71.105 59.890 71.425 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 59.480 71.425 59.800 ;
      LAYER met4 ;
        RECT 71.105 59.480 71.425 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 59.070 71.425 59.390 ;
      LAYER met4 ;
        RECT 71.105 59.070 71.425 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 58.660 71.425 58.980 ;
      LAYER met4 ;
        RECT 71.105 58.660 71.425 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.105 58.250 71.425 58.570 ;
      LAYER met4 ;
        RECT 71.105 58.250 71.425 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 62.350 71.020 62.670 ;
      LAYER met4 ;
        RECT 70.700 62.350 71.020 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 61.940 71.020 62.260 ;
      LAYER met4 ;
        RECT 70.700 61.940 71.020 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 61.530 71.020 61.850 ;
      LAYER met4 ;
        RECT 70.700 61.530 71.020 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 61.120 71.020 61.440 ;
      LAYER met4 ;
        RECT 70.700 61.120 71.020 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 60.710 71.020 61.030 ;
      LAYER met4 ;
        RECT 70.700 60.710 71.020 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 60.300 71.020 60.620 ;
      LAYER met4 ;
        RECT 70.700 60.300 71.020 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 59.890 71.020 60.210 ;
      LAYER met4 ;
        RECT 70.700 59.890 71.020 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 59.480 71.020 59.800 ;
      LAYER met4 ;
        RECT 70.700 59.480 71.020 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 59.070 71.020 59.390 ;
      LAYER met4 ;
        RECT 70.700 59.070 71.020 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 58.660 71.020 58.980 ;
      LAYER met4 ;
        RECT 70.700 58.660 71.020 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.700 58.250 71.020 58.570 ;
      LAYER met4 ;
        RECT 70.700 58.250 71.020 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 62.350 70.615 62.670 ;
      LAYER met4 ;
        RECT 70.295 62.350 70.615 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 61.940 70.615 62.260 ;
      LAYER met4 ;
        RECT 70.295 61.940 70.615 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 61.530 70.615 61.850 ;
      LAYER met4 ;
        RECT 70.295 61.530 70.615 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 61.120 70.615 61.440 ;
      LAYER met4 ;
        RECT 70.295 61.120 70.615 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 60.710 70.615 61.030 ;
      LAYER met4 ;
        RECT 70.295 60.710 70.615 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 60.300 70.615 60.620 ;
      LAYER met4 ;
        RECT 70.295 60.300 70.615 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 59.890 70.615 60.210 ;
      LAYER met4 ;
        RECT 70.295 59.890 70.615 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 59.480 70.615 59.800 ;
      LAYER met4 ;
        RECT 70.295 59.480 70.615 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 59.070 70.615 59.390 ;
      LAYER met4 ;
        RECT 70.295 59.070 70.615 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 58.660 70.615 58.980 ;
      LAYER met4 ;
        RECT 70.295 58.660 70.615 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.295 58.250 70.615 58.570 ;
      LAYER met4 ;
        RECT 70.295 58.250 70.615 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 62.350 70.210 62.670 ;
      LAYER met4 ;
        RECT 69.890 62.350 70.210 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 61.940 70.210 62.260 ;
      LAYER met4 ;
        RECT 69.890 61.940 70.210 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 61.530 70.210 61.850 ;
      LAYER met4 ;
        RECT 69.890 61.530 70.210 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 61.120 70.210 61.440 ;
      LAYER met4 ;
        RECT 69.890 61.120 70.210 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 60.710 70.210 61.030 ;
      LAYER met4 ;
        RECT 69.890 60.710 70.210 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 60.300 70.210 60.620 ;
      LAYER met4 ;
        RECT 69.890 60.300 70.210 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 59.890 70.210 60.210 ;
      LAYER met4 ;
        RECT 69.890 59.890 70.210 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 59.480 70.210 59.800 ;
      LAYER met4 ;
        RECT 69.890 59.480 70.210 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 59.070 70.210 59.390 ;
      LAYER met4 ;
        RECT 69.890 59.070 70.210 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 58.660 70.210 58.980 ;
      LAYER met4 ;
        RECT 69.890 58.660 70.210 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.890 58.250 70.210 58.570 ;
      LAYER met4 ;
        RECT 69.890 58.250 70.210 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 62.350 69.805 62.670 ;
      LAYER met4 ;
        RECT 69.485 62.350 69.805 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 61.940 69.805 62.260 ;
      LAYER met4 ;
        RECT 69.485 61.940 69.805 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 61.530 69.805 61.850 ;
      LAYER met4 ;
        RECT 69.485 61.530 69.805 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 61.120 69.805 61.440 ;
      LAYER met4 ;
        RECT 69.485 61.120 69.805 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 60.710 69.805 61.030 ;
      LAYER met4 ;
        RECT 69.485 60.710 69.805 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 60.300 69.805 60.620 ;
      LAYER met4 ;
        RECT 69.485 60.300 69.805 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 59.890 69.805 60.210 ;
      LAYER met4 ;
        RECT 69.485 59.890 69.805 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 59.480 69.805 59.800 ;
      LAYER met4 ;
        RECT 69.485 59.480 69.805 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 59.070 69.805 59.390 ;
      LAYER met4 ;
        RECT 69.485 59.070 69.805 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 58.660 69.805 58.980 ;
      LAYER met4 ;
        RECT 69.485 58.660 69.805 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.485 58.250 69.805 58.570 ;
      LAYER met4 ;
        RECT 69.485 58.250 69.805 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 62.350 69.400 62.670 ;
      LAYER met4 ;
        RECT 69.080 62.350 69.400 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 61.940 69.400 62.260 ;
      LAYER met4 ;
        RECT 69.080 61.940 69.400 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 61.530 69.400 61.850 ;
      LAYER met4 ;
        RECT 69.080 61.530 69.400 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 61.120 69.400 61.440 ;
      LAYER met4 ;
        RECT 69.080 61.120 69.400 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 60.710 69.400 61.030 ;
      LAYER met4 ;
        RECT 69.080 60.710 69.400 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 60.300 69.400 60.620 ;
      LAYER met4 ;
        RECT 69.080 60.300 69.400 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 59.890 69.400 60.210 ;
      LAYER met4 ;
        RECT 69.080 59.890 69.400 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 59.480 69.400 59.800 ;
      LAYER met4 ;
        RECT 69.080 59.480 69.400 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 59.070 69.400 59.390 ;
      LAYER met4 ;
        RECT 69.080 59.070 69.400 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 58.660 69.400 58.980 ;
      LAYER met4 ;
        RECT 69.080 58.660 69.400 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.080 58.250 69.400 58.570 ;
      LAYER met4 ;
        RECT 69.080 58.250 69.400 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 62.350 68.995 62.670 ;
      LAYER met4 ;
        RECT 68.675 62.350 68.995 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 61.940 68.995 62.260 ;
      LAYER met4 ;
        RECT 68.675 61.940 68.995 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 61.530 68.995 61.850 ;
      LAYER met4 ;
        RECT 68.675 61.530 68.995 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 61.120 68.995 61.440 ;
      LAYER met4 ;
        RECT 68.675 61.120 68.995 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 60.710 68.995 61.030 ;
      LAYER met4 ;
        RECT 68.675 60.710 68.995 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 60.300 68.995 60.620 ;
      LAYER met4 ;
        RECT 68.675 60.300 68.995 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 59.890 68.995 60.210 ;
      LAYER met4 ;
        RECT 68.675 59.890 68.995 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 59.480 68.995 59.800 ;
      LAYER met4 ;
        RECT 68.675 59.480 68.995 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 59.070 68.995 59.390 ;
      LAYER met4 ;
        RECT 68.675 59.070 68.995 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 58.660 68.995 58.980 ;
      LAYER met4 ;
        RECT 68.675 58.660 68.995 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.675 58.250 68.995 58.570 ;
      LAYER met4 ;
        RECT 68.675 58.250 68.995 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 62.350 68.590 62.670 ;
      LAYER met4 ;
        RECT 68.270 62.350 68.590 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 61.940 68.590 62.260 ;
      LAYER met4 ;
        RECT 68.270 61.940 68.590 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 61.530 68.590 61.850 ;
      LAYER met4 ;
        RECT 68.270 61.530 68.590 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 61.120 68.590 61.440 ;
      LAYER met4 ;
        RECT 68.270 61.120 68.590 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 60.710 68.590 61.030 ;
      LAYER met4 ;
        RECT 68.270 60.710 68.590 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 60.300 68.590 60.620 ;
      LAYER met4 ;
        RECT 68.270 60.300 68.590 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 59.890 68.590 60.210 ;
      LAYER met4 ;
        RECT 68.270 59.890 68.590 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 59.480 68.590 59.800 ;
      LAYER met4 ;
        RECT 68.270 59.480 68.590 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 59.070 68.590 59.390 ;
      LAYER met4 ;
        RECT 68.270 59.070 68.590 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 58.660 68.590 58.980 ;
      LAYER met4 ;
        RECT 68.270 58.660 68.590 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.270 58.250 68.590 58.570 ;
      LAYER met4 ;
        RECT 68.270 58.250 68.590 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 62.350 68.185 62.670 ;
      LAYER met4 ;
        RECT 67.865 62.350 68.185 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 61.940 68.185 62.260 ;
      LAYER met4 ;
        RECT 67.865 61.940 68.185 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 61.530 68.185 61.850 ;
      LAYER met4 ;
        RECT 67.865 61.530 68.185 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 61.120 68.185 61.440 ;
      LAYER met4 ;
        RECT 67.865 61.120 68.185 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 60.710 68.185 61.030 ;
      LAYER met4 ;
        RECT 67.865 60.710 68.185 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 60.300 68.185 60.620 ;
      LAYER met4 ;
        RECT 67.865 60.300 68.185 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 59.890 68.185 60.210 ;
      LAYER met4 ;
        RECT 67.865 59.890 68.185 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 59.480 68.185 59.800 ;
      LAYER met4 ;
        RECT 67.865 59.480 68.185 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 59.070 68.185 59.390 ;
      LAYER met4 ;
        RECT 67.865 59.070 68.185 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 58.660 68.185 58.980 ;
      LAYER met4 ;
        RECT 67.865 58.660 68.185 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.865 58.250 68.185 58.570 ;
      LAYER met4 ;
        RECT 67.865 58.250 68.185 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 62.350 67.780 62.670 ;
      LAYER met4 ;
        RECT 67.460 62.350 67.780 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 61.940 67.780 62.260 ;
      LAYER met4 ;
        RECT 67.460 61.940 67.780 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 61.530 67.780 61.850 ;
      LAYER met4 ;
        RECT 67.460 61.530 67.780 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 61.120 67.780 61.440 ;
      LAYER met4 ;
        RECT 67.460 61.120 67.780 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 60.710 67.780 61.030 ;
      LAYER met4 ;
        RECT 67.460 60.710 67.780 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 60.300 67.780 60.620 ;
      LAYER met4 ;
        RECT 67.460 60.300 67.780 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 59.890 67.780 60.210 ;
      LAYER met4 ;
        RECT 67.460 59.890 67.780 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 59.480 67.780 59.800 ;
      LAYER met4 ;
        RECT 67.460 59.480 67.780 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 59.070 67.780 59.390 ;
      LAYER met4 ;
        RECT 67.460 59.070 67.780 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 58.660 67.780 58.980 ;
      LAYER met4 ;
        RECT 67.460 58.660 67.780 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.460 58.250 67.780 58.570 ;
      LAYER met4 ;
        RECT 67.460 58.250 67.780 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 62.350 67.375 62.670 ;
      LAYER met4 ;
        RECT 67.055 62.350 67.375 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 61.940 67.375 62.260 ;
      LAYER met4 ;
        RECT 67.055 61.940 67.375 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 61.530 67.375 61.850 ;
      LAYER met4 ;
        RECT 67.055 61.530 67.375 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 61.120 67.375 61.440 ;
      LAYER met4 ;
        RECT 67.055 61.120 67.375 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 60.710 67.375 61.030 ;
      LAYER met4 ;
        RECT 67.055 60.710 67.375 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 60.300 67.375 60.620 ;
      LAYER met4 ;
        RECT 67.055 60.300 67.375 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 59.890 67.375 60.210 ;
      LAYER met4 ;
        RECT 67.055 59.890 67.375 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 59.480 67.375 59.800 ;
      LAYER met4 ;
        RECT 67.055 59.480 67.375 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 59.070 67.375 59.390 ;
      LAYER met4 ;
        RECT 67.055 59.070 67.375 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 58.660 67.375 58.980 ;
      LAYER met4 ;
        RECT 67.055 58.660 67.375 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.055 58.250 67.375 58.570 ;
      LAYER met4 ;
        RECT 67.055 58.250 67.375 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 62.350 66.970 62.670 ;
      LAYER met4 ;
        RECT 66.650 62.350 66.970 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 61.940 66.970 62.260 ;
      LAYER met4 ;
        RECT 66.650 61.940 66.970 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 61.530 66.970 61.850 ;
      LAYER met4 ;
        RECT 66.650 61.530 66.970 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 61.120 66.970 61.440 ;
      LAYER met4 ;
        RECT 66.650 61.120 66.970 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 60.710 66.970 61.030 ;
      LAYER met4 ;
        RECT 66.650 60.710 66.970 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 60.300 66.970 60.620 ;
      LAYER met4 ;
        RECT 66.650 60.300 66.970 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 59.890 66.970 60.210 ;
      LAYER met4 ;
        RECT 66.650 59.890 66.970 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 59.480 66.970 59.800 ;
      LAYER met4 ;
        RECT 66.650 59.480 66.970 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 59.070 66.970 59.390 ;
      LAYER met4 ;
        RECT 66.650 59.070 66.970 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 58.660 66.970 58.980 ;
      LAYER met4 ;
        RECT 66.650 58.660 66.970 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 58.250 66.970 58.570 ;
      LAYER met4 ;
        RECT 66.650 58.250 66.970 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 62.350 66.565 62.670 ;
      LAYER met4 ;
        RECT 66.245 62.350 66.565 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 61.940 66.565 62.260 ;
      LAYER met4 ;
        RECT 66.245 61.940 66.565 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 61.530 66.565 61.850 ;
      LAYER met4 ;
        RECT 66.245 61.530 66.565 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 61.120 66.565 61.440 ;
      LAYER met4 ;
        RECT 66.245 61.120 66.565 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 60.710 66.565 61.030 ;
      LAYER met4 ;
        RECT 66.245 60.710 66.565 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 60.300 66.565 60.620 ;
      LAYER met4 ;
        RECT 66.245 60.300 66.565 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 59.890 66.565 60.210 ;
      LAYER met4 ;
        RECT 66.245 59.890 66.565 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 59.480 66.565 59.800 ;
      LAYER met4 ;
        RECT 66.245 59.480 66.565 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 59.070 66.565 59.390 ;
      LAYER met4 ;
        RECT 66.245 59.070 66.565 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 58.660 66.565 58.980 ;
      LAYER met4 ;
        RECT 66.245 58.660 66.565 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.245 58.250 66.565 58.570 ;
      LAYER met4 ;
        RECT 66.245 58.250 66.565 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 62.350 66.160 62.670 ;
      LAYER met4 ;
        RECT 65.840 62.350 66.160 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 61.940 66.160 62.260 ;
      LAYER met4 ;
        RECT 65.840 61.940 66.160 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 61.530 66.160 61.850 ;
      LAYER met4 ;
        RECT 65.840 61.530 66.160 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 61.120 66.160 61.440 ;
      LAYER met4 ;
        RECT 65.840 61.120 66.160 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 60.710 66.160 61.030 ;
      LAYER met4 ;
        RECT 65.840 60.710 66.160 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 60.300 66.160 60.620 ;
      LAYER met4 ;
        RECT 65.840 60.300 66.160 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 59.890 66.160 60.210 ;
      LAYER met4 ;
        RECT 65.840 59.890 66.160 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 59.480 66.160 59.800 ;
      LAYER met4 ;
        RECT 65.840 59.480 66.160 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 59.070 66.160 59.390 ;
      LAYER met4 ;
        RECT 65.840 59.070 66.160 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 58.660 66.160 58.980 ;
      LAYER met4 ;
        RECT 65.840 58.660 66.160 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.840 58.250 66.160 58.570 ;
      LAYER met4 ;
        RECT 65.840 58.250 66.160 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 62.350 65.755 62.670 ;
      LAYER met4 ;
        RECT 65.435 62.350 65.755 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 61.940 65.755 62.260 ;
      LAYER met4 ;
        RECT 65.435 61.940 65.755 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 61.530 65.755 61.850 ;
      LAYER met4 ;
        RECT 65.435 61.530 65.755 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 61.120 65.755 61.440 ;
      LAYER met4 ;
        RECT 65.435 61.120 65.755 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 60.710 65.755 61.030 ;
      LAYER met4 ;
        RECT 65.435 60.710 65.755 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 60.300 65.755 60.620 ;
      LAYER met4 ;
        RECT 65.435 60.300 65.755 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 59.890 65.755 60.210 ;
      LAYER met4 ;
        RECT 65.435 59.890 65.755 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 59.480 65.755 59.800 ;
      LAYER met4 ;
        RECT 65.435 59.480 65.755 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 59.070 65.755 59.390 ;
      LAYER met4 ;
        RECT 65.435 59.070 65.755 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 58.660 65.755 58.980 ;
      LAYER met4 ;
        RECT 65.435 58.660 65.755 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.435 58.250 65.755 58.570 ;
      LAYER met4 ;
        RECT 65.435 58.250 65.755 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 62.350 65.350 62.670 ;
      LAYER met4 ;
        RECT 65.030 62.350 65.350 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 61.940 65.350 62.260 ;
      LAYER met4 ;
        RECT 65.030 61.940 65.350 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 61.530 65.350 61.850 ;
      LAYER met4 ;
        RECT 65.030 61.530 65.350 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 61.120 65.350 61.440 ;
      LAYER met4 ;
        RECT 65.030 61.120 65.350 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 60.710 65.350 61.030 ;
      LAYER met4 ;
        RECT 65.030 60.710 65.350 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 60.300 65.350 60.620 ;
      LAYER met4 ;
        RECT 65.030 60.300 65.350 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 59.890 65.350 60.210 ;
      LAYER met4 ;
        RECT 65.030 59.890 65.350 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 59.480 65.350 59.800 ;
      LAYER met4 ;
        RECT 65.030 59.480 65.350 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 59.070 65.350 59.390 ;
      LAYER met4 ;
        RECT 65.030 59.070 65.350 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 58.660 65.350 58.980 ;
      LAYER met4 ;
        RECT 65.030 58.660 65.350 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.030 58.250 65.350 58.570 ;
      LAYER met4 ;
        RECT 65.030 58.250 65.350 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 62.350 64.945 62.670 ;
      LAYER met4 ;
        RECT 64.625 62.350 64.945 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 61.940 64.945 62.260 ;
      LAYER met4 ;
        RECT 64.625 61.940 64.945 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 61.530 64.945 61.850 ;
      LAYER met4 ;
        RECT 64.625 61.530 64.945 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 61.120 64.945 61.440 ;
      LAYER met4 ;
        RECT 64.625 61.120 64.945 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 60.710 64.945 61.030 ;
      LAYER met4 ;
        RECT 64.625 60.710 64.945 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 60.300 64.945 60.620 ;
      LAYER met4 ;
        RECT 64.625 60.300 64.945 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 59.890 64.945 60.210 ;
      LAYER met4 ;
        RECT 64.625 59.890 64.945 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 59.480 64.945 59.800 ;
      LAYER met4 ;
        RECT 64.625 59.480 64.945 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 59.070 64.945 59.390 ;
      LAYER met4 ;
        RECT 64.625 59.070 64.945 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 58.660 64.945 58.980 ;
      LAYER met4 ;
        RECT 64.625 58.660 64.945 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.625 58.250 64.945 58.570 ;
      LAYER met4 ;
        RECT 64.625 58.250 64.945 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 62.350 64.540 62.670 ;
      LAYER met4 ;
        RECT 64.220 62.350 64.540 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 61.940 64.540 62.260 ;
      LAYER met4 ;
        RECT 64.220 61.940 64.540 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 61.530 64.540 61.850 ;
      LAYER met4 ;
        RECT 64.220 61.530 64.540 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 61.120 64.540 61.440 ;
      LAYER met4 ;
        RECT 64.220 61.120 64.540 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 60.710 64.540 61.030 ;
      LAYER met4 ;
        RECT 64.220 60.710 64.540 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 60.300 64.540 60.620 ;
      LAYER met4 ;
        RECT 64.220 60.300 64.540 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 59.890 64.540 60.210 ;
      LAYER met4 ;
        RECT 64.220 59.890 64.540 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 59.480 64.540 59.800 ;
      LAYER met4 ;
        RECT 64.220 59.480 64.540 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 59.070 64.540 59.390 ;
      LAYER met4 ;
        RECT 64.220 59.070 64.540 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 58.660 64.540 58.980 ;
      LAYER met4 ;
        RECT 64.220 58.660 64.540 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.220 58.250 64.540 58.570 ;
      LAYER met4 ;
        RECT 64.220 58.250 64.540 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 62.350 64.135 62.670 ;
      LAYER met4 ;
        RECT 63.815 62.350 64.135 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 61.940 64.135 62.260 ;
      LAYER met4 ;
        RECT 63.815 61.940 64.135 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 61.530 64.135 61.850 ;
      LAYER met4 ;
        RECT 63.815 61.530 64.135 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 61.120 64.135 61.440 ;
      LAYER met4 ;
        RECT 63.815 61.120 64.135 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 60.710 64.135 61.030 ;
      LAYER met4 ;
        RECT 63.815 60.710 64.135 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 60.300 64.135 60.620 ;
      LAYER met4 ;
        RECT 63.815 60.300 64.135 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 59.890 64.135 60.210 ;
      LAYER met4 ;
        RECT 63.815 59.890 64.135 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 59.480 64.135 59.800 ;
      LAYER met4 ;
        RECT 63.815 59.480 64.135 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 59.070 64.135 59.390 ;
      LAYER met4 ;
        RECT 63.815 59.070 64.135 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 58.660 64.135 58.980 ;
      LAYER met4 ;
        RECT 63.815 58.660 64.135 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.815 58.250 64.135 58.570 ;
      LAYER met4 ;
        RECT 63.815 58.250 64.135 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 62.350 63.730 62.670 ;
      LAYER met4 ;
        RECT 63.410 62.350 63.730 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 61.940 63.730 62.260 ;
      LAYER met4 ;
        RECT 63.410 61.940 63.730 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 61.530 63.730 61.850 ;
      LAYER met4 ;
        RECT 63.410 61.530 63.730 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 61.120 63.730 61.440 ;
      LAYER met4 ;
        RECT 63.410 61.120 63.730 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 60.710 63.730 61.030 ;
      LAYER met4 ;
        RECT 63.410 60.710 63.730 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 60.300 63.730 60.620 ;
      LAYER met4 ;
        RECT 63.410 60.300 63.730 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 59.890 63.730 60.210 ;
      LAYER met4 ;
        RECT 63.410 59.890 63.730 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 59.480 63.730 59.800 ;
      LAYER met4 ;
        RECT 63.410 59.480 63.730 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 59.070 63.730 59.390 ;
      LAYER met4 ;
        RECT 63.410 59.070 63.730 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 58.660 63.730 58.980 ;
      LAYER met4 ;
        RECT 63.410 58.660 63.730 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.410 58.250 63.730 58.570 ;
      LAYER met4 ;
        RECT 63.410 58.250 63.730 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 62.350 63.325 62.670 ;
      LAYER met4 ;
        RECT 63.005 62.350 63.325 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 61.940 63.325 62.260 ;
      LAYER met4 ;
        RECT 63.005 61.940 63.325 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 61.530 63.325 61.850 ;
      LAYER met4 ;
        RECT 63.005 61.530 63.325 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 61.120 63.325 61.440 ;
      LAYER met4 ;
        RECT 63.005 61.120 63.325 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 60.710 63.325 61.030 ;
      LAYER met4 ;
        RECT 63.005 60.710 63.325 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 60.300 63.325 60.620 ;
      LAYER met4 ;
        RECT 63.005 60.300 63.325 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 59.890 63.325 60.210 ;
      LAYER met4 ;
        RECT 63.005 59.890 63.325 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 59.480 63.325 59.800 ;
      LAYER met4 ;
        RECT 63.005 59.480 63.325 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 59.070 63.325 59.390 ;
      LAYER met4 ;
        RECT 63.005 59.070 63.325 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 58.660 63.325 58.980 ;
      LAYER met4 ;
        RECT 63.005 58.660 63.325 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.005 58.250 63.325 58.570 ;
      LAYER met4 ;
        RECT 63.005 58.250 63.325 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 62.350 62.920 62.670 ;
      LAYER met4 ;
        RECT 62.600 62.350 62.920 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 61.940 62.920 62.260 ;
      LAYER met4 ;
        RECT 62.600 61.940 62.920 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 61.530 62.920 61.850 ;
      LAYER met4 ;
        RECT 62.600 61.530 62.920 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 61.120 62.920 61.440 ;
      LAYER met4 ;
        RECT 62.600 61.120 62.920 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 60.710 62.920 61.030 ;
      LAYER met4 ;
        RECT 62.600 60.710 62.920 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 60.300 62.920 60.620 ;
      LAYER met4 ;
        RECT 62.600 60.300 62.920 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 59.890 62.920 60.210 ;
      LAYER met4 ;
        RECT 62.600 59.890 62.920 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 59.480 62.920 59.800 ;
      LAYER met4 ;
        RECT 62.600 59.480 62.920 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 59.070 62.920 59.390 ;
      LAYER met4 ;
        RECT 62.600 59.070 62.920 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 58.660 62.920 58.980 ;
      LAYER met4 ;
        RECT 62.600 58.660 62.920 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.600 58.250 62.920 58.570 ;
      LAYER met4 ;
        RECT 62.600 58.250 62.920 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 62.350 62.515 62.670 ;
      LAYER met4 ;
        RECT 62.195 62.350 62.515 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 61.940 62.515 62.260 ;
      LAYER met4 ;
        RECT 62.195 61.940 62.515 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 61.530 62.515 61.850 ;
      LAYER met4 ;
        RECT 62.195 61.530 62.515 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 61.120 62.515 61.440 ;
      LAYER met4 ;
        RECT 62.195 61.120 62.515 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 60.710 62.515 61.030 ;
      LAYER met4 ;
        RECT 62.195 60.710 62.515 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 60.300 62.515 60.620 ;
      LAYER met4 ;
        RECT 62.195 60.300 62.515 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 59.890 62.515 60.210 ;
      LAYER met4 ;
        RECT 62.195 59.890 62.515 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 59.480 62.515 59.800 ;
      LAYER met4 ;
        RECT 62.195 59.480 62.515 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 59.070 62.515 59.390 ;
      LAYER met4 ;
        RECT 62.195 59.070 62.515 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 58.660 62.515 58.980 ;
      LAYER met4 ;
        RECT 62.195 58.660 62.515 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.195 58.250 62.515 58.570 ;
      LAYER met4 ;
        RECT 62.195 58.250 62.515 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 62.350 62.110 62.670 ;
      LAYER met4 ;
        RECT 61.790 62.350 62.110 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 61.940 62.110 62.260 ;
      LAYER met4 ;
        RECT 61.790 61.940 62.110 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 61.530 62.110 61.850 ;
      LAYER met4 ;
        RECT 61.790 61.530 62.110 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 61.120 62.110 61.440 ;
      LAYER met4 ;
        RECT 61.790 61.120 62.110 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 60.710 62.110 61.030 ;
      LAYER met4 ;
        RECT 61.790 60.710 62.110 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 60.300 62.110 60.620 ;
      LAYER met4 ;
        RECT 61.790 60.300 62.110 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 59.890 62.110 60.210 ;
      LAYER met4 ;
        RECT 61.790 59.890 62.110 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 59.480 62.110 59.800 ;
      LAYER met4 ;
        RECT 61.790 59.480 62.110 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 59.070 62.110 59.390 ;
      LAYER met4 ;
        RECT 61.790 59.070 62.110 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 58.660 62.110 58.980 ;
      LAYER met4 ;
        RECT 61.790 58.660 62.110 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.790 58.250 62.110 58.570 ;
      LAYER met4 ;
        RECT 61.790 58.250 62.110 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 62.350 61.705 62.670 ;
      LAYER met4 ;
        RECT 61.385 62.350 61.705 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 61.940 61.705 62.260 ;
      LAYER met4 ;
        RECT 61.385 61.940 61.705 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 61.530 61.705 61.850 ;
      LAYER met4 ;
        RECT 61.385 61.530 61.705 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 61.120 61.705 61.440 ;
      LAYER met4 ;
        RECT 61.385 61.120 61.705 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 60.710 61.705 61.030 ;
      LAYER met4 ;
        RECT 61.385 60.710 61.705 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 60.300 61.705 60.620 ;
      LAYER met4 ;
        RECT 61.385 60.300 61.705 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 59.890 61.705 60.210 ;
      LAYER met4 ;
        RECT 61.385 59.890 61.705 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 59.480 61.705 59.800 ;
      LAYER met4 ;
        RECT 61.385 59.480 61.705 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 59.070 61.705 59.390 ;
      LAYER met4 ;
        RECT 61.385 59.070 61.705 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 58.660 61.705 58.980 ;
      LAYER met4 ;
        RECT 61.385 58.660 61.705 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.385 58.250 61.705 58.570 ;
      LAYER met4 ;
        RECT 61.385 58.250 61.705 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 62.350 61.300 62.670 ;
      LAYER met4 ;
        RECT 60.980 62.350 61.300 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 61.940 61.300 62.260 ;
      LAYER met4 ;
        RECT 60.980 61.940 61.300 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 61.530 61.300 61.850 ;
      LAYER met4 ;
        RECT 60.980 61.530 61.300 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 61.120 61.300 61.440 ;
      LAYER met4 ;
        RECT 60.980 61.120 61.300 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 60.710 61.300 61.030 ;
      LAYER met4 ;
        RECT 60.980 60.710 61.300 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 60.300 61.300 60.620 ;
      LAYER met4 ;
        RECT 60.980 60.300 61.300 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 59.890 61.300 60.210 ;
      LAYER met4 ;
        RECT 60.980 59.890 61.300 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 59.480 61.300 59.800 ;
      LAYER met4 ;
        RECT 60.980 59.480 61.300 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 59.070 61.300 59.390 ;
      LAYER met4 ;
        RECT 60.980 59.070 61.300 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 58.660 61.300 58.980 ;
      LAYER met4 ;
        RECT 60.980 58.660 61.300 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.980 58.250 61.300 58.570 ;
      LAYER met4 ;
        RECT 60.980 58.250 61.300 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 62.350 60.895 62.670 ;
      LAYER met4 ;
        RECT 60.575 62.350 60.895 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 61.940 60.895 62.260 ;
      LAYER met4 ;
        RECT 60.575 61.940 60.895 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 61.530 60.895 61.850 ;
      LAYER met4 ;
        RECT 60.575 61.530 60.895 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 61.120 60.895 61.440 ;
      LAYER met4 ;
        RECT 60.575 61.120 60.895 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 60.710 60.895 61.030 ;
      LAYER met4 ;
        RECT 60.575 60.710 60.895 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 60.300 60.895 60.620 ;
      LAYER met4 ;
        RECT 60.575 60.300 60.895 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 59.890 60.895 60.210 ;
      LAYER met4 ;
        RECT 60.575 59.890 60.895 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 59.480 60.895 59.800 ;
      LAYER met4 ;
        RECT 60.575 59.480 60.895 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 59.070 60.895 59.390 ;
      LAYER met4 ;
        RECT 60.575 59.070 60.895 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 58.660 60.895 58.980 ;
      LAYER met4 ;
        RECT 60.575 58.660 60.895 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.575 58.250 60.895 58.570 ;
      LAYER met4 ;
        RECT 60.575 58.250 60.895 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 62.350 60.490 62.670 ;
      LAYER met4 ;
        RECT 60.170 62.350 60.490 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 61.940 60.490 62.260 ;
      LAYER met4 ;
        RECT 60.170 61.940 60.490 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 61.530 60.490 61.850 ;
      LAYER met4 ;
        RECT 60.170 61.530 60.490 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 61.120 60.490 61.440 ;
      LAYER met4 ;
        RECT 60.170 61.120 60.490 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 60.710 60.490 61.030 ;
      LAYER met4 ;
        RECT 60.170 60.710 60.490 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 60.300 60.490 60.620 ;
      LAYER met4 ;
        RECT 60.170 60.300 60.490 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 59.890 60.490 60.210 ;
      LAYER met4 ;
        RECT 60.170 59.890 60.490 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 59.480 60.490 59.800 ;
      LAYER met4 ;
        RECT 60.170 59.480 60.490 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 59.070 60.490 59.390 ;
      LAYER met4 ;
        RECT 60.170 59.070 60.490 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 58.660 60.490 58.980 ;
      LAYER met4 ;
        RECT 60.170 58.660 60.490 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.170 58.250 60.490 58.570 ;
      LAYER met4 ;
        RECT 60.170 58.250 60.490 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 62.350 60.085 62.670 ;
      LAYER met4 ;
        RECT 59.765 62.350 60.085 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 61.940 60.085 62.260 ;
      LAYER met4 ;
        RECT 59.765 61.940 60.085 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 61.530 60.085 61.850 ;
      LAYER met4 ;
        RECT 59.765 61.530 60.085 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 61.120 60.085 61.440 ;
      LAYER met4 ;
        RECT 59.765 61.120 60.085 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 60.710 60.085 61.030 ;
      LAYER met4 ;
        RECT 59.765 60.710 60.085 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 60.300 60.085 60.620 ;
      LAYER met4 ;
        RECT 59.765 60.300 60.085 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 59.890 60.085 60.210 ;
      LAYER met4 ;
        RECT 59.765 59.890 60.085 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 59.480 60.085 59.800 ;
      LAYER met4 ;
        RECT 59.765 59.480 60.085 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 59.070 60.085 59.390 ;
      LAYER met4 ;
        RECT 59.765 59.070 60.085 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 58.660 60.085 58.980 ;
      LAYER met4 ;
        RECT 59.765 58.660 60.085 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.765 58.250 60.085 58.570 ;
      LAYER met4 ;
        RECT 59.765 58.250 60.085 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 62.350 59.680 62.670 ;
      LAYER met4 ;
        RECT 59.360 62.350 59.680 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 61.940 59.680 62.260 ;
      LAYER met4 ;
        RECT 59.360 61.940 59.680 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 61.530 59.680 61.850 ;
      LAYER met4 ;
        RECT 59.360 61.530 59.680 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 61.120 59.680 61.440 ;
      LAYER met4 ;
        RECT 59.360 61.120 59.680 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 60.710 59.680 61.030 ;
      LAYER met4 ;
        RECT 59.360 60.710 59.680 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 60.300 59.680 60.620 ;
      LAYER met4 ;
        RECT 59.360 60.300 59.680 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 59.890 59.680 60.210 ;
      LAYER met4 ;
        RECT 59.360 59.890 59.680 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 59.480 59.680 59.800 ;
      LAYER met4 ;
        RECT 59.360 59.480 59.680 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 59.070 59.680 59.390 ;
      LAYER met4 ;
        RECT 59.360 59.070 59.680 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 58.660 59.680 58.980 ;
      LAYER met4 ;
        RECT 59.360 58.660 59.680 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.360 58.250 59.680 58.570 ;
      LAYER met4 ;
        RECT 59.360 58.250 59.680 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 62.350 59.275 62.670 ;
      LAYER met4 ;
        RECT 58.955 62.350 59.275 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 61.940 59.275 62.260 ;
      LAYER met4 ;
        RECT 58.955 61.940 59.275 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 61.530 59.275 61.850 ;
      LAYER met4 ;
        RECT 58.955 61.530 59.275 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 61.120 59.275 61.440 ;
      LAYER met4 ;
        RECT 58.955 61.120 59.275 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 60.710 59.275 61.030 ;
      LAYER met4 ;
        RECT 58.955 60.710 59.275 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 60.300 59.275 60.620 ;
      LAYER met4 ;
        RECT 58.955 60.300 59.275 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 59.890 59.275 60.210 ;
      LAYER met4 ;
        RECT 58.955 59.890 59.275 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 59.480 59.275 59.800 ;
      LAYER met4 ;
        RECT 58.955 59.480 59.275 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 59.070 59.275 59.390 ;
      LAYER met4 ;
        RECT 58.955 59.070 59.275 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 58.660 59.275 58.980 ;
      LAYER met4 ;
        RECT 58.955 58.660 59.275 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.955 58.250 59.275 58.570 ;
      LAYER met4 ;
        RECT 58.955 58.250 59.275 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 62.350 58.870 62.670 ;
      LAYER met4 ;
        RECT 58.550 62.350 58.870 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 61.940 58.870 62.260 ;
      LAYER met4 ;
        RECT 58.550 61.940 58.870 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 61.530 58.870 61.850 ;
      LAYER met4 ;
        RECT 58.550 61.530 58.870 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 61.120 58.870 61.440 ;
      LAYER met4 ;
        RECT 58.550 61.120 58.870 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 60.710 58.870 61.030 ;
      LAYER met4 ;
        RECT 58.550 60.710 58.870 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 60.300 58.870 60.620 ;
      LAYER met4 ;
        RECT 58.550 60.300 58.870 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 59.890 58.870 60.210 ;
      LAYER met4 ;
        RECT 58.550 59.890 58.870 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 59.480 58.870 59.800 ;
      LAYER met4 ;
        RECT 58.550 59.480 58.870 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 59.070 58.870 59.390 ;
      LAYER met4 ;
        RECT 58.550 59.070 58.870 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 58.660 58.870 58.980 ;
      LAYER met4 ;
        RECT 58.550 58.660 58.870 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.550 58.250 58.870 58.570 ;
      LAYER met4 ;
        RECT 58.550 58.250 58.870 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 62.350 58.465 62.670 ;
      LAYER met4 ;
        RECT 58.145 62.350 58.465 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 61.940 58.465 62.260 ;
      LAYER met4 ;
        RECT 58.145 61.940 58.465 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 61.530 58.465 61.850 ;
      LAYER met4 ;
        RECT 58.145 61.530 58.465 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 61.120 58.465 61.440 ;
      LAYER met4 ;
        RECT 58.145 61.120 58.465 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 60.710 58.465 61.030 ;
      LAYER met4 ;
        RECT 58.145 60.710 58.465 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 60.300 58.465 60.620 ;
      LAYER met4 ;
        RECT 58.145 60.300 58.465 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 59.890 58.465 60.210 ;
      LAYER met4 ;
        RECT 58.145 59.890 58.465 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 59.480 58.465 59.800 ;
      LAYER met4 ;
        RECT 58.145 59.480 58.465 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 59.070 58.465 59.390 ;
      LAYER met4 ;
        RECT 58.145 59.070 58.465 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 58.660 58.465 58.980 ;
      LAYER met4 ;
        RECT 58.145 58.660 58.465 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.145 58.250 58.465 58.570 ;
      LAYER met4 ;
        RECT 58.145 58.250 58.465 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 62.350 58.060 62.670 ;
      LAYER met4 ;
        RECT 57.740 62.350 58.060 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 61.940 58.060 62.260 ;
      LAYER met4 ;
        RECT 57.740 61.940 58.060 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 61.530 58.060 61.850 ;
      LAYER met4 ;
        RECT 57.740 61.530 58.060 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 61.120 58.060 61.440 ;
      LAYER met4 ;
        RECT 57.740 61.120 58.060 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 60.710 58.060 61.030 ;
      LAYER met4 ;
        RECT 57.740 60.710 58.060 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 60.300 58.060 60.620 ;
      LAYER met4 ;
        RECT 57.740 60.300 58.060 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 59.890 58.060 60.210 ;
      LAYER met4 ;
        RECT 57.740 59.890 58.060 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 59.480 58.060 59.800 ;
      LAYER met4 ;
        RECT 57.740 59.480 58.060 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 59.070 58.060 59.390 ;
      LAYER met4 ;
        RECT 57.740 59.070 58.060 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 58.660 58.060 58.980 ;
      LAYER met4 ;
        RECT 57.740 58.660 58.060 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.740 58.250 58.060 58.570 ;
      LAYER met4 ;
        RECT 57.740 58.250 58.060 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 62.350 57.655 62.670 ;
      LAYER met4 ;
        RECT 57.335 62.350 57.655 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 61.940 57.655 62.260 ;
      LAYER met4 ;
        RECT 57.335 61.940 57.655 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 61.530 57.655 61.850 ;
      LAYER met4 ;
        RECT 57.335 61.530 57.655 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 61.120 57.655 61.440 ;
      LAYER met4 ;
        RECT 57.335 61.120 57.655 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 60.710 57.655 61.030 ;
      LAYER met4 ;
        RECT 57.335 60.710 57.655 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 60.300 57.655 60.620 ;
      LAYER met4 ;
        RECT 57.335 60.300 57.655 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 59.890 57.655 60.210 ;
      LAYER met4 ;
        RECT 57.335 59.890 57.655 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 59.480 57.655 59.800 ;
      LAYER met4 ;
        RECT 57.335 59.480 57.655 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 59.070 57.655 59.390 ;
      LAYER met4 ;
        RECT 57.335 59.070 57.655 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 58.660 57.655 58.980 ;
      LAYER met4 ;
        RECT 57.335 58.660 57.655 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.335 58.250 57.655 58.570 ;
      LAYER met4 ;
        RECT 57.335 58.250 57.655 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 62.350 57.250 62.670 ;
      LAYER met4 ;
        RECT 56.930 62.350 57.250 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 61.940 57.250 62.260 ;
      LAYER met4 ;
        RECT 56.930 61.940 57.250 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 61.530 57.250 61.850 ;
      LAYER met4 ;
        RECT 56.930 61.530 57.250 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 61.120 57.250 61.440 ;
      LAYER met4 ;
        RECT 56.930 61.120 57.250 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 60.710 57.250 61.030 ;
      LAYER met4 ;
        RECT 56.930 60.710 57.250 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 60.300 57.250 60.620 ;
      LAYER met4 ;
        RECT 56.930 60.300 57.250 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 59.890 57.250 60.210 ;
      LAYER met4 ;
        RECT 56.930 59.890 57.250 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 59.480 57.250 59.800 ;
      LAYER met4 ;
        RECT 56.930 59.480 57.250 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 59.070 57.250 59.390 ;
      LAYER met4 ;
        RECT 56.930 59.070 57.250 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 58.660 57.250 58.980 ;
      LAYER met4 ;
        RECT 56.930 58.660 57.250 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.930 58.250 57.250 58.570 ;
      LAYER met4 ;
        RECT 56.930 58.250 57.250 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 62.350 56.845 62.670 ;
      LAYER met4 ;
        RECT 56.525 62.350 56.845 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 61.940 56.845 62.260 ;
      LAYER met4 ;
        RECT 56.525 61.940 56.845 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 61.530 56.845 61.850 ;
      LAYER met4 ;
        RECT 56.525 61.530 56.845 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 61.120 56.845 61.440 ;
      LAYER met4 ;
        RECT 56.525 61.120 56.845 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 60.710 56.845 61.030 ;
      LAYER met4 ;
        RECT 56.525 60.710 56.845 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 60.300 56.845 60.620 ;
      LAYER met4 ;
        RECT 56.525 60.300 56.845 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 59.890 56.845 60.210 ;
      LAYER met4 ;
        RECT 56.525 59.890 56.845 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 59.480 56.845 59.800 ;
      LAYER met4 ;
        RECT 56.525 59.480 56.845 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 59.070 56.845 59.390 ;
      LAYER met4 ;
        RECT 56.525 59.070 56.845 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 58.660 56.845 58.980 ;
      LAYER met4 ;
        RECT 56.525 58.660 56.845 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.525 58.250 56.845 58.570 ;
      LAYER met4 ;
        RECT 56.525 58.250 56.845 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 62.350 56.440 62.670 ;
      LAYER met4 ;
        RECT 56.120 62.350 56.440 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 61.940 56.440 62.260 ;
      LAYER met4 ;
        RECT 56.120 61.940 56.440 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 61.530 56.440 61.850 ;
      LAYER met4 ;
        RECT 56.120 61.530 56.440 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 61.120 56.440 61.440 ;
      LAYER met4 ;
        RECT 56.120 61.120 56.440 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 60.710 56.440 61.030 ;
      LAYER met4 ;
        RECT 56.120 60.710 56.440 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 60.300 56.440 60.620 ;
      LAYER met4 ;
        RECT 56.120 60.300 56.440 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 59.890 56.440 60.210 ;
      LAYER met4 ;
        RECT 56.120 59.890 56.440 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 59.480 56.440 59.800 ;
      LAYER met4 ;
        RECT 56.120 59.480 56.440 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 59.070 56.440 59.390 ;
      LAYER met4 ;
        RECT 56.120 59.070 56.440 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 58.660 56.440 58.980 ;
      LAYER met4 ;
        RECT 56.120 58.660 56.440 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.120 58.250 56.440 58.570 ;
      LAYER met4 ;
        RECT 56.120 58.250 56.440 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 62.350 56.035 62.670 ;
      LAYER met4 ;
        RECT 55.715 62.350 56.035 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 61.940 56.035 62.260 ;
      LAYER met4 ;
        RECT 55.715 61.940 56.035 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 61.530 56.035 61.850 ;
      LAYER met4 ;
        RECT 55.715 61.530 56.035 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 61.120 56.035 61.440 ;
      LAYER met4 ;
        RECT 55.715 61.120 56.035 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 60.710 56.035 61.030 ;
      LAYER met4 ;
        RECT 55.715 60.710 56.035 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 60.300 56.035 60.620 ;
      LAYER met4 ;
        RECT 55.715 60.300 56.035 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 59.890 56.035 60.210 ;
      LAYER met4 ;
        RECT 55.715 59.890 56.035 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 59.480 56.035 59.800 ;
      LAYER met4 ;
        RECT 55.715 59.480 56.035 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 59.070 56.035 59.390 ;
      LAYER met4 ;
        RECT 55.715 59.070 56.035 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 58.660 56.035 58.980 ;
      LAYER met4 ;
        RECT 55.715 58.660 56.035 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.715 58.250 56.035 58.570 ;
      LAYER met4 ;
        RECT 55.715 58.250 56.035 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 62.350 55.630 62.670 ;
      LAYER met4 ;
        RECT 55.310 62.350 55.630 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 61.940 55.630 62.260 ;
      LAYER met4 ;
        RECT 55.310 61.940 55.630 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 61.530 55.630 61.850 ;
      LAYER met4 ;
        RECT 55.310 61.530 55.630 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 61.120 55.630 61.440 ;
      LAYER met4 ;
        RECT 55.310 61.120 55.630 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 60.710 55.630 61.030 ;
      LAYER met4 ;
        RECT 55.310 60.710 55.630 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 60.300 55.630 60.620 ;
      LAYER met4 ;
        RECT 55.310 60.300 55.630 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 59.890 55.630 60.210 ;
      LAYER met4 ;
        RECT 55.310 59.890 55.630 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 59.480 55.630 59.800 ;
      LAYER met4 ;
        RECT 55.310 59.480 55.630 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 59.070 55.630 59.390 ;
      LAYER met4 ;
        RECT 55.310 59.070 55.630 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 58.660 55.630 58.980 ;
      LAYER met4 ;
        RECT 55.310 58.660 55.630 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.310 58.250 55.630 58.570 ;
      LAYER met4 ;
        RECT 55.310 58.250 55.630 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 62.350 55.225 62.670 ;
      LAYER met4 ;
        RECT 54.905 62.350 55.225 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 61.940 55.225 62.260 ;
      LAYER met4 ;
        RECT 54.905 61.940 55.225 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 61.530 55.225 61.850 ;
      LAYER met4 ;
        RECT 54.905 61.530 55.225 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 61.120 55.225 61.440 ;
      LAYER met4 ;
        RECT 54.905 61.120 55.225 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 60.710 55.225 61.030 ;
      LAYER met4 ;
        RECT 54.905 60.710 55.225 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 60.300 55.225 60.620 ;
      LAYER met4 ;
        RECT 54.905 60.300 55.225 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 59.890 55.225 60.210 ;
      LAYER met4 ;
        RECT 54.905 59.890 55.225 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 59.480 55.225 59.800 ;
      LAYER met4 ;
        RECT 54.905 59.480 55.225 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 59.070 55.225 59.390 ;
      LAYER met4 ;
        RECT 54.905 59.070 55.225 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 58.660 55.225 58.980 ;
      LAYER met4 ;
        RECT 54.905 58.660 55.225 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.905 58.250 55.225 58.570 ;
      LAYER met4 ;
        RECT 54.905 58.250 55.225 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 62.350 54.820 62.670 ;
      LAYER met4 ;
        RECT 54.500 62.350 54.820 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 61.940 54.820 62.260 ;
      LAYER met4 ;
        RECT 54.500 61.940 54.820 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 61.530 54.820 61.850 ;
      LAYER met4 ;
        RECT 54.500 61.530 54.820 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 61.120 54.820 61.440 ;
      LAYER met4 ;
        RECT 54.500 61.120 54.820 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 60.710 54.820 61.030 ;
      LAYER met4 ;
        RECT 54.500 60.710 54.820 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 60.300 54.820 60.620 ;
      LAYER met4 ;
        RECT 54.500 60.300 54.820 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 59.890 54.820 60.210 ;
      LAYER met4 ;
        RECT 54.500 59.890 54.820 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 59.480 54.820 59.800 ;
      LAYER met4 ;
        RECT 54.500 59.480 54.820 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 59.070 54.820 59.390 ;
      LAYER met4 ;
        RECT 54.500 59.070 54.820 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 58.660 54.820 58.980 ;
      LAYER met4 ;
        RECT 54.500 58.660 54.820 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.500 58.250 54.820 58.570 ;
      LAYER met4 ;
        RECT 54.500 58.250 54.820 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 62.350 54.415 62.670 ;
      LAYER met4 ;
        RECT 54.095 62.350 54.415 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 61.940 54.415 62.260 ;
      LAYER met4 ;
        RECT 54.095 61.940 54.415 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 61.530 54.415 61.850 ;
      LAYER met4 ;
        RECT 54.095 61.530 54.415 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 61.120 54.415 61.440 ;
      LAYER met4 ;
        RECT 54.095 61.120 54.415 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 60.710 54.415 61.030 ;
      LAYER met4 ;
        RECT 54.095 60.710 54.415 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 60.300 54.415 60.620 ;
      LAYER met4 ;
        RECT 54.095 60.300 54.415 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 59.890 54.415 60.210 ;
      LAYER met4 ;
        RECT 54.095 59.890 54.415 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 59.480 54.415 59.800 ;
      LAYER met4 ;
        RECT 54.095 59.480 54.415 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 59.070 54.415 59.390 ;
      LAYER met4 ;
        RECT 54.095 59.070 54.415 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 58.660 54.415 58.980 ;
      LAYER met4 ;
        RECT 54.095 58.660 54.415 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.095 58.250 54.415 58.570 ;
      LAYER met4 ;
        RECT 54.095 58.250 54.415 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 62.350 54.010 62.670 ;
      LAYER met4 ;
        RECT 53.690 62.350 54.010 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 61.940 54.010 62.260 ;
      LAYER met4 ;
        RECT 53.690 61.940 54.010 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 61.530 54.010 61.850 ;
      LAYER met4 ;
        RECT 53.690 61.530 54.010 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 61.120 54.010 61.440 ;
      LAYER met4 ;
        RECT 53.690 61.120 54.010 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 60.710 54.010 61.030 ;
      LAYER met4 ;
        RECT 53.690 60.710 54.010 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 60.300 54.010 60.620 ;
      LAYER met4 ;
        RECT 53.690 60.300 54.010 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 59.890 54.010 60.210 ;
      LAYER met4 ;
        RECT 53.690 59.890 54.010 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 59.480 54.010 59.800 ;
      LAYER met4 ;
        RECT 53.690 59.480 54.010 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 59.070 54.010 59.390 ;
      LAYER met4 ;
        RECT 53.690 59.070 54.010 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 58.660 54.010 58.980 ;
      LAYER met4 ;
        RECT 53.690 58.660 54.010 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.690 58.250 54.010 58.570 ;
      LAYER met4 ;
        RECT 53.690 58.250 54.010 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 62.350 53.605 62.670 ;
      LAYER met4 ;
        RECT 53.285 62.350 53.605 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 61.940 53.605 62.260 ;
      LAYER met4 ;
        RECT 53.285 61.940 53.605 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 61.530 53.605 61.850 ;
      LAYER met4 ;
        RECT 53.285 61.530 53.605 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 61.120 53.605 61.440 ;
      LAYER met4 ;
        RECT 53.285 61.120 53.605 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 60.710 53.605 61.030 ;
      LAYER met4 ;
        RECT 53.285 60.710 53.605 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 60.300 53.605 60.620 ;
      LAYER met4 ;
        RECT 53.285 60.300 53.605 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 59.890 53.605 60.210 ;
      LAYER met4 ;
        RECT 53.285 59.890 53.605 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 59.480 53.605 59.800 ;
      LAYER met4 ;
        RECT 53.285 59.480 53.605 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 59.070 53.605 59.390 ;
      LAYER met4 ;
        RECT 53.285 59.070 53.605 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 58.660 53.605 58.980 ;
      LAYER met4 ;
        RECT 53.285 58.660 53.605 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 58.250 53.605 58.570 ;
      LAYER met4 ;
        RECT 53.285 58.250 53.605 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 62.350 53.200 62.670 ;
      LAYER met4 ;
        RECT 52.880 62.350 53.200 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 61.940 53.200 62.260 ;
      LAYER met4 ;
        RECT 52.880 61.940 53.200 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 61.530 53.200 61.850 ;
      LAYER met4 ;
        RECT 52.880 61.530 53.200 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 61.120 53.200 61.440 ;
      LAYER met4 ;
        RECT 52.880 61.120 53.200 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 60.710 53.200 61.030 ;
      LAYER met4 ;
        RECT 52.880 60.710 53.200 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 60.300 53.200 60.620 ;
      LAYER met4 ;
        RECT 52.880 60.300 53.200 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 59.890 53.200 60.210 ;
      LAYER met4 ;
        RECT 52.880 59.890 53.200 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 59.480 53.200 59.800 ;
      LAYER met4 ;
        RECT 52.880 59.480 53.200 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 59.070 53.200 59.390 ;
      LAYER met4 ;
        RECT 52.880 59.070 53.200 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 58.660 53.200 58.980 ;
      LAYER met4 ;
        RECT 52.880 58.660 53.200 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.880 58.250 53.200 58.570 ;
      LAYER met4 ;
        RECT 52.880 58.250 53.200 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 62.350 52.790 62.670 ;
      LAYER met4 ;
        RECT 52.470 62.350 52.790 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 61.940 52.790 62.260 ;
      LAYER met4 ;
        RECT 52.470 61.940 52.790 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 61.530 52.790 61.850 ;
      LAYER met4 ;
        RECT 52.470 61.530 52.790 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 61.120 52.790 61.440 ;
      LAYER met4 ;
        RECT 52.470 61.120 52.790 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 60.710 52.790 61.030 ;
      LAYER met4 ;
        RECT 52.470 60.710 52.790 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 60.300 52.790 60.620 ;
      LAYER met4 ;
        RECT 52.470 60.300 52.790 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 59.890 52.790 60.210 ;
      LAYER met4 ;
        RECT 52.470 59.890 52.790 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 59.480 52.790 59.800 ;
      LAYER met4 ;
        RECT 52.470 59.480 52.790 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 59.070 52.790 59.390 ;
      LAYER met4 ;
        RECT 52.470 59.070 52.790 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 58.660 52.790 58.980 ;
      LAYER met4 ;
        RECT 52.470 58.660 52.790 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.470 58.250 52.790 58.570 ;
      LAYER met4 ;
        RECT 52.470 58.250 52.790 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 62.350 52.380 62.670 ;
      LAYER met4 ;
        RECT 52.060 62.350 52.380 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 61.940 52.380 62.260 ;
      LAYER met4 ;
        RECT 52.060 61.940 52.380 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 61.530 52.380 61.850 ;
      LAYER met4 ;
        RECT 52.060 61.530 52.380 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 61.120 52.380 61.440 ;
      LAYER met4 ;
        RECT 52.060 61.120 52.380 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 60.710 52.380 61.030 ;
      LAYER met4 ;
        RECT 52.060 60.710 52.380 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 60.300 52.380 60.620 ;
      LAYER met4 ;
        RECT 52.060 60.300 52.380 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 59.890 52.380 60.210 ;
      LAYER met4 ;
        RECT 52.060 59.890 52.380 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 59.480 52.380 59.800 ;
      LAYER met4 ;
        RECT 52.060 59.480 52.380 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 59.070 52.380 59.390 ;
      LAYER met4 ;
        RECT 52.060 59.070 52.380 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 58.660 52.380 58.980 ;
      LAYER met4 ;
        RECT 52.060 58.660 52.380 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.060 58.250 52.380 58.570 ;
      LAYER met4 ;
        RECT 52.060 58.250 52.380 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 62.350 51.970 62.670 ;
      LAYER met4 ;
        RECT 51.650 62.350 51.970 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 61.940 51.970 62.260 ;
      LAYER met4 ;
        RECT 51.650 61.940 51.970 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 61.530 51.970 61.850 ;
      LAYER met4 ;
        RECT 51.650 61.530 51.970 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 61.120 51.970 61.440 ;
      LAYER met4 ;
        RECT 51.650 61.120 51.970 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 60.710 51.970 61.030 ;
      LAYER met4 ;
        RECT 51.650 60.710 51.970 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 60.300 51.970 60.620 ;
      LAYER met4 ;
        RECT 51.650 60.300 51.970 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 59.890 51.970 60.210 ;
      LAYER met4 ;
        RECT 51.650 59.890 51.970 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 59.480 51.970 59.800 ;
      LAYER met4 ;
        RECT 51.650 59.480 51.970 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 59.070 51.970 59.390 ;
      LAYER met4 ;
        RECT 51.650 59.070 51.970 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 58.660 51.970 58.980 ;
      LAYER met4 ;
        RECT 51.650 58.660 51.970 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.650 58.250 51.970 58.570 ;
      LAYER met4 ;
        RECT 51.650 58.250 51.970 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 62.350 51.560 62.670 ;
      LAYER met4 ;
        RECT 51.240 62.350 51.560 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 61.940 51.560 62.260 ;
      LAYER met4 ;
        RECT 51.240 61.940 51.560 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 61.530 51.560 61.850 ;
      LAYER met4 ;
        RECT 51.240 61.530 51.560 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 61.120 51.560 61.440 ;
      LAYER met4 ;
        RECT 51.240 61.120 51.560 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 60.710 51.560 61.030 ;
      LAYER met4 ;
        RECT 51.240 60.710 51.560 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 60.300 51.560 60.620 ;
      LAYER met4 ;
        RECT 51.240 60.300 51.560 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 59.890 51.560 60.210 ;
      LAYER met4 ;
        RECT 51.240 59.890 51.560 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 59.480 51.560 59.800 ;
      LAYER met4 ;
        RECT 51.240 59.480 51.560 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 59.070 51.560 59.390 ;
      LAYER met4 ;
        RECT 51.240 59.070 51.560 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 58.660 51.560 58.980 ;
      LAYER met4 ;
        RECT 51.240 58.660 51.560 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.240 58.250 51.560 58.570 ;
      LAYER met4 ;
        RECT 51.240 58.250 51.560 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 62.350 51.150 62.670 ;
      LAYER met4 ;
        RECT 50.830 62.350 51.150 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 61.940 51.150 62.260 ;
      LAYER met4 ;
        RECT 50.830 61.940 51.150 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 61.530 51.150 61.850 ;
      LAYER met4 ;
        RECT 50.830 61.530 51.150 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 61.120 51.150 61.440 ;
      LAYER met4 ;
        RECT 50.830 61.120 51.150 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 60.710 51.150 61.030 ;
      LAYER met4 ;
        RECT 50.830 60.710 51.150 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 60.300 51.150 60.620 ;
      LAYER met4 ;
        RECT 50.830 60.300 51.150 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 59.890 51.150 60.210 ;
      LAYER met4 ;
        RECT 50.830 59.890 51.150 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 59.480 51.150 59.800 ;
      LAYER met4 ;
        RECT 50.830 59.480 51.150 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 59.070 51.150 59.390 ;
      LAYER met4 ;
        RECT 50.830 59.070 51.150 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 58.660 51.150 58.980 ;
      LAYER met4 ;
        RECT 50.830 58.660 51.150 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.830 58.250 51.150 58.570 ;
      LAYER met4 ;
        RECT 50.830 58.250 51.150 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 62.350 50.740 62.670 ;
      LAYER met4 ;
        RECT 50.420 62.350 50.740 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 61.940 50.740 62.260 ;
      LAYER met4 ;
        RECT 50.420 61.940 50.740 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 61.530 50.740 61.850 ;
      LAYER met4 ;
        RECT 50.420 61.530 50.740 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 61.120 50.740 61.440 ;
      LAYER met4 ;
        RECT 50.420 61.120 50.740 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 60.710 50.740 61.030 ;
      LAYER met4 ;
        RECT 50.420 60.710 50.740 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 60.300 50.740 60.620 ;
      LAYER met4 ;
        RECT 50.420 60.300 50.740 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 59.890 50.740 60.210 ;
      LAYER met4 ;
        RECT 50.420 59.890 50.740 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 59.480 50.740 59.800 ;
      LAYER met4 ;
        RECT 50.420 59.480 50.740 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 59.070 50.740 59.390 ;
      LAYER met4 ;
        RECT 50.420 59.070 50.740 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 58.660 50.740 58.980 ;
      LAYER met4 ;
        RECT 50.420 58.660 50.740 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.420 58.250 50.740 58.570 ;
      LAYER met4 ;
        RECT 50.420 58.250 50.740 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 62.350 24.365 62.670 ;
      LAYER met4 ;
        RECT 24.045 62.350 24.365 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 61.940 24.365 62.260 ;
      LAYER met4 ;
        RECT 24.045 61.940 24.365 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 61.530 24.365 61.850 ;
      LAYER met4 ;
        RECT 24.045 61.530 24.365 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 61.120 24.365 61.440 ;
      LAYER met4 ;
        RECT 24.045 61.120 24.365 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 60.710 24.365 61.030 ;
      LAYER met4 ;
        RECT 24.045 60.710 24.365 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 60.300 24.365 60.620 ;
      LAYER met4 ;
        RECT 24.045 60.300 24.365 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 59.890 24.365 60.210 ;
      LAYER met4 ;
        RECT 24.045 59.890 24.365 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 59.480 24.365 59.800 ;
      LAYER met4 ;
        RECT 24.045 59.480 24.365 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 59.070 24.365 59.390 ;
      LAYER met4 ;
        RECT 24.045 59.070 24.365 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 58.660 24.365 58.980 ;
      LAYER met4 ;
        RECT 24.045 58.660 24.365 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.045 58.250 24.365 58.570 ;
      LAYER met4 ;
        RECT 24.045 58.250 24.365 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 62.350 23.960 62.670 ;
      LAYER met4 ;
        RECT 23.640 62.350 23.960 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 61.940 23.960 62.260 ;
      LAYER met4 ;
        RECT 23.640 61.940 23.960 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 61.530 23.960 61.850 ;
      LAYER met4 ;
        RECT 23.640 61.530 23.960 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 61.120 23.960 61.440 ;
      LAYER met4 ;
        RECT 23.640 61.120 23.960 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 60.710 23.960 61.030 ;
      LAYER met4 ;
        RECT 23.640 60.710 23.960 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 60.300 23.960 60.620 ;
      LAYER met4 ;
        RECT 23.640 60.300 23.960 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 59.890 23.960 60.210 ;
      LAYER met4 ;
        RECT 23.640 59.890 23.960 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 59.480 23.960 59.800 ;
      LAYER met4 ;
        RECT 23.640 59.480 23.960 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 59.070 23.960 59.390 ;
      LAYER met4 ;
        RECT 23.640 59.070 23.960 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 58.660 23.960 58.980 ;
      LAYER met4 ;
        RECT 23.640 58.660 23.960 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.640 58.250 23.960 58.570 ;
      LAYER met4 ;
        RECT 23.640 58.250 23.960 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 62.350 23.555 62.670 ;
      LAYER met4 ;
        RECT 23.235 62.350 23.555 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 61.940 23.555 62.260 ;
      LAYER met4 ;
        RECT 23.235 61.940 23.555 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 61.530 23.555 61.850 ;
      LAYER met4 ;
        RECT 23.235 61.530 23.555 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 61.120 23.555 61.440 ;
      LAYER met4 ;
        RECT 23.235 61.120 23.555 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 60.710 23.555 61.030 ;
      LAYER met4 ;
        RECT 23.235 60.710 23.555 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 60.300 23.555 60.620 ;
      LAYER met4 ;
        RECT 23.235 60.300 23.555 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 59.890 23.555 60.210 ;
      LAYER met4 ;
        RECT 23.235 59.890 23.555 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 59.480 23.555 59.800 ;
      LAYER met4 ;
        RECT 23.235 59.480 23.555 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 59.070 23.555 59.390 ;
      LAYER met4 ;
        RECT 23.235 59.070 23.555 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 58.660 23.555 58.980 ;
      LAYER met4 ;
        RECT 23.235 58.660 23.555 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.235 58.250 23.555 58.570 ;
      LAYER met4 ;
        RECT 23.235 58.250 23.555 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 62.350 23.150 62.670 ;
      LAYER met4 ;
        RECT 22.830 62.350 23.150 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 61.940 23.150 62.260 ;
      LAYER met4 ;
        RECT 22.830 61.940 23.150 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 61.530 23.150 61.850 ;
      LAYER met4 ;
        RECT 22.830 61.530 23.150 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 61.120 23.150 61.440 ;
      LAYER met4 ;
        RECT 22.830 61.120 23.150 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 60.710 23.150 61.030 ;
      LAYER met4 ;
        RECT 22.830 60.710 23.150 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 60.300 23.150 60.620 ;
      LAYER met4 ;
        RECT 22.830 60.300 23.150 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 59.890 23.150 60.210 ;
      LAYER met4 ;
        RECT 22.830 59.890 23.150 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 59.480 23.150 59.800 ;
      LAYER met4 ;
        RECT 22.830 59.480 23.150 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 59.070 23.150 59.390 ;
      LAYER met4 ;
        RECT 22.830 59.070 23.150 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 58.660 23.150 58.980 ;
      LAYER met4 ;
        RECT 22.830 58.660 23.150 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.830 58.250 23.150 58.570 ;
      LAYER met4 ;
        RECT 22.830 58.250 23.150 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 62.350 22.745 62.670 ;
      LAYER met4 ;
        RECT 22.425 62.350 22.745 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 61.940 22.745 62.260 ;
      LAYER met4 ;
        RECT 22.425 61.940 22.745 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 61.530 22.745 61.850 ;
      LAYER met4 ;
        RECT 22.425 61.530 22.745 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 61.120 22.745 61.440 ;
      LAYER met4 ;
        RECT 22.425 61.120 22.745 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 60.710 22.745 61.030 ;
      LAYER met4 ;
        RECT 22.425 60.710 22.745 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 60.300 22.745 60.620 ;
      LAYER met4 ;
        RECT 22.425 60.300 22.745 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 59.890 22.745 60.210 ;
      LAYER met4 ;
        RECT 22.425 59.890 22.745 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 59.480 22.745 59.800 ;
      LAYER met4 ;
        RECT 22.425 59.480 22.745 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 59.070 22.745 59.390 ;
      LAYER met4 ;
        RECT 22.425 59.070 22.745 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 58.660 22.745 58.980 ;
      LAYER met4 ;
        RECT 22.425 58.660 22.745 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.425 58.250 22.745 58.570 ;
      LAYER met4 ;
        RECT 22.425 58.250 22.745 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 62.350 22.340 62.670 ;
      LAYER met4 ;
        RECT 22.020 62.350 22.340 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 61.940 22.340 62.260 ;
      LAYER met4 ;
        RECT 22.020 61.940 22.340 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 61.530 22.340 61.850 ;
      LAYER met4 ;
        RECT 22.020 61.530 22.340 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 61.120 22.340 61.440 ;
      LAYER met4 ;
        RECT 22.020 61.120 22.340 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 60.710 22.340 61.030 ;
      LAYER met4 ;
        RECT 22.020 60.710 22.340 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 60.300 22.340 60.620 ;
      LAYER met4 ;
        RECT 22.020 60.300 22.340 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 59.890 22.340 60.210 ;
      LAYER met4 ;
        RECT 22.020 59.890 22.340 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 59.480 22.340 59.800 ;
      LAYER met4 ;
        RECT 22.020 59.480 22.340 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 59.070 22.340 59.390 ;
      LAYER met4 ;
        RECT 22.020 59.070 22.340 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 58.660 22.340 58.980 ;
      LAYER met4 ;
        RECT 22.020 58.660 22.340 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.020 58.250 22.340 58.570 ;
      LAYER met4 ;
        RECT 22.020 58.250 22.340 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 62.350 21.935 62.670 ;
      LAYER met4 ;
        RECT 21.615 62.350 21.935 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 61.940 21.935 62.260 ;
      LAYER met4 ;
        RECT 21.615 61.940 21.935 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 61.530 21.935 61.850 ;
      LAYER met4 ;
        RECT 21.615 61.530 21.935 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 61.120 21.935 61.440 ;
      LAYER met4 ;
        RECT 21.615 61.120 21.935 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 60.710 21.935 61.030 ;
      LAYER met4 ;
        RECT 21.615 60.710 21.935 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 60.300 21.935 60.620 ;
      LAYER met4 ;
        RECT 21.615 60.300 21.935 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 59.890 21.935 60.210 ;
      LAYER met4 ;
        RECT 21.615 59.890 21.935 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 59.480 21.935 59.800 ;
      LAYER met4 ;
        RECT 21.615 59.480 21.935 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 59.070 21.935 59.390 ;
      LAYER met4 ;
        RECT 21.615 59.070 21.935 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 58.660 21.935 58.980 ;
      LAYER met4 ;
        RECT 21.615 58.660 21.935 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.615 58.250 21.935 58.570 ;
      LAYER met4 ;
        RECT 21.615 58.250 21.935 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 62.350 21.530 62.670 ;
      LAYER met4 ;
        RECT 21.210 62.350 21.530 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 61.940 21.530 62.260 ;
      LAYER met4 ;
        RECT 21.210 61.940 21.530 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 61.530 21.530 61.850 ;
      LAYER met4 ;
        RECT 21.210 61.530 21.530 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 61.120 21.530 61.440 ;
      LAYER met4 ;
        RECT 21.210 61.120 21.530 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 60.710 21.530 61.030 ;
      LAYER met4 ;
        RECT 21.210 60.710 21.530 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 60.300 21.530 60.620 ;
      LAYER met4 ;
        RECT 21.210 60.300 21.530 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 59.890 21.530 60.210 ;
      LAYER met4 ;
        RECT 21.210 59.890 21.530 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 59.480 21.530 59.800 ;
      LAYER met4 ;
        RECT 21.210 59.480 21.530 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 59.070 21.530 59.390 ;
      LAYER met4 ;
        RECT 21.210 59.070 21.530 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 58.660 21.530 58.980 ;
      LAYER met4 ;
        RECT 21.210 58.660 21.530 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.210 58.250 21.530 58.570 ;
      LAYER met4 ;
        RECT 21.210 58.250 21.530 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 62.350 21.125 62.670 ;
      LAYER met4 ;
        RECT 20.805 62.350 21.125 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 61.940 21.125 62.260 ;
      LAYER met4 ;
        RECT 20.805 61.940 21.125 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 61.530 21.125 61.850 ;
      LAYER met4 ;
        RECT 20.805 61.530 21.125 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 61.120 21.125 61.440 ;
      LAYER met4 ;
        RECT 20.805 61.120 21.125 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 60.710 21.125 61.030 ;
      LAYER met4 ;
        RECT 20.805 60.710 21.125 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 60.300 21.125 60.620 ;
      LAYER met4 ;
        RECT 20.805 60.300 21.125 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 59.890 21.125 60.210 ;
      LAYER met4 ;
        RECT 20.805 59.890 21.125 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 59.480 21.125 59.800 ;
      LAYER met4 ;
        RECT 20.805 59.480 21.125 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 59.070 21.125 59.390 ;
      LAYER met4 ;
        RECT 20.805 59.070 21.125 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 58.660 21.125 58.980 ;
      LAYER met4 ;
        RECT 20.805 58.660 21.125 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.805 58.250 21.125 58.570 ;
      LAYER met4 ;
        RECT 20.805 58.250 21.125 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 62.350 20.720 62.670 ;
      LAYER met4 ;
        RECT 20.400 62.350 20.720 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 61.940 20.720 62.260 ;
      LAYER met4 ;
        RECT 20.400 61.940 20.720 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 61.530 20.720 61.850 ;
      LAYER met4 ;
        RECT 20.400 61.530 20.720 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 61.120 20.720 61.440 ;
      LAYER met4 ;
        RECT 20.400 61.120 20.720 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 60.710 20.720 61.030 ;
      LAYER met4 ;
        RECT 20.400 60.710 20.720 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 60.300 20.720 60.620 ;
      LAYER met4 ;
        RECT 20.400 60.300 20.720 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 59.890 20.720 60.210 ;
      LAYER met4 ;
        RECT 20.400 59.890 20.720 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 59.480 20.720 59.800 ;
      LAYER met4 ;
        RECT 20.400 59.480 20.720 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 59.070 20.720 59.390 ;
      LAYER met4 ;
        RECT 20.400 59.070 20.720 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 58.660 20.720 58.980 ;
      LAYER met4 ;
        RECT 20.400 58.660 20.720 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.400 58.250 20.720 58.570 ;
      LAYER met4 ;
        RECT 20.400 58.250 20.720 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 62.350 20.315 62.670 ;
      LAYER met4 ;
        RECT 19.995 62.350 20.315 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 61.940 20.315 62.260 ;
      LAYER met4 ;
        RECT 19.995 61.940 20.315 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 61.530 20.315 61.850 ;
      LAYER met4 ;
        RECT 19.995 61.530 20.315 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 61.120 20.315 61.440 ;
      LAYER met4 ;
        RECT 19.995 61.120 20.315 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 60.710 20.315 61.030 ;
      LAYER met4 ;
        RECT 19.995 60.710 20.315 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 60.300 20.315 60.620 ;
      LAYER met4 ;
        RECT 19.995 60.300 20.315 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 59.890 20.315 60.210 ;
      LAYER met4 ;
        RECT 19.995 59.890 20.315 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 59.480 20.315 59.800 ;
      LAYER met4 ;
        RECT 19.995 59.480 20.315 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 59.070 20.315 59.390 ;
      LAYER met4 ;
        RECT 19.995 59.070 20.315 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 58.660 20.315 58.980 ;
      LAYER met4 ;
        RECT 19.995 58.660 20.315 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 58.250 20.315 58.570 ;
      LAYER met4 ;
        RECT 19.995 58.250 20.315 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 62.350 19.910 62.670 ;
      LAYER met4 ;
        RECT 19.590 62.350 19.910 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 61.940 19.910 62.260 ;
      LAYER met4 ;
        RECT 19.590 61.940 19.910 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 61.530 19.910 61.850 ;
      LAYER met4 ;
        RECT 19.590 61.530 19.910 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 61.120 19.910 61.440 ;
      LAYER met4 ;
        RECT 19.590 61.120 19.910 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 60.710 19.910 61.030 ;
      LAYER met4 ;
        RECT 19.590 60.710 19.910 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 60.300 19.910 60.620 ;
      LAYER met4 ;
        RECT 19.590 60.300 19.910 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 59.890 19.910 60.210 ;
      LAYER met4 ;
        RECT 19.590 59.890 19.910 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 59.480 19.910 59.800 ;
      LAYER met4 ;
        RECT 19.590 59.480 19.910 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 59.070 19.910 59.390 ;
      LAYER met4 ;
        RECT 19.590 59.070 19.910 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 58.660 19.910 58.980 ;
      LAYER met4 ;
        RECT 19.590 58.660 19.910 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.590 58.250 19.910 58.570 ;
      LAYER met4 ;
        RECT 19.590 58.250 19.910 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 62.350 19.505 62.670 ;
      LAYER met4 ;
        RECT 19.185 62.350 19.505 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 61.940 19.505 62.260 ;
      LAYER met4 ;
        RECT 19.185 61.940 19.505 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 61.530 19.505 61.850 ;
      LAYER met4 ;
        RECT 19.185 61.530 19.505 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 61.120 19.505 61.440 ;
      LAYER met4 ;
        RECT 19.185 61.120 19.505 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 60.710 19.505 61.030 ;
      LAYER met4 ;
        RECT 19.185 60.710 19.505 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 60.300 19.505 60.620 ;
      LAYER met4 ;
        RECT 19.185 60.300 19.505 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 59.890 19.505 60.210 ;
      LAYER met4 ;
        RECT 19.185 59.890 19.505 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 59.480 19.505 59.800 ;
      LAYER met4 ;
        RECT 19.185 59.480 19.505 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 59.070 19.505 59.390 ;
      LAYER met4 ;
        RECT 19.185 59.070 19.505 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 58.660 19.505 58.980 ;
      LAYER met4 ;
        RECT 19.185 58.660 19.505 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.185 58.250 19.505 58.570 ;
      LAYER met4 ;
        RECT 19.185 58.250 19.505 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 62.350 19.100 62.670 ;
      LAYER met4 ;
        RECT 18.780 62.350 19.100 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 61.940 19.100 62.260 ;
      LAYER met4 ;
        RECT 18.780 61.940 19.100 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 61.530 19.100 61.850 ;
      LAYER met4 ;
        RECT 18.780 61.530 19.100 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 61.120 19.100 61.440 ;
      LAYER met4 ;
        RECT 18.780 61.120 19.100 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 60.710 19.100 61.030 ;
      LAYER met4 ;
        RECT 18.780 60.710 19.100 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 60.300 19.100 60.620 ;
      LAYER met4 ;
        RECT 18.780 60.300 19.100 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 59.890 19.100 60.210 ;
      LAYER met4 ;
        RECT 18.780 59.890 19.100 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 59.480 19.100 59.800 ;
      LAYER met4 ;
        RECT 18.780 59.480 19.100 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 59.070 19.100 59.390 ;
      LAYER met4 ;
        RECT 18.780 59.070 19.100 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 58.660 19.100 58.980 ;
      LAYER met4 ;
        RECT 18.780 58.660 19.100 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.780 58.250 19.100 58.570 ;
      LAYER met4 ;
        RECT 18.780 58.250 19.100 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 62.350 18.695 62.670 ;
      LAYER met4 ;
        RECT 18.375 62.350 18.695 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 61.940 18.695 62.260 ;
      LAYER met4 ;
        RECT 18.375 61.940 18.695 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 61.530 18.695 61.850 ;
      LAYER met4 ;
        RECT 18.375 61.530 18.695 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 61.120 18.695 61.440 ;
      LAYER met4 ;
        RECT 18.375 61.120 18.695 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 60.710 18.695 61.030 ;
      LAYER met4 ;
        RECT 18.375 60.710 18.695 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 60.300 18.695 60.620 ;
      LAYER met4 ;
        RECT 18.375 60.300 18.695 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 59.890 18.695 60.210 ;
      LAYER met4 ;
        RECT 18.375 59.890 18.695 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 59.480 18.695 59.800 ;
      LAYER met4 ;
        RECT 18.375 59.480 18.695 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 59.070 18.695 59.390 ;
      LAYER met4 ;
        RECT 18.375 59.070 18.695 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 58.660 18.695 58.980 ;
      LAYER met4 ;
        RECT 18.375 58.660 18.695 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.375 58.250 18.695 58.570 ;
      LAYER met4 ;
        RECT 18.375 58.250 18.695 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 62.350 18.290 62.670 ;
      LAYER met4 ;
        RECT 17.970 62.350 18.290 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 61.940 18.290 62.260 ;
      LAYER met4 ;
        RECT 17.970 61.940 18.290 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 61.530 18.290 61.850 ;
      LAYER met4 ;
        RECT 17.970 61.530 18.290 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 61.120 18.290 61.440 ;
      LAYER met4 ;
        RECT 17.970 61.120 18.290 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 60.710 18.290 61.030 ;
      LAYER met4 ;
        RECT 17.970 60.710 18.290 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 60.300 18.290 60.620 ;
      LAYER met4 ;
        RECT 17.970 60.300 18.290 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 59.890 18.290 60.210 ;
      LAYER met4 ;
        RECT 17.970 59.890 18.290 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 59.480 18.290 59.800 ;
      LAYER met4 ;
        RECT 17.970 59.480 18.290 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 59.070 18.290 59.390 ;
      LAYER met4 ;
        RECT 17.970 59.070 18.290 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 58.660 18.290 58.980 ;
      LAYER met4 ;
        RECT 17.970 58.660 18.290 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.970 58.250 18.290 58.570 ;
      LAYER met4 ;
        RECT 17.970 58.250 18.290 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 62.350 17.885 62.670 ;
      LAYER met4 ;
        RECT 17.565 62.350 17.885 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 61.940 17.885 62.260 ;
      LAYER met4 ;
        RECT 17.565 61.940 17.885 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 61.530 17.885 61.850 ;
      LAYER met4 ;
        RECT 17.565 61.530 17.885 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 61.120 17.885 61.440 ;
      LAYER met4 ;
        RECT 17.565 61.120 17.885 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 60.710 17.885 61.030 ;
      LAYER met4 ;
        RECT 17.565 60.710 17.885 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 60.300 17.885 60.620 ;
      LAYER met4 ;
        RECT 17.565 60.300 17.885 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 59.890 17.885 60.210 ;
      LAYER met4 ;
        RECT 17.565 59.890 17.885 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 59.480 17.885 59.800 ;
      LAYER met4 ;
        RECT 17.565 59.480 17.885 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 59.070 17.885 59.390 ;
      LAYER met4 ;
        RECT 17.565 59.070 17.885 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 58.660 17.885 58.980 ;
      LAYER met4 ;
        RECT 17.565 58.660 17.885 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.565 58.250 17.885 58.570 ;
      LAYER met4 ;
        RECT 17.565 58.250 17.885 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 62.350 17.480 62.670 ;
      LAYER met4 ;
        RECT 17.160 62.350 17.480 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 61.940 17.480 62.260 ;
      LAYER met4 ;
        RECT 17.160 61.940 17.480 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 61.530 17.480 61.850 ;
      LAYER met4 ;
        RECT 17.160 61.530 17.480 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 61.120 17.480 61.440 ;
      LAYER met4 ;
        RECT 17.160 61.120 17.480 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 60.710 17.480 61.030 ;
      LAYER met4 ;
        RECT 17.160 60.710 17.480 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 60.300 17.480 60.620 ;
      LAYER met4 ;
        RECT 17.160 60.300 17.480 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 59.890 17.480 60.210 ;
      LAYER met4 ;
        RECT 17.160 59.890 17.480 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 59.480 17.480 59.800 ;
      LAYER met4 ;
        RECT 17.160 59.480 17.480 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 59.070 17.480 59.390 ;
      LAYER met4 ;
        RECT 17.160 59.070 17.480 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 58.660 17.480 58.980 ;
      LAYER met4 ;
        RECT 17.160 58.660 17.480 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.160 58.250 17.480 58.570 ;
      LAYER met4 ;
        RECT 17.160 58.250 17.480 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 62.350 17.075 62.670 ;
      LAYER met4 ;
        RECT 16.755 62.350 17.075 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 61.940 17.075 62.260 ;
      LAYER met4 ;
        RECT 16.755 61.940 17.075 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 61.530 17.075 61.850 ;
      LAYER met4 ;
        RECT 16.755 61.530 17.075 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 61.120 17.075 61.440 ;
      LAYER met4 ;
        RECT 16.755 61.120 17.075 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 60.710 17.075 61.030 ;
      LAYER met4 ;
        RECT 16.755 60.710 17.075 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 60.300 17.075 60.620 ;
      LAYER met4 ;
        RECT 16.755 60.300 17.075 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 59.890 17.075 60.210 ;
      LAYER met4 ;
        RECT 16.755 59.890 17.075 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 59.480 17.075 59.800 ;
      LAYER met4 ;
        RECT 16.755 59.480 17.075 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 59.070 17.075 59.390 ;
      LAYER met4 ;
        RECT 16.755 59.070 17.075 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 58.660 17.075 58.980 ;
      LAYER met4 ;
        RECT 16.755 58.660 17.075 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.755 58.250 17.075 58.570 ;
      LAYER met4 ;
        RECT 16.755 58.250 17.075 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 62.350 16.670 62.670 ;
      LAYER met4 ;
        RECT 16.350 62.350 16.670 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 61.940 16.670 62.260 ;
      LAYER met4 ;
        RECT 16.350 61.940 16.670 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 61.530 16.670 61.850 ;
      LAYER met4 ;
        RECT 16.350 61.530 16.670 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 61.120 16.670 61.440 ;
      LAYER met4 ;
        RECT 16.350 61.120 16.670 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 60.710 16.670 61.030 ;
      LAYER met4 ;
        RECT 16.350 60.710 16.670 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 60.300 16.670 60.620 ;
      LAYER met4 ;
        RECT 16.350 60.300 16.670 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 59.890 16.670 60.210 ;
      LAYER met4 ;
        RECT 16.350 59.890 16.670 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 59.480 16.670 59.800 ;
      LAYER met4 ;
        RECT 16.350 59.480 16.670 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 59.070 16.670 59.390 ;
      LAYER met4 ;
        RECT 16.350 59.070 16.670 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 58.660 16.670 58.980 ;
      LAYER met4 ;
        RECT 16.350 58.660 16.670 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.350 58.250 16.670 58.570 ;
      LAYER met4 ;
        RECT 16.350 58.250 16.670 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 62.350 16.265 62.670 ;
      LAYER met4 ;
        RECT 15.945 62.350 16.265 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 61.940 16.265 62.260 ;
      LAYER met4 ;
        RECT 15.945 61.940 16.265 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 61.530 16.265 61.850 ;
      LAYER met4 ;
        RECT 15.945 61.530 16.265 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 61.120 16.265 61.440 ;
      LAYER met4 ;
        RECT 15.945 61.120 16.265 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 60.710 16.265 61.030 ;
      LAYER met4 ;
        RECT 15.945 60.710 16.265 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 60.300 16.265 60.620 ;
      LAYER met4 ;
        RECT 15.945 60.300 16.265 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 59.890 16.265 60.210 ;
      LAYER met4 ;
        RECT 15.945 59.890 16.265 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 59.480 16.265 59.800 ;
      LAYER met4 ;
        RECT 15.945 59.480 16.265 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 59.070 16.265 59.390 ;
      LAYER met4 ;
        RECT 15.945 59.070 16.265 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 58.660 16.265 58.980 ;
      LAYER met4 ;
        RECT 15.945 58.660 16.265 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 58.250 16.265 58.570 ;
      LAYER met4 ;
        RECT 15.945 58.250 16.265 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 62.350 15.860 62.670 ;
      LAYER met4 ;
        RECT 15.540 62.350 15.860 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 61.940 15.860 62.260 ;
      LAYER met4 ;
        RECT 15.540 61.940 15.860 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 61.530 15.860 61.850 ;
      LAYER met4 ;
        RECT 15.540 61.530 15.860 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 61.120 15.860 61.440 ;
      LAYER met4 ;
        RECT 15.540 61.120 15.860 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 60.710 15.860 61.030 ;
      LAYER met4 ;
        RECT 15.540 60.710 15.860 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 60.300 15.860 60.620 ;
      LAYER met4 ;
        RECT 15.540 60.300 15.860 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 59.890 15.860 60.210 ;
      LAYER met4 ;
        RECT 15.540 59.890 15.860 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 59.480 15.860 59.800 ;
      LAYER met4 ;
        RECT 15.540 59.480 15.860 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 59.070 15.860 59.390 ;
      LAYER met4 ;
        RECT 15.540 59.070 15.860 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 58.660 15.860 58.980 ;
      LAYER met4 ;
        RECT 15.540 58.660 15.860 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.540 58.250 15.860 58.570 ;
      LAYER met4 ;
        RECT 15.540 58.250 15.860 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 62.350 15.455 62.670 ;
      LAYER met4 ;
        RECT 15.135 62.350 15.455 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 61.940 15.455 62.260 ;
      LAYER met4 ;
        RECT 15.135 61.940 15.455 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 61.530 15.455 61.850 ;
      LAYER met4 ;
        RECT 15.135 61.530 15.455 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 61.120 15.455 61.440 ;
      LAYER met4 ;
        RECT 15.135 61.120 15.455 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 60.710 15.455 61.030 ;
      LAYER met4 ;
        RECT 15.135 60.710 15.455 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 60.300 15.455 60.620 ;
      LAYER met4 ;
        RECT 15.135 60.300 15.455 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 59.890 15.455 60.210 ;
      LAYER met4 ;
        RECT 15.135 59.890 15.455 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 59.480 15.455 59.800 ;
      LAYER met4 ;
        RECT 15.135 59.480 15.455 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 59.070 15.455 59.390 ;
      LAYER met4 ;
        RECT 15.135 59.070 15.455 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 58.660 15.455 58.980 ;
      LAYER met4 ;
        RECT 15.135 58.660 15.455 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.135 58.250 15.455 58.570 ;
      LAYER met4 ;
        RECT 15.135 58.250 15.455 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 62.350 15.050 62.670 ;
      LAYER met4 ;
        RECT 14.730 62.350 15.050 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 61.940 15.050 62.260 ;
      LAYER met4 ;
        RECT 14.730 61.940 15.050 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 61.530 15.050 61.850 ;
      LAYER met4 ;
        RECT 14.730 61.530 15.050 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 61.120 15.050 61.440 ;
      LAYER met4 ;
        RECT 14.730 61.120 15.050 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 60.710 15.050 61.030 ;
      LAYER met4 ;
        RECT 14.730 60.710 15.050 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 60.300 15.050 60.620 ;
      LAYER met4 ;
        RECT 14.730 60.300 15.050 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 59.890 15.050 60.210 ;
      LAYER met4 ;
        RECT 14.730 59.890 15.050 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 59.480 15.050 59.800 ;
      LAYER met4 ;
        RECT 14.730 59.480 15.050 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 59.070 15.050 59.390 ;
      LAYER met4 ;
        RECT 14.730 59.070 15.050 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 58.660 15.050 58.980 ;
      LAYER met4 ;
        RECT 14.730 58.660 15.050 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.730 58.250 15.050 58.570 ;
      LAYER met4 ;
        RECT 14.730 58.250 15.050 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 62.350 14.645 62.670 ;
      LAYER met4 ;
        RECT 14.325 62.350 14.645 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 61.940 14.645 62.260 ;
      LAYER met4 ;
        RECT 14.325 61.940 14.645 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 61.530 14.645 61.850 ;
      LAYER met4 ;
        RECT 14.325 61.530 14.645 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 61.120 14.645 61.440 ;
      LAYER met4 ;
        RECT 14.325 61.120 14.645 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 60.710 14.645 61.030 ;
      LAYER met4 ;
        RECT 14.325 60.710 14.645 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 60.300 14.645 60.620 ;
      LAYER met4 ;
        RECT 14.325 60.300 14.645 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 59.890 14.645 60.210 ;
      LAYER met4 ;
        RECT 14.325 59.890 14.645 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 59.480 14.645 59.800 ;
      LAYER met4 ;
        RECT 14.325 59.480 14.645 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 59.070 14.645 59.390 ;
      LAYER met4 ;
        RECT 14.325 59.070 14.645 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 58.660 14.645 58.980 ;
      LAYER met4 ;
        RECT 14.325 58.660 14.645 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.325 58.250 14.645 58.570 ;
      LAYER met4 ;
        RECT 14.325 58.250 14.645 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 62.350 14.240 62.670 ;
      LAYER met4 ;
        RECT 13.920 62.350 14.240 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 61.940 14.240 62.260 ;
      LAYER met4 ;
        RECT 13.920 61.940 14.240 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 61.530 14.240 61.850 ;
      LAYER met4 ;
        RECT 13.920 61.530 14.240 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 61.120 14.240 61.440 ;
      LAYER met4 ;
        RECT 13.920 61.120 14.240 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 60.710 14.240 61.030 ;
      LAYER met4 ;
        RECT 13.920 60.710 14.240 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 60.300 14.240 60.620 ;
      LAYER met4 ;
        RECT 13.920 60.300 14.240 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 59.890 14.240 60.210 ;
      LAYER met4 ;
        RECT 13.920 59.890 14.240 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 59.480 14.240 59.800 ;
      LAYER met4 ;
        RECT 13.920 59.480 14.240 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 59.070 14.240 59.390 ;
      LAYER met4 ;
        RECT 13.920 59.070 14.240 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 58.660 14.240 58.980 ;
      LAYER met4 ;
        RECT 13.920 58.660 14.240 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.920 58.250 14.240 58.570 ;
      LAYER met4 ;
        RECT 13.920 58.250 14.240 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 62.350 13.835 62.670 ;
      LAYER met4 ;
        RECT 13.515 62.350 13.835 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 61.940 13.835 62.260 ;
      LAYER met4 ;
        RECT 13.515 61.940 13.835 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 61.530 13.835 61.850 ;
      LAYER met4 ;
        RECT 13.515 61.530 13.835 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 61.120 13.835 61.440 ;
      LAYER met4 ;
        RECT 13.515 61.120 13.835 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 60.710 13.835 61.030 ;
      LAYER met4 ;
        RECT 13.515 60.710 13.835 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 60.300 13.835 60.620 ;
      LAYER met4 ;
        RECT 13.515 60.300 13.835 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 59.890 13.835 60.210 ;
      LAYER met4 ;
        RECT 13.515 59.890 13.835 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 59.480 13.835 59.800 ;
      LAYER met4 ;
        RECT 13.515 59.480 13.835 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 59.070 13.835 59.390 ;
      LAYER met4 ;
        RECT 13.515 59.070 13.835 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 58.660 13.835 58.980 ;
      LAYER met4 ;
        RECT 13.515 58.660 13.835 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.515 58.250 13.835 58.570 ;
      LAYER met4 ;
        RECT 13.515 58.250 13.835 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 62.350 13.430 62.670 ;
      LAYER met4 ;
        RECT 13.110 62.350 13.430 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 61.940 13.430 62.260 ;
      LAYER met4 ;
        RECT 13.110 61.940 13.430 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 61.530 13.430 61.850 ;
      LAYER met4 ;
        RECT 13.110 61.530 13.430 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 61.120 13.430 61.440 ;
      LAYER met4 ;
        RECT 13.110 61.120 13.430 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 60.710 13.430 61.030 ;
      LAYER met4 ;
        RECT 13.110 60.710 13.430 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 60.300 13.430 60.620 ;
      LAYER met4 ;
        RECT 13.110 60.300 13.430 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 59.890 13.430 60.210 ;
      LAYER met4 ;
        RECT 13.110 59.890 13.430 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 59.480 13.430 59.800 ;
      LAYER met4 ;
        RECT 13.110 59.480 13.430 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 59.070 13.430 59.390 ;
      LAYER met4 ;
        RECT 13.110 59.070 13.430 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 58.660 13.430 58.980 ;
      LAYER met4 ;
        RECT 13.110 58.660 13.430 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.110 58.250 13.430 58.570 ;
      LAYER met4 ;
        RECT 13.110 58.250 13.430 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 62.350 13.025 62.670 ;
      LAYER met4 ;
        RECT 12.705 62.350 13.025 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 61.940 13.025 62.260 ;
      LAYER met4 ;
        RECT 12.705 61.940 13.025 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 61.530 13.025 61.850 ;
      LAYER met4 ;
        RECT 12.705 61.530 13.025 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 61.120 13.025 61.440 ;
      LAYER met4 ;
        RECT 12.705 61.120 13.025 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 60.710 13.025 61.030 ;
      LAYER met4 ;
        RECT 12.705 60.710 13.025 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 60.300 13.025 60.620 ;
      LAYER met4 ;
        RECT 12.705 60.300 13.025 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 59.890 13.025 60.210 ;
      LAYER met4 ;
        RECT 12.705 59.890 13.025 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 59.480 13.025 59.800 ;
      LAYER met4 ;
        RECT 12.705 59.480 13.025 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 59.070 13.025 59.390 ;
      LAYER met4 ;
        RECT 12.705 59.070 13.025 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 58.660 13.025 58.980 ;
      LAYER met4 ;
        RECT 12.705 58.660 13.025 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.705 58.250 13.025 58.570 ;
      LAYER met4 ;
        RECT 12.705 58.250 13.025 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 62.350 12.620 62.670 ;
      LAYER met4 ;
        RECT 12.300 62.350 12.620 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 61.940 12.620 62.260 ;
      LAYER met4 ;
        RECT 12.300 61.940 12.620 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 61.530 12.620 61.850 ;
      LAYER met4 ;
        RECT 12.300 61.530 12.620 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 61.120 12.620 61.440 ;
      LAYER met4 ;
        RECT 12.300 61.120 12.620 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 60.710 12.620 61.030 ;
      LAYER met4 ;
        RECT 12.300 60.710 12.620 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 60.300 12.620 60.620 ;
      LAYER met4 ;
        RECT 12.300 60.300 12.620 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 59.890 12.620 60.210 ;
      LAYER met4 ;
        RECT 12.300 59.890 12.620 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 59.480 12.620 59.800 ;
      LAYER met4 ;
        RECT 12.300 59.480 12.620 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 59.070 12.620 59.390 ;
      LAYER met4 ;
        RECT 12.300 59.070 12.620 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 58.660 12.620 58.980 ;
      LAYER met4 ;
        RECT 12.300 58.660 12.620 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.300 58.250 12.620 58.570 ;
      LAYER met4 ;
        RECT 12.300 58.250 12.620 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 62.350 12.215 62.670 ;
      LAYER met4 ;
        RECT 11.895 62.350 12.215 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 61.940 12.215 62.260 ;
      LAYER met4 ;
        RECT 11.895 61.940 12.215 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 61.530 12.215 61.850 ;
      LAYER met4 ;
        RECT 11.895 61.530 12.215 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 61.120 12.215 61.440 ;
      LAYER met4 ;
        RECT 11.895 61.120 12.215 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 60.710 12.215 61.030 ;
      LAYER met4 ;
        RECT 11.895 60.710 12.215 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 60.300 12.215 60.620 ;
      LAYER met4 ;
        RECT 11.895 60.300 12.215 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 59.890 12.215 60.210 ;
      LAYER met4 ;
        RECT 11.895 59.890 12.215 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 59.480 12.215 59.800 ;
      LAYER met4 ;
        RECT 11.895 59.480 12.215 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 59.070 12.215 59.390 ;
      LAYER met4 ;
        RECT 11.895 59.070 12.215 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 58.660 12.215 58.980 ;
      LAYER met4 ;
        RECT 11.895 58.660 12.215 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.895 58.250 12.215 58.570 ;
      LAYER met4 ;
        RECT 11.895 58.250 12.215 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 62.350 11.810 62.670 ;
      LAYER met4 ;
        RECT 11.490 62.350 11.810 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 61.940 11.810 62.260 ;
      LAYER met4 ;
        RECT 11.490 61.940 11.810 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 61.530 11.810 61.850 ;
      LAYER met4 ;
        RECT 11.490 61.530 11.810 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 61.120 11.810 61.440 ;
      LAYER met4 ;
        RECT 11.490 61.120 11.810 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 60.710 11.810 61.030 ;
      LAYER met4 ;
        RECT 11.490 60.710 11.810 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 60.300 11.810 60.620 ;
      LAYER met4 ;
        RECT 11.490 60.300 11.810 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 59.890 11.810 60.210 ;
      LAYER met4 ;
        RECT 11.490 59.890 11.810 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 59.480 11.810 59.800 ;
      LAYER met4 ;
        RECT 11.490 59.480 11.810 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 59.070 11.810 59.390 ;
      LAYER met4 ;
        RECT 11.490 59.070 11.810 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 58.660 11.810 58.980 ;
      LAYER met4 ;
        RECT 11.490 58.660 11.810 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.490 58.250 11.810 58.570 ;
      LAYER met4 ;
        RECT 11.490 58.250 11.810 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 62.350 11.405 62.670 ;
      LAYER met4 ;
        RECT 11.085 62.350 11.405 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 61.940 11.405 62.260 ;
      LAYER met4 ;
        RECT 11.085 61.940 11.405 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 61.530 11.405 61.850 ;
      LAYER met4 ;
        RECT 11.085 61.530 11.405 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 61.120 11.405 61.440 ;
      LAYER met4 ;
        RECT 11.085 61.120 11.405 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 60.710 11.405 61.030 ;
      LAYER met4 ;
        RECT 11.085 60.710 11.405 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 60.300 11.405 60.620 ;
      LAYER met4 ;
        RECT 11.085 60.300 11.405 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 59.890 11.405 60.210 ;
      LAYER met4 ;
        RECT 11.085 59.890 11.405 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 59.480 11.405 59.800 ;
      LAYER met4 ;
        RECT 11.085 59.480 11.405 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 59.070 11.405 59.390 ;
      LAYER met4 ;
        RECT 11.085 59.070 11.405 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 58.660 11.405 58.980 ;
      LAYER met4 ;
        RECT 11.085 58.660 11.405 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.085 58.250 11.405 58.570 ;
      LAYER met4 ;
        RECT 11.085 58.250 11.405 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 62.350 11.000 62.670 ;
      LAYER met4 ;
        RECT 10.680 62.350 11.000 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 61.940 11.000 62.260 ;
      LAYER met4 ;
        RECT 10.680 61.940 11.000 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 61.530 11.000 61.850 ;
      LAYER met4 ;
        RECT 10.680 61.530 11.000 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 61.120 11.000 61.440 ;
      LAYER met4 ;
        RECT 10.680 61.120 11.000 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 60.710 11.000 61.030 ;
      LAYER met4 ;
        RECT 10.680 60.710 11.000 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 60.300 11.000 60.620 ;
      LAYER met4 ;
        RECT 10.680 60.300 11.000 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 59.890 11.000 60.210 ;
      LAYER met4 ;
        RECT 10.680 59.890 11.000 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 59.480 11.000 59.800 ;
      LAYER met4 ;
        RECT 10.680 59.480 11.000 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 59.070 11.000 59.390 ;
      LAYER met4 ;
        RECT 10.680 59.070 11.000 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 58.660 11.000 58.980 ;
      LAYER met4 ;
        RECT 10.680 58.660 11.000 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.680 58.250 11.000 58.570 ;
      LAYER met4 ;
        RECT 10.680 58.250 11.000 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 62.350 10.595 62.670 ;
      LAYER met4 ;
        RECT 10.275 62.350 10.595 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 61.940 10.595 62.260 ;
      LAYER met4 ;
        RECT 10.275 61.940 10.595 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 61.530 10.595 61.850 ;
      LAYER met4 ;
        RECT 10.275 61.530 10.595 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 61.120 10.595 61.440 ;
      LAYER met4 ;
        RECT 10.275 61.120 10.595 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 60.710 10.595 61.030 ;
      LAYER met4 ;
        RECT 10.275 60.710 10.595 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 60.300 10.595 60.620 ;
      LAYER met4 ;
        RECT 10.275 60.300 10.595 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 59.890 10.595 60.210 ;
      LAYER met4 ;
        RECT 10.275 59.890 10.595 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 59.480 10.595 59.800 ;
      LAYER met4 ;
        RECT 10.275 59.480 10.595 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 59.070 10.595 59.390 ;
      LAYER met4 ;
        RECT 10.275 59.070 10.595 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 58.660 10.595 58.980 ;
      LAYER met4 ;
        RECT 10.275 58.660 10.595 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.275 58.250 10.595 58.570 ;
      LAYER met4 ;
        RECT 10.275 58.250 10.595 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 62.350 10.190 62.670 ;
      LAYER met4 ;
        RECT 9.870 62.350 10.190 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 61.940 10.190 62.260 ;
      LAYER met4 ;
        RECT 9.870 61.940 10.190 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 61.530 10.190 61.850 ;
      LAYER met4 ;
        RECT 9.870 61.530 10.190 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 61.120 10.190 61.440 ;
      LAYER met4 ;
        RECT 9.870 61.120 10.190 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 60.710 10.190 61.030 ;
      LAYER met4 ;
        RECT 9.870 60.710 10.190 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 60.300 10.190 60.620 ;
      LAYER met4 ;
        RECT 9.870 60.300 10.190 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 59.890 10.190 60.210 ;
      LAYER met4 ;
        RECT 9.870 59.890 10.190 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 59.480 10.190 59.800 ;
      LAYER met4 ;
        RECT 9.870 59.480 10.190 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 59.070 10.190 59.390 ;
      LAYER met4 ;
        RECT 9.870 59.070 10.190 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 58.660 10.190 58.980 ;
      LAYER met4 ;
        RECT 9.870 58.660 10.190 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.870 58.250 10.190 58.570 ;
      LAYER met4 ;
        RECT 9.870 58.250 10.190 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 62.350 9.785 62.670 ;
      LAYER met4 ;
        RECT 9.465 62.350 9.785 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 61.940 9.785 62.260 ;
      LAYER met4 ;
        RECT 9.465 61.940 9.785 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 61.530 9.785 61.850 ;
      LAYER met4 ;
        RECT 9.465 61.530 9.785 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 61.120 9.785 61.440 ;
      LAYER met4 ;
        RECT 9.465 61.120 9.785 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 60.710 9.785 61.030 ;
      LAYER met4 ;
        RECT 9.465 60.710 9.785 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 60.300 9.785 60.620 ;
      LAYER met4 ;
        RECT 9.465 60.300 9.785 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 59.890 9.785 60.210 ;
      LAYER met4 ;
        RECT 9.465 59.890 9.785 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 59.480 9.785 59.800 ;
      LAYER met4 ;
        RECT 9.465 59.480 9.785 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 59.070 9.785 59.390 ;
      LAYER met4 ;
        RECT 9.465 59.070 9.785 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 58.660 9.785 58.980 ;
      LAYER met4 ;
        RECT 9.465 58.660 9.785 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.465 58.250 9.785 58.570 ;
      LAYER met4 ;
        RECT 9.465 58.250 9.785 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 62.350 9.380 62.670 ;
      LAYER met4 ;
        RECT 9.060 62.350 9.380 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 61.940 9.380 62.260 ;
      LAYER met4 ;
        RECT 9.060 61.940 9.380 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 61.530 9.380 61.850 ;
      LAYER met4 ;
        RECT 9.060 61.530 9.380 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 61.120 9.380 61.440 ;
      LAYER met4 ;
        RECT 9.060 61.120 9.380 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 60.710 9.380 61.030 ;
      LAYER met4 ;
        RECT 9.060 60.710 9.380 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 60.300 9.380 60.620 ;
      LAYER met4 ;
        RECT 9.060 60.300 9.380 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 59.890 9.380 60.210 ;
      LAYER met4 ;
        RECT 9.060 59.890 9.380 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 59.480 9.380 59.800 ;
      LAYER met4 ;
        RECT 9.060 59.480 9.380 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 59.070 9.380 59.390 ;
      LAYER met4 ;
        RECT 9.060 59.070 9.380 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 58.660 9.380 58.980 ;
      LAYER met4 ;
        RECT 9.060 58.660 9.380 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.060 58.250 9.380 58.570 ;
      LAYER met4 ;
        RECT 9.060 58.250 9.380 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 62.350 8.975 62.670 ;
      LAYER met4 ;
        RECT 8.655 62.350 8.975 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 61.940 8.975 62.260 ;
      LAYER met4 ;
        RECT 8.655 61.940 8.975 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 61.530 8.975 61.850 ;
      LAYER met4 ;
        RECT 8.655 61.530 8.975 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 61.120 8.975 61.440 ;
      LAYER met4 ;
        RECT 8.655 61.120 8.975 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 60.710 8.975 61.030 ;
      LAYER met4 ;
        RECT 8.655 60.710 8.975 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 60.300 8.975 60.620 ;
      LAYER met4 ;
        RECT 8.655 60.300 8.975 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 59.890 8.975 60.210 ;
      LAYER met4 ;
        RECT 8.655 59.890 8.975 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 59.480 8.975 59.800 ;
      LAYER met4 ;
        RECT 8.655 59.480 8.975 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 59.070 8.975 59.390 ;
      LAYER met4 ;
        RECT 8.655 59.070 8.975 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 58.660 8.975 58.980 ;
      LAYER met4 ;
        RECT 8.655 58.660 8.975 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.655 58.250 8.975 58.570 ;
      LAYER met4 ;
        RECT 8.655 58.250 8.975 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 62.350 8.570 62.670 ;
      LAYER met4 ;
        RECT 8.250 62.350 8.570 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 61.940 8.570 62.260 ;
      LAYER met4 ;
        RECT 8.250 61.940 8.570 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 61.530 8.570 61.850 ;
      LAYER met4 ;
        RECT 8.250 61.530 8.570 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 61.120 8.570 61.440 ;
      LAYER met4 ;
        RECT 8.250 61.120 8.570 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 60.710 8.570 61.030 ;
      LAYER met4 ;
        RECT 8.250 60.710 8.570 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 60.300 8.570 60.620 ;
      LAYER met4 ;
        RECT 8.250 60.300 8.570 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 59.890 8.570 60.210 ;
      LAYER met4 ;
        RECT 8.250 59.890 8.570 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 59.480 8.570 59.800 ;
      LAYER met4 ;
        RECT 8.250 59.480 8.570 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 59.070 8.570 59.390 ;
      LAYER met4 ;
        RECT 8.250 59.070 8.570 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 58.660 8.570 58.980 ;
      LAYER met4 ;
        RECT 8.250 58.660 8.570 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.250 58.250 8.570 58.570 ;
      LAYER met4 ;
        RECT 8.250 58.250 8.570 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 62.350 8.165 62.670 ;
      LAYER met4 ;
        RECT 7.845 62.350 8.165 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 61.940 8.165 62.260 ;
      LAYER met4 ;
        RECT 7.845 61.940 8.165 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 61.530 8.165 61.850 ;
      LAYER met4 ;
        RECT 7.845 61.530 8.165 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 61.120 8.165 61.440 ;
      LAYER met4 ;
        RECT 7.845 61.120 8.165 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 60.710 8.165 61.030 ;
      LAYER met4 ;
        RECT 7.845 60.710 8.165 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 60.300 8.165 60.620 ;
      LAYER met4 ;
        RECT 7.845 60.300 8.165 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 59.890 8.165 60.210 ;
      LAYER met4 ;
        RECT 7.845 59.890 8.165 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 59.480 8.165 59.800 ;
      LAYER met4 ;
        RECT 7.845 59.480 8.165 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 59.070 8.165 59.390 ;
      LAYER met4 ;
        RECT 7.845 59.070 8.165 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 58.660 8.165 58.980 ;
      LAYER met4 ;
        RECT 7.845 58.660 8.165 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.845 58.250 8.165 58.570 ;
      LAYER met4 ;
        RECT 7.845 58.250 8.165 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 62.350 7.760 62.670 ;
      LAYER met4 ;
        RECT 7.440 62.350 7.760 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 61.940 7.760 62.260 ;
      LAYER met4 ;
        RECT 7.440 61.940 7.760 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 61.530 7.760 61.850 ;
      LAYER met4 ;
        RECT 7.440 61.530 7.760 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 61.120 7.760 61.440 ;
      LAYER met4 ;
        RECT 7.440 61.120 7.760 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 60.710 7.760 61.030 ;
      LAYER met4 ;
        RECT 7.440 60.710 7.760 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 60.300 7.760 60.620 ;
      LAYER met4 ;
        RECT 7.440 60.300 7.760 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 59.890 7.760 60.210 ;
      LAYER met4 ;
        RECT 7.440 59.890 7.760 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 59.480 7.760 59.800 ;
      LAYER met4 ;
        RECT 7.440 59.480 7.760 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 59.070 7.760 59.390 ;
      LAYER met4 ;
        RECT 7.440 59.070 7.760 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 58.660 7.760 58.980 ;
      LAYER met4 ;
        RECT 7.440 58.660 7.760 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.440 58.250 7.760 58.570 ;
      LAYER met4 ;
        RECT 7.440 58.250 7.760 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 62.350 7.355 62.670 ;
      LAYER met4 ;
        RECT 7.035 62.350 7.355 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 61.940 7.355 62.260 ;
      LAYER met4 ;
        RECT 7.035 61.940 7.355 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 61.530 7.355 61.850 ;
      LAYER met4 ;
        RECT 7.035 61.530 7.355 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 61.120 7.355 61.440 ;
      LAYER met4 ;
        RECT 7.035 61.120 7.355 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 60.710 7.355 61.030 ;
      LAYER met4 ;
        RECT 7.035 60.710 7.355 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 60.300 7.355 60.620 ;
      LAYER met4 ;
        RECT 7.035 60.300 7.355 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 59.890 7.355 60.210 ;
      LAYER met4 ;
        RECT 7.035 59.890 7.355 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 59.480 7.355 59.800 ;
      LAYER met4 ;
        RECT 7.035 59.480 7.355 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 59.070 7.355 59.390 ;
      LAYER met4 ;
        RECT 7.035 59.070 7.355 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 58.660 7.355 58.980 ;
      LAYER met4 ;
        RECT 7.035 58.660 7.355 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.035 58.250 7.355 58.570 ;
      LAYER met4 ;
        RECT 7.035 58.250 7.355 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 62.350 6.950 62.670 ;
      LAYER met4 ;
        RECT 6.630 62.350 6.950 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 61.940 6.950 62.260 ;
      LAYER met4 ;
        RECT 6.630 61.940 6.950 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 61.530 6.950 61.850 ;
      LAYER met4 ;
        RECT 6.630 61.530 6.950 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 61.120 6.950 61.440 ;
      LAYER met4 ;
        RECT 6.630 61.120 6.950 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 60.710 6.950 61.030 ;
      LAYER met4 ;
        RECT 6.630 60.710 6.950 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 60.300 6.950 60.620 ;
      LAYER met4 ;
        RECT 6.630 60.300 6.950 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 59.890 6.950 60.210 ;
      LAYER met4 ;
        RECT 6.630 59.890 6.950 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 59.480 6.950 59.800 ;
      LAYER met4 ;
        RECT 6.630 59.480 6.950 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 59.070 6.950 59.390 ;
      LAYER met4 ;
        RECT 6.630 59.070 6.950 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 58.660 6.950 58.980 ;
      LAYER met4 ;
        RECT 6.630 58.660 6.950 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.630 58.250 6.950 58.570 ;
      LAYER met4 ;
        RECT 6.630 58.250 6.950 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 62.350 6.545 62.670 ;
      LAYER met4 ;
        RECT 6.225 62.350 6.545 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 61.940 6.545 62.260 ;
      LAYER met4 ;
        RECT 6.225 61.940 6.545 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 61.530 6.545 61.850 ;
      LAYER met4 ;
        RECT 6.225 61.530 6.545 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 61.120 6.545 61.440 ;
      LAYER met4 ;
        RECT 6.225 61.120 6.545 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 60.710 6.545 61.030 ;
      LAYER met4 ;
        RECT 6.225 60.710 6.545 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 60.300 6.545 60.620 ;
      LAYER met4 ;
        RECT 6.225 60.300 6.545 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 59.890 6.545 60.210 ;
      LAYER met4 ;
        RECT 6.225 59.890 6.545 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 59.480 6.545 59.800 ;
      LAYER met4 ;
        RECT 6.225 59.480 6.545 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 59.070 6.545 59.390 ;
      LAYER met4 ;
        RECT 6.225 59.070 6.545 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 58.660 6.545 58.980 ;
      LAYER met4 ;
        RECT 6.225 58.660 6.545 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.225 58.250 6.545 58.570 ;
      LAYER met4 ;
        RECT 6.225 58.250 6.545 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 62.350 6.140 62.670 ;
      LAYER met4 ;
        RECT 5.820 62.350 6.140 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 61.940 6.140 62.260 ;
      LAYER met4 ;
        RECT 5.820 61.940 6.140 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 61.530 6.140 61.850 ;
      LAYER met4 ;
        RECT 5.820 61.530 6.140 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 61.120 6.140 61.440 ;
      LAYER met4 ;
        RECT 5.820 61.120 6.140 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 60.710 6.140 61.030 ;
      LAYER met4 ;
        RECT 5.820 60.710 6.140 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 60.300 6.140 60.620 ;
      LAYER met4 ;
        RECT 5.820 60.300 6.140 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 59.890 6.140 60.210 ;
      LAYER met4 ;
        RECT 5.820 59.890 6.140 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 59.480 6.140 59.800 ;
      LAYER met4 ;
        RECT 5.820 59.480 6.140 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 59.070 6.140 59.390 ;
      LAYER met4 ;
        RECT 5.820 59.070 6.140 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 58.660 6.140 58.980 ;
      LAYER met4 ;
        RECT 5.820 58.660 6.140 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.820 58.250 6.140 58.570 ;
      LAYER met4 ;
        RECT 5.820 58.250 6.140 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 62.350 5.735 62.670 ;
      LAYER met4 ;
        RECT 5.415 62.350 5.735 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 61.940 5.735 62.260 ;
      LAYER met4 ;
        RECT 5.415 61.940 5.735 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 61.530 5.735 61.850 ;
      LAYER met4 ;
        RECT 5.415 61.530 5.735 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 61.120 5.735 61.440 ;
      LAYER met4 ;
        RECT 5.415 61.120 5.735 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 60.710 5.735 61.030 ;
      LAYER met4 ;
        RECT 5.415 60.710 5.735 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 60.300 5.735 60.620 ;
      LAYER met4 ;
        RECT 5.415 60.300 5.735 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 59.890 5.735 60.210 ;
      LAYER met4 ;
        RECT 5.415 59.890 5.735 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 59.480 5.735 59.800 ;
      LAYER met4 ;
        RECT 5.415 59.480 5.735 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 59.070 5.735 59.390 ;
      LAYER met4 ;
        RECT 5.415 59.070 5.735 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 58.660 5.735 58.980 ;
      LAYER met4 ;
        RECT 5.415 58.660 5.735 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.415 58.250 5.735 58.570 ;
      LAYER met4 ;
        RECT 5.415 58.250 5.735 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 62.350 5.330 62.670 ;
      LAYER met4 ;
        RECT 5.010 62.350 5.330 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 61.940 5.330 62.260 ;
      LAYER met4 ;
        RECT 5.010 61.940 5.330 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 61.530 5.330 61.850 ;
      LAYER met4 ;
        RECT 5.010 61.530 5.330 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 61.120 5.330 61.440 ;
      LAYER met4 ;
        RECT 5.010 61.120 5.330 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 60.710 5.330 61.030 ;
      LAYER met4 ;
        RECT 5.010 60.710 5.330 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 60.300 5.330 60.620 ;
      LAYER met4 ;
        RECT 5.010 60.300 5.330 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 59.890 5.330 60.210 ;
      LAYER met4 ;
        RECT 5.010 59.890 5.330 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 59.480 5.330 59.800 ;
      LAYER met4 ;
        RECT 5.010 59.480 5.330 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 59.070 5.330 59.390 ;
      LAYER met4 ;
        RECT 5.010 59.070 5.330 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 58.660 5.330 58.980 ;
      LAYER met4 ;
        RECT 5.010 58.660 5.330 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.010 58.250 5.330 58.570 ;
      LAYER met4 ;
        RECT 5.010 58.250 5.330 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 62.350 4.925 62.670 ;
      LAYER met4 ;
        RECT 4.605 62.350 4.925 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 61.940 4.925 62.260 ;
      LAYER met4 ;
        RECT 4.605 61.940 4.925 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 61.530 4.925 61.850 ;
      LAYER met4 ;
        RECT 4.605 61.530 4.925 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 61.120 4.925 61.440 ;
      LAYER met4 ;
        RECT 4.605 61.120 4.925 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 60.710 4.925 61.030 ;
      LAYER met4 ;
        RECT 4.605 60.710 4.925 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 60.300 4.925 60.620 ;
      LAYER met4 ;
        RECT 4.605 60.300 4.925 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 59.890 4.925 60.210 ;
      LAYER met4 ;
        RECT 4.605 59.890 4.925 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 59.480 4.925 59.800 ;
      LAYER met4 ;
        RECT 4.605 59.480 4.925 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 59.070 4.925 59.390 ;
      LAYER met4 ;
        RECT 4.605 59.070 4.925 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 58.660 4.925 58.980 ;
      LAYER met4 ;
        RECT 4.605 58.660 4.925 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.605 58.250 4.925 58.570 ;
      LAYER met4 ;
        RECT 4.605 58.250 4.925 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 62.350 4.520 62.670 ;
      LAYER met4 ;
        RECT 4.200 62.350 4.520 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 61.940 4.520 62.260 ;
      LAYER met4 ;
        RECT 4.200 61.940 4.520 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 61.530 4.520 61.850 ;
      LAYER met4 ;
        RECT 4.200 61.530 4.520 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 61.120 4.520 61.440 ;
      LAYER met4 ;
        RECT 4.200 61.120 4.520 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 60.710 4.520 61.030 ;
      LAYER met4 ;
        RECT 4.200 60.710 4.520 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 60.300 4.520 60.620 ;
      LAYER met4 ;
        RECT 4.200 60.300 4.520 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 59.890 4.520 60.210 ;
      LAYER met4 ;
        RECT 4.200 59.890 4.520 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 59.480 4.520 59.800 ;
      LAYER met4 ;
        RECT 4.200 59.480 4.520 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 59.070 4.520 59.390 ;
      LAYER met4 ;
        RECT 4.200 59.070 4.520 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 58.660 4.520 58.980 ;
      LAYER met4 ;
        RECT 4.200 58.660 4.520 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.200 58.250 4.520 58.570 ;
      LAYER met4 ;
        RECT 4.200 58.250 4.520 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 62.350 4.115 62.670 ;
      LAYER met4 ;
        RECT 3.795 62.350 4.115 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 61.940 4.115 62.260 ;
      LAYER met4 ;
        RECT 3.795 61.940 4.115 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 61.530 4.115 61.850 ;
      LAYER met4 ;
        RECT 3.795 61.530 4.115 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 61.120 4.115 61.440 ;
      LAYER met4 ;
        RECT 3.795 61.120 4.115 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 60.710 4.115 61.030 ;
      LAYER met4 ;
        RECT 3.795 60.710 4.115 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 60.300 4.115 60.620 ;
      LAYER met4 ;
        RECT 3.795 60.300 4.115 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 59.890 4.115 60.210 ;
      LAYER met4 ;
        RECT 3.795 59.890 4.115 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 59.480 4.115 59.800 ;
      LAYER met4 ;
        RECT 3.795 59.480 4.115 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 59.070 4.115 59.390 ;
      LAYER met4 ;
        RECT 3.795 59.070 4.115 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 58.660 4.115 58.980 ;
      LAYER met4 ;
        RECT 3.795 58.660 4.115 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.795 58.250 4.115 58.570 ;
      LAYER met4 ;
        RECT 3.795 58.250 4.115 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 62.350 3.710 62.670 ;
      LAYER met4 ;
        RECT 3.390 62.350 3.710 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 61.940 3.710 62.260 ;
      LAYER met4 ;
        RECT 3.390 61.940 3.710 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 61.530 3.710 61.850 ;
      LAYER met4 ;
        RECT 3.390 61.530 3.710 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 61.120 3.710 61.440 ;
      LAYER met4 ;
        RECT 3.390 61.120 3.710 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 60.710 3.710 61.030 ;
      LAYER met4 ;
        RECT 3.390 60.710 3.710 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 60.300 3.710 60.620 ;
      LAYER met4 ;
        RECT 3.390 60.300 3.710 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 59.890 3.710 60.210 ;
      LAYER met4 ;
        RECT 3.390 59.890 3.710 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 59.480 3.710 59.800 ;
      LAYER met4 ;
        RECT 3.390 59.480 3.710 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 59.070 3.710 59.390 ;
      LAYER met4 ;
        RECT 3.390 59.070 3.710 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 58.660 3.710 58.980 ;
      LAYER met4 ;
        RECT 3.390 58.660 3.710 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.390 58.250 3.710 58.570 ;
      LAYER met4 ;
        RECT 3.390 58.250 3.710 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 62.350 3.305 62.670 ;
      LAYER met4 ;
        RECT 2.985 62.350 3.305 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 61.940 3.305 62.260 ;
      LAYER met4 ;
        RECT 2.985 61.940 3.305 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 61.530 3.305 61.850 ;
      LAYER met4 ;
        RECT 2.985 61.530 3.305 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 61.120 3.305 61.440 ;
      LAYER met4 ;
        RECT 2.985 61.120 3.305 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 60.710 3.305 61.030 ;
      LAYER met4 ;
        RECT 2.985 60.710 3.305 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 60.300 3.305 60.620 ;
      LAYER met4 ;
        RECT 2.985 60.300 3.305 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 59.890 3.305 60.210 ;
      LAYER met4 ;
        RECT 2.985 59.890 3.305 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 59.480 3.305 59.800 ;
      LAYER met4 ;
        RECT 2.985 59.480 3.305 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 59.070 3.305 59.390 ;
      LAYER met4 ;
        RECT 2.985 59.070 3.305 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 58.660 3.305 58.980 ;
      LAYER met4 ;
        RECT 2.985 58.660 3.305 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.985 58.250 3.305 58.570 ;
      LAYER met4 ;
        RECT 2.985 58.250 3.305 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 62.350 2.895 62.670 ;
      LAYER met4 ;
        RECT 2.575 62.350 2.895 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 61.940 2.895 62.260 ;
      LAYER met4 ;
        RECT 2.575 61.940 2.895 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 61.530 2.895 61.850 ;
      LAYER met4 ;
        RECT 2.575 61.530 2.895 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 61.120 2.895 61.440 ;
      LAYER met4 ;
        RECT 2.575 61.120 2.895 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 60.710 2.895 61.030 ;
      LAYER met4 ;
        RECT 2.575 60.710 2.895 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 60.300 2.895 60.620 ;
      LAYER met4 ;
        RECT 2.575 60.300 2.895 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 59.890 2.895 60.210 ;
      LAYER met4 ;
        RECT 2.575 59.890 2.895 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 59.480 2.895 59.800 ;
      LAYER met4 ;
        RECT 2.575 59.480 2.895 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 59.070 2.895 59.390 ;
      LAYER met4 ;
        RECT 2.575 59.070 2.895 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 58.660 2.895 58.980 ;
      LAYER met4 ;
        RECT 2.575 58.660 2.895 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.575 58.250 2.895 58.570 ;
      LAYER met4 ;
        RECT 2.575 58.250 2.895 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 62.350 2.485 62.670 ;
      LAYER met4 ;
        RECT 2.165 62.350 2.485 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 61.940 2.485 62.260 ;
      LAYER met4 ;
        RECT 2.165 61.940 2.485 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 61.530 2.485 61.850 ;
      LAYER met4 ;
        RECT 2.165 61.530 2.485 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 61.120 2.485 61.440 ;
      LAYER met4 ;
        RECT 2.165 61.120 2.485 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 60.710 2.485 61.030 ;
      LAYER met4 ;
        RECT 2.165 60.710 2.485 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 60.300 2.485 60.620 ;
      LAYER met4 ;
        RECT 2.165 60.300 2.485 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 59.890 2.485 60.210 ;
      LAYER met4 ;
        RECT 2.165 59.890 2.485 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 59.480 2.485 59.800 ;
      LAYER met4 ;
        RECT 2.165 59.480 2.485 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 59.070 2.485 59.390 ;
      LAYER met4 ;
        RECT 2.165 59.070 2.485 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 58.660 2.485 58.980 ;
      LAYER met4 ;
        RECT 2.165 58.660 2.485 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.165 58.250 2.485 58.570 ;
      LAYER met4 ;
        RECT 2.165 58.250 2.485 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 62.350 2.075 62.670 ;
      LAYER met4 ;
        RECT 1.755 62.350 2.075 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 61.940 2.075 62.260 ;
      LAYER met4 ;
        RECT 1.755 61.940 2.075 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 61.530 2.075 61.850 ;
      LAYER met4 ;
        RECT 1.755 61.530 2.075 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 61.120 2.075 61.440 ;
      LAYER met4 ;
        RECT 1.755 61.120 2.075 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 60.710 2.075 61.030 ;
      LAYER met4 ;
        RECT 1.755 60.710 2.075 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 60.300 2.075 60.620 ;
      LAYER met4 ;
        RECT 1.755 60.300 2.075 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 59.890 2.075 60.210 ;
      LAYER met4 ;
        RECT 1.755 59.890 2.075 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 59.480 2.075 59.800 ;
      LAYER met4 ;
        RECT 1.755 59.480 2.075 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 59.070 2.075 59.390 ;
      LAYER met4 ;
        RECT 1.755 59.070 2.075 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 58.660 2.075 58.980 ;
      LAYER met4 ;
        RECT 1.755 58.660 2.075 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 58.250 2.075 58.570 ;
      LAYER met4 ;
        RECT 1.755 58.250 2.075 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 62.350 1.665 62.670 ;
      LAYER met4 ;
        RECT 1.345 62.350 1.665 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 61.940 1.665 62.260 ;
      LAYER met4 ;
        RECT 1.345 61.940 1.665 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 61.530 1.665 61.850 ;
      LAYER met4 ;
        RECT 1.345 61.530 1.665 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 61.120 1.665 61.440 ;
      LAYER met4 ;
        RECT 1.345 61.120 1.665 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 60.710 1.665 61.030 ;
      LAYER met4 ;
        RECT 1.345 60.710 1.665 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 60.300 1.665 60.620 ;
      LAYER met4 ;
        RECT 1.345 60.300 1.665 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 59.890 1.665 60.210 ;
      LAYER met4 ;
        RECT 1.345 59.890 1.665 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 59.480 1.665 59.800 ;
      LAYER met4 ;
        RECT 1.345 59.480 1.665 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 59.070 1.665 59.390 ;
      LAYER met4 ;
        RECT 1.345 59.070 1.665 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 58.660 1.665 58.980 ;
      LAYER met4 ;
        RECT 1.345 58.660 1.665 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.345 58.250 1.665 58.570 ;
      LAYER met4 ;
        RECT 1.345 58.250 1.665 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 62.350 1.255 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 61.940 1.255 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 61.530 1.255 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 61.120 1.255 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 60.710 1.255 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 60.300 1.255 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 59.890 1.255 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 59.480 1.255 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 59.070 1.255 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 58.660 1.255 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.935 58.250 1.255 58.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 62.350 0.845 62.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 61.940 0.845 62.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 61.530 0.845 61.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 61.120 0.845 61.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 60.710 0.845 61.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 60.300 0.845 60.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 59.890 0.845 60.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 59.480 0.845 59.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 59.070 0.845 59.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 58.660 0.845 58.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.525 58.250 0.845 58.570 ;
    END
  END VSSIO_Q
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
  END VCCHIB
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  OBS
      LAYER met3 ;
        RECT 0.495 58.240 74.290 200.000 ;
      LAYER met4 ;
        RECT 1.670 197.370 13.230 200.000 ;
        RECT 61.725 197.370 73.330 200.000 ;
        RECT 1.670 195.830 13.195 197.370 ;
        RECT 14.655 195.830 60.280 196.770 ;
        RECT 61.740 195.830 73.330 197.370 ;
        RECT 1.670 175.385 73.330 195.830 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 96.585 75.000 174.185 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__overlay_vssio_hvc

#--------EOF---------

MACRO sky130_fd_io__overlay_vssio_lvc
  CLASS PAD ;
  FOREIGN sky130_fd_io__overlay_vssio_lvc ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
  END VCCD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
  END VSSA
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
  END VDDA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 23.840 24.400 28.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 23.840 74.290 28.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.045 171.195 74.700 198.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 197.705 74.640 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 197.300 74.640 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 196.895 74.640 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 196.490 74.640 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 196.085 74.640 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 195.680 74.640 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 195.275 74.640 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 194.870 74.640 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 194.465 74.640 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 194.060 74.640 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 193.655 74.640 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 193.250 74.640 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 192.845 74.640 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 192.440 74.640 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 192.035 74.640 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 191.630 74.640 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 191.225 74.640 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 190.820 74.640 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 190.415 74.640 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 190.010 74.640 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 189.605 74.640 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 189.200 74.640 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 188.795 74.640 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 188.390 74.640 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 187.985 74.640 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 187.580 74.640 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 187.175 74.640 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 186.770 74.640 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 186.365 74.640 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 185.960 74.640 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 185.555 74.640 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 185.150 74.640 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 184.745 74.640 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 184.340 74.640 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 183.935 74.640 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 183.530 74.640 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 183.125 74.640 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 182.720 74.640 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 182.315 74.640 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 181.910 74.640 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 181.505 74.640 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 181.100 74.640 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 180.700 74.640 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 180.300 74.640 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 179.900 74.640 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 179.500 74.640 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 179.100 74.640 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 178.700 74.640 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 178.300 74.640 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 177.900 74.640 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 177.500 74.640 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 177.100 74.640 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 176.700 74.640 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 176.300 74.640 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 175.900 74.640 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 175.500 74.640 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 175.100 74.640 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 174.700 74.640 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 174.300 74.640 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.440 173.900 74.640 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 197.705 74.230 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 197.300 74.230 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 196.895 74.230 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 196.490 74.230 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 196.085 74.230 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 195.680 74.230 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 195.275 74.230 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 194.870 74.230 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 194.465 74.230 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 194.060 74.230 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 193.655 74.230 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 193.250 74.230 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 192.845 74.230 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 192.440 74.230 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 192.035 74.230 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 191.630 74.230 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 191.225 74.230 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 190.820 74.230 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 190.415 74.230 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 190.010 74.230 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 189.605 74.230 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 189.200 74.230 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 188.795 74.230 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 188.390 74.230 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 187.985 74.230 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 187.580 74.230 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 187.175 74.230 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 186.770 74.230 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 186.365 74.230 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 185.960 74.230 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 185.555 74.230 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 185.150 74.230 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 184.745 74.230 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 184.340 74.230 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 183.935 74.230 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 183.530 74.230 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 183.125 74.230 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 182.720 74.230 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 182.315 74.230 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 181.910 74.230 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 181.505 74.230 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 181.100 74.230 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 180.700 74.230 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 180.300 74.230 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 179.900 74.230 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 179.500 74.230 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 179.100 74.230 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 178.700 74.230 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 178.300 74.230 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 177.900 74.230 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 177.500 74.230 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 177.100 74.230 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 176.700 74.230 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 176.300 74.230 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 175.900 74.230 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 175.500 74.230 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 175.100 74.230 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 174.700 74.230 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 174.300 74.230 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.030 173.900 74.230 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 28.210 74.200 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 27.780 74.200 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 27.350 74.200 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 26.920 74.200 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 26.490 74.200 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 26.060 74.200 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 25.630 74.200 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 25.200 74.200 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 24.770 74.200 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 24.340 74.200 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 23.910 74.200 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 197.705 73.820 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 197.300 73.820 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 196.895 73.820 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 196.490 73.820 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 196.085 73.820 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 195.680 73.820 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 195.275 73.820 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 194.870 73.820 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 194.465 73.820 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 194.060 73.820 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 193.655 73.820 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 193.250 73.820 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 192.845 73.820 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 192.440 73.820 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 192.035 73.820 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 191.630 73.820 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 191.225 73.820 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 190.820 73.820 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 190.415 73.820 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 190.010 73.820 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 189.605 73.820 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 189.200 73.820 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 188.795 73.820 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 188.390 73.820 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 187.985 73.820 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 187.580 73.820 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 187.175 73.820 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 186.770 73.820 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 186.365 73.820 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 185.960 73.820 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 185.555 73.820 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 185.150 73.820 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 184.745 73.820 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 184.340 73.820 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 183.935 73.820 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 183.530 73.820 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 183.125 73.820 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 182.720 73.820 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 182.315 73.820 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 181.910 73.820 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 181.505 73.820 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 181.100 73.820 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 180.700 73.820 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 180.300 73.820 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 179.900 73.820 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 179.500 73.820 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 179.100 73.820 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 178.700 73.820 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 178.300 73.820 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 177.900 73.820 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 177.500 73.820 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 177.100 73.820 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 176.700 73.820 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 176.300 73.820 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 175.900 73.820 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 175.500 73.820 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 175.100 73.820 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 174.700 73.820 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 174.300 73.820 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.620 173.900 73.820 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 28.210 73.795 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 27.780 73.795 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 27.350 73.795 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 26.920 73.795 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 26.490 73.795 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 26.060 73.795 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 25.630 73.795 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 25.200 73.795 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 24.770 73.795 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 24.340 73.795 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 23.910 73.795 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 197.705 73.410 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 197.300 73.410 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 196.895 73.410 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 196.490 73.410 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 196.085 73.410 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 195.680 73.410 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 195.275 73.410 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 194.870 73.410 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 194.465 73.410 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 194.060 73.410 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 193.655 73.410 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 193.250 73.410 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 192.845 73.410 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 192.440 73.410 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 192.035 73.410 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 191.630 73.410 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 191.225 73.410 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 190.820 73.410 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 190.415 73.410 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 190.010 73.410 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 189.605 73.410 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 189.200 73.410 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 188.795 73.410 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 188.390 73.410 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 187.985 73.410 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 187.580 73.410 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 187.175 73.410 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 186.770 73.410 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 186.365 73.410 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 185.960 73.410 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 185.555 73.410 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 185.150 73.410 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 184.745 73.410 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 184.340 73.410 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 183.935 73.410 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 183.530 73.410 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 183.125 73.410 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 182.720 73.410 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 182.315 73.410 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 181.910 73.410 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 181.505 73.410 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 181.100 73.410 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 180.700 73.410 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 180.300 73.410 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 179.900 73.410 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 179.500 73.410 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 179.100 73.410 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 178.700 73.410 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 178.300 73.410 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 177.900 73.410 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 177.500 73.410 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 177.100 73.410 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 176.700 73.410 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 176.300 73.410 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 175.900 73.410 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 175.500 73.410 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 175.100 73.410 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 174.700 73.410 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 174.300 73.410 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.210 173.900 73.410 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 28.210 73.390 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 27.780 73.390 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 27.350 73.390 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 26.920 73.390 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 26.490 73.390 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 26.060 73.390 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 25.630 73.390 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 25.200 73.390 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 24.770 73.390 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 24.340 73.390 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 23.910 73.390 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 197.705 73.000 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 197.300 73.000 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 196.895 73.000 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 196.490 73.000 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 196.085 73.000 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 195.680 73.000 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 195.275 73.000 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 194.870 73.000 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 194.465 73.000 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 194.060 73.000 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 193.655 73.000 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 193.250 73.000 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 192.845 73.000 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 192.440 73.000 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 192.035 73.000 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 191.630 73.000 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 191.225 73.000 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 190.820 73.000 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 190.415 73.000 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 190.010 73.000 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 189.605 73.000 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 189.200 73.000 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 188.795 73.000 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 188.390 73.000 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 187.985 73.000 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 187.580 73.000 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 187.175 73.000 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 186.770 73.000 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 186.365 73.000 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 185.960 73.000 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 185.555 73.000 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 185.150 73.000 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 184.745 73.000 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 184.340 73.000 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 183.935 73.000 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 183.530 73.000 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 183.125 73.000 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 182.720 73.000 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 182.315 73.000 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 181.910 73.000 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 181.505 73.000 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 181.100 73.000 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 180.700 73.000 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 180.300 73.000 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 179.900 73.000 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 179.500 73.000 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 179.100 73.000 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 178.700 73.000 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 178.300 73.000 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 177.900 73.000 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 177.500 73.000 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 177.100 73.000 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 176.700 73.000 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 176.300 73.000 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 175.900 73.000 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 175.500 73.000 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 175.100 73.000 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 174.700 73.000 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 174.300 73.000 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.800 173.900 73.000 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 28.210 72.985 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 27.780 72.985 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 27.350 72.985 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 26.920 72.985 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 26.490 72.985 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 26.060 72.985 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 25.630 72.985 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 25.200 72.985 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 24.770 72.985 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 24.340 72.985 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 23.910 72.985 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 197.705 72.590 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 197.300 72.590 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 196.895 72.590 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 196.490 72.590 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 196.085 72.590 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 195.680 72.590 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 195.275 72.590 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 194.870 72.590 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 194.465 72.590 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 194.060 72.590 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 193.655 72.590 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 193.250 72.590 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 192.845 72.590 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 192.440 72.590 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 192.035 72.590 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 191.630 72.590 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 191.225 72.590 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 190.820 72.590 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 190.415 72.590 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 190.010 72.590 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 189.605 72.590 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 189.200 72.590 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 188.795 72.590 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 188.390 72.590 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 187.985 72.590 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 187.580 72.590 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 187.175 72.590 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 186.770 72.590 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 186.365 72.590 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 185.960 72.590 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 185.555 72.590 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 185.150 72.590 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 184.745 72.590 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 184.340 72.590 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 183.935 72.590 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 183.530 72.590 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 183.125 72.590 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 182.720 72.590 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 182.315 72.590 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 181.910 72.590 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 181.505 72.590 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 181.100 72.590 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 180.700 72.590 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 180.300 72.590 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 179.900 72.590 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 179.500 72.590 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 179.100 72.590 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 178.700 72.590 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 178.300 72.590 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 177.900 72.590 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 177.500 72.590 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 177.100 72.590 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 176.700 72.590 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 176.300 72.590 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 175.900 72.590 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 175.500 72.590 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 175.100 72.590 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 174.700 72.590 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 174.300 72.590 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.390 173.900 72.590 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 28.210 72.580 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 27.780 72.580 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 27.350 72.580 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 26.920 72.580 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 26.490 72.580 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 26.060 72.580 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 25.630 72.580 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 25.200 72.580 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 24.770 72.580 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 24.340 72.580 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 23.910 72.580 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 197.705 72.180 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 197.300 72.180 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 196.895 72.180 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 196.490 72.180 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 196.085 72.180 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 195.680 72.180 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 195.275 72.180 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 194.870 72.180 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 194.465 72.180 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 194.060 72.180 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 193.655 72.180 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 193.250 72.180 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 192.845 72.180 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 192.440 72.180 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 192.035 72.180 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 191.630 72.180 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 191.225 72.180 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 190.820 72.180 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 190.415 72.180 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 190.010 72.180 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 189.605 72.180 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 189.200 72.180 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 188.795 72.180 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 188.390 72.180 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 187.985 72.180 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 187.580 72.180 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 187.175 72.180 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 186.770 72.180 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 186.365 72.180 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 185.960 72.180 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 185.555 72.180 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 185.150 72.180 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 184.745 72.180 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 184.340 72.180 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 183.935 72.180 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 183.530 72.180 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 183.125 72.180 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 182.720 72.180 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 182.315 72.180 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 181.910 72.180 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 181.505 72.180 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 181.100 72.180 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 180.700 72.180 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 180.300 72.180 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 179.900 72.180 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 179.500 72.180 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 179.100 72.180 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 178.700 72.180 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 178.300 72.180 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 177.900 72.180 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 177.500 72.180 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 177.100 72.180 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 176.700 72.180 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 176.300 72.180 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 175.900 72.180 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 175.500 72.180 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 175.100 72.180 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 174.700 72.180 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 174.300 72.180 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.980 173.900 72.180 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 28.210 72.175 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 27.780 72.175 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 27.350 72.175 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 26.920 72.175 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 26.490 72.175 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 26.060 72.175 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 25.630 72.175 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 25.200 72.175 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 24.770 72.175 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 24.340 72.175 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 23.910 72.175 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 197.705 71.770 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 197.300 71.770 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 196.895 71.770 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 196.490 71.770 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 196.085 71.770 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 195.680 71.770 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 195.275 71.770 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 194.870 71.770 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 194.465 71.770 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 194.060 71.770 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 193.655 71.770 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 193.250 71.770 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 192.845 71.770 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 192.440 71.770 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 192.035 71.770 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 191.630 71.770 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 191.225 71.770 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 190.820 71.770 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 190.415 71.770 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 190.010 71.770 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 189.605 71.770 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 189.200 71.770 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 188.795 71.770 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 188.390 71.770 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 187.985 71.770 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 187.580 71.770 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 187.175 71.770 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 186.770 71.770 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 186.365 71.770 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 185.960 71.770 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 185.555 71.770 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 185.150 71.770 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 184.745 71.770 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 184.340 71.770 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 183.935 71.770 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 183.530 71.770 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 183.125 71.770 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 182.720 71.770 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 182.315 71.770 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 181.910 71.770 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 181.505 71.770 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 181.100 71.770 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 180.700 71.770 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 180.300 71.770 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 179.900 71.770 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 179.500 71.770 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 179.100 71.770 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 178.700 71.770 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 178.300 71.770 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 177.900 71.770 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 177.500 71.770 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 177.100 71.770 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 176.700 71.770 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 176.300 71.770 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 175.900 71.770 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 175.500 71.770 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 175.100 71.770 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 174.700 71.770 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 174.300 71.770 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 173.900 71.770 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 28.210 71.770 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 27.780 71.770 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 27.350 71.770 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 26.920 71.770 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 26.490 71.770 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 26.060 71.770 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 25.630 71.770 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 25.200 71.770 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 24.770 71.770 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 24.340 71.770 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 23.910 71.770 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 28.210 71.365 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 27.780 71.365 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 27.350 71.365 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 26.920 71.365 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 26.490 71.365 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 26.060 71.365 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 25.630 71.365 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 25.200 71.365 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 24.770 71.365 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 24.340 71.365 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 23.910 71.365 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 197.705 71.360 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 197.300 71.360 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 196.895 71.360 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 196.490 71.360 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 196.085 71.360 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 195.680 71.360 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 195.275 71.360 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 194.870 71.360 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 194.465 71.360 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 194.060 71.360 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 193.655 71.360 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 193.250 71.360 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 192.845 71.360 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 192.440 71.360 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 192.035 71.360 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 191.630 71.360 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 191.225 71.360 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 190.820 71.360 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 190.415 71.360 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 190.010 71.360 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 189.605 71.360 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 189.200 71.360 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 188.795 71.360 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 188.390 71.360 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 187.985 71.360 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 187.580 71.360 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 187.175 71.360 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 186.770 71.360 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 186.365 71.360 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 185.960 71.360 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 185.555 71.360 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 185.150 71.360 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 184.745 71.360 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 184.340 71.360 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 183.935 71.360 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 183.530 71.360 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 183.125 71.360 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 182.720 71.360 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 182.315 71.360 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 181.910 71.360 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 181.505 71.360 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 181.100 71.360 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 180.700 71.360 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 180.300 71.360 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 179.900 71.360 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 179.500 71.360 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 179.100 71.360 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 178.700 71.360 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 178.300 71.360 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 177.900 71.360 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 177.500 71.360 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 177.100 71.360 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 176.700 71.360 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 176.300 71.360 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 175.900 71.360 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 175.500 71.360 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 175.100 71.360 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 174.700 71.360 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 174.300 71.360 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.160 173.900 71.360 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 28.210 70.960 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 27.780 70.960 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 27.350 70.960 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 26.920 70.960 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 26.490 70.960 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 26.060 70.960 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 25.630 70.960 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 25.200 70.960 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 24.770 70.960 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 24.340 70.960 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 23.910 70.960 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 197.705 70.950 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 197.300 70.950 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 196.895 70.950 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 196.490 70.950 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 196.085 70.950 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 195.680 70.950 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 195.275 70.950 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 194.870 70.950 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 194.465 70.950 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 194.060 70.950 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 193.655 70.950 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 193.250 70.950 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 192.845 70.950 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 192.440 70.950 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 192.035 70.950 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 191.630 70.950 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 191.225 70.950 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 190.820 70.950 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 190.415 70.950 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 190.010 70.950 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 189.605 70.950 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 189.200 70.950 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 188.795 70.950 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 188.390 70.950 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 187.985 70.950 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 187.580 70.950 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 187.175 70.950 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 186.770 70.950 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 186.365 70.950 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 185.960 70.950 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 185.555 70.950 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 185.150 70.950 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 184.745 70.950 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 184.340 70.950 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 183.935 70.950 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 183.530 70.950 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 183.125 70.950 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 182.720 70.950 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 182.315 70.950 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 181.910 70.950 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 181.505 70.950 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 181.100 70.950 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 180.700 70.950 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 180.300 70.950 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 179.900 70.950 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 179.500 70.950 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 179.100 70.950 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 178.700 70.950 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 178.300 70.950 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 177.900 70.950 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 177.500 70.950 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 177.100 70.950 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 176.700 70.950 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 176.300 70.950 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 175.900 70.950 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 175.500 70.950 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 175.100 70.950 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 174.700 70.950 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 174.300 70.950 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.750 173.900 70.950 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 28.210 70.555 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 27.780 70.555 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 27.350 70.555 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 26.920 70.555 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 26.490 70.555 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 26.060 70.555 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 25.630 70.555 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 25.200 70.555 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 24.770 70.555 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 24.340 70.555 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 23.910 70.555 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 197.705 70.540 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 197.300 70.540 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 196.895 70.540 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 196.490 70.540 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 196.085 70.540 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 195.680 70.540 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 195.275 70.540 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 194.870 70.540 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 194.465 70.540 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 194.060 70.540 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 193.655 70.540 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 193.250 70.540 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 192.845 70.540 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 192.440 70.540 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 192.035 70.540 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 191.630 70.540 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 191.225 70.540 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 190.820 70.540 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 190.415 70.540 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 190.010 70.540 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 189.605 70.540 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 189.200 70.540 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 188.795 70.540 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 188.390 70.540 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 187.985 70.540 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 187.580 70.540 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 187.175 70.540 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 186.770 70.540 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 186.365 70.540 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 185.960 70.540 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 185.555 70.540 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 185.150 70.540 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 184.745 70.540 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 184.340 70.540 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 183.935 70.540 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 183.530 70.540 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 183.125 70.540 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 182.720 70.540 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 182.315 70.540 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 181.910 70.540 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 181.505 70.540 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 181.100 70.540 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 180.700 70.540 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 180.300 70.540 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 179.900 70.540 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 179.500 70.540 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 179.100 70.540 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 178.700 70.540 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 178.300 70.540 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 177.900 70.540 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 177.500 70.540 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 177.100 70.540 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 176.700 70.540 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 176.300 70.540 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 175.900 70.540 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 175.500 70.540 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 175.100 70.540 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 174.700 70.540 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 174.300 70.540 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.340 173.900 70.540 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 28.210 70.150 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 27.780 70.150 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 27.350 70.150 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 26.920 70.150 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 26.490 70.150 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 26.060 70.150 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 25.630 70.150 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 25.200 70.150 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 24.770 70.150 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 24.340 70.150 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 23.910 70.150 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 197.705 70.130 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 197.300 70.130 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 196.895 70.130 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 196.490 70.130 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 196.085 70.130 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 195.680 70.130 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 195.275 70.130 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 194.870 70.130 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 194.465 70.130 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 194.060 70.130 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 193.655 70.130 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 193.250 70.130 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 192.845 70.130 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 192.440 70.130 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 192.035 70.130 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 191.630 70.130 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 191.225 70.130 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 190.820 70.130 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 190.415 70.130 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 190.010 70.130 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 189.605 70.130 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 189.200 70.130 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 188.795 70.130 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 188.390 70.130 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 187.985 70.130 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 187.580 70.130 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 187.175 70.130 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 186.770 70.130 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 186.365 70.130 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 185.960 70.130 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 185.555 70.130 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 185.150 70.130 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 184.745 70.130 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 184.340 70.130 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 183.935 70.130 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 183.530 70.130 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 183.125 70.130 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 182.720 70.130 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 182.315 70.130 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 181.910 70.130 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 181.505 70.130 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 181.100 70.130 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 180.700 70.130 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 180.300 70.130 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 179.900 70.130 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 179.500 70.130 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 179.100 70.130 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 178.700 70.130 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 178.300 70.130 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 177.900 70.130 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 177.500 70.130 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 177.100 70.130 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 176.700 70.130 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 176.300 70.130 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 175.900 70.130 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 175.500 70.130 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 175.100 70.130 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 174.700 70.130 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 174.300 70.130 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.930 173.900 70.130 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 28.210 69.745 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 27.780 69.745 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 27.350 69.745 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 26.920 69.745 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 26.490 69.745 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 26.060 69.745 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 25.630 69.745 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 25.200 69.745 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 24.770 69.745 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 24.340 69.745 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 23.910 69.745 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 197.705 69.720 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 197.300 69.720 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 196.895 69.720 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 196.490 69.720 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 196.085 69.720 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 195.680 69.720 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 195.275 69.720 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 194.870 69.720 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 194.465 69.720 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 194.060 69.720 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 193.655 69.720 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 193.250 69.720 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 192.845 69.720 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 192.440 69.720 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 192.035 69.720 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 191.630 69.720 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 191.225 69.720 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 190.820 69.720 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 190.415 69.720 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 190.010 69.720 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 189.605 69.720 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 189.200 69.720 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 188.795 69.720 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 188.390 69.720 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 187.985 69.720 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 187.580 69.720 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 187.175 69.720 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 186.770 69.720 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 186.365 69.720 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 185.960 69.720 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 185.555 69.720 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 185.150 69.720 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 184.745 69.720 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 184.340 69.720 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 183.935 69.720 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 183.530 69.720 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 183.125 69.720 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 182.720 69.720 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 182.315 69.720 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 181.910 69.720 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 181.505 69.720 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 181.100 69.720 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 180.700 69.720 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 180.300 69.720 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 179.900 69.720 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 179.500 69.720 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 179.100 69.720 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 178.700 69.720 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 178.300 69.720 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 177.900 69.720 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 177.500 69.720 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 177.100 69.720 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 176.700 69.720 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 176.300 69.720 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 175.900 69.720 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 175.500 69.720 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 175.100 69.720 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 174.700 69.720 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 174.300 69.720 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.520 173.900 69.720 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 28.210 69.340 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 27.780 69.340 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 27.350 69.340 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 26.920 69.340 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 26.490 69.340 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 26.060 69.340 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 25.630 69.340 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 25.200 69.340 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 24.770 69.340 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 24.340 69.340 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 23.910 69.340 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 197.705 69.310 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 197.300 69.310 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 196.895 69.310 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 196.490 69.310 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 196.085 69.310 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 195.680 69.310 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 195.275 69.310 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 194.870 69.310 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 194.465 69.310 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 194.060 69.310 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 193.655 69.310 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 193.250 69.310 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 192.845 69.310 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 192.440 69.310 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 192.035 69.310 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 191.630 69.310 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 191.225 69.310 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 190.820 69.310 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 190.415 69.310 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 190.010 69.310 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 189.605 69.310 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 189.200 69.310 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 188.795 69.310 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 188.390 69.310 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 187.985 69.310 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 187.580 69.310 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 187.175 69.310 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 186.770 69.310 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 186.365 69.310 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 185.960 69.310 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 185.555 69.310 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 185.150 69.310 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 184.745 69.310 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 184.340 69.310 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 183.935 69.310 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 183.530 69.310 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 183.125 69.310 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 182.720 69.310 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 182.315 69.310 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 181.910 69.310 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 181.505 69.310 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 181.100 69.310 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 180.700 69.310 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 180.300 69.310 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 179.900 69.310 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 179.500 69.310 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 179.100 69.310 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 178.700 69.310 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 178.300 69.310 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 177.900 69.310 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 177.500 69.310 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 177.100 69.310 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 176.700 69.310 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 176.300 69.310 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 175.900 69.310 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 175.500 69.310 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 175.100 69.310 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 174.700 69.310 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 174.300 69.310 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.110 173.900 69.310 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 28.210 68.935 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 27.780 68.935 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 27.350 68.935 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 26.920 68.935 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 26.490 68.935 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 26.060 68.935 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 25.630 68.935 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 25.200 68.935 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 24.770 68.935 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 24.340 68.935 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 23.910 68.935 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 197.705 68.900 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 197.300 68.900 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 196.895 68.900 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 196.490 68.900 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 196.085 68.900 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 195.680 68.900 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 195.275 68.900 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 194.870 68.900 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 194.465 68.900 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 194.060 68.900 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 193.655 68.900 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 193.250 68.900 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 192.845 68.900 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 192.440 68.900 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 192.035 68.900 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 191.630 68.900 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 191.225 68.900 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 190.820 68.900 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 190.415 68.900 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 190.010 68.900 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 189.605 68.900 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 189.200 68.900 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 188.795 68.900 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 188.390 68.900 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 187.985 68.900 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 187.580 68.900 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 187.175 68.900 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 186.770 68.900 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 186.365 68.900 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 185.960 68.900 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 185.555 68.900 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 185.150 68.900 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 184.745 68.900 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 184.340 68.900 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 183.935 68.900 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 183.530 68.900 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 183.125 68.900 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 182.720 68.900 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 182.315 68.900 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 181.910 68.900 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 181.505 68.900 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 181.100 68.900 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 180.700 68.900 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 180.300 68.900 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 179.900 68.900 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 179.500 68.900 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 179.100 68.900 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 178.700 68.900 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 178.300 68.900 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 177.900 68.900 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 177.500 68.900 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 177.100 68.900 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 176.700 68.900 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 176.300 68.900 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 175.900 68.900 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 175.500 68.900 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 175.100 68.900 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 174.700 68.900 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 174.300 68.900 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.700 173.900 68.900 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 28.210 68.530 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 27.780 68.530 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 27.350 68.530 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 26.920 68.530 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 26.490 68.530 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 26.060 68.530 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 25.630 68.530 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 25.200 68.530 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 24.770 68.530 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 24.340 68.530 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 23.910 68.530 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 197.705 68.490 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 197.300 68.490 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 196.895 68.490 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 196.490 68.490 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 196.085 68.490 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 195.680 68.490 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 195.275 68.490 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 194.870 68.490 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 194.465 68.490 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 194.060 68.490 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 193.655 68.490 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 193.250 68.490 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 192.845 68.490 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 192.440 68.490 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 192.035 68.490 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 191.630 68.490 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 191.225 68.490 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 190.820 68.490 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 190.415 68.490 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 190.010 68.490 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 189.605 68.490 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 189.200 68.490 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 188.795 68.490 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 188.390 68.490 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 187.985 68.490 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 187.580 68.490 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 187.175 68.490 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 186.770 68.490 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 186.365 68.490 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 185.960 68.490 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 185.555 68.490 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 185.150 68.490 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 184.745 68.490 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 184.340 68.490 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 183.935 68.490 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 183.530 68.490 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 183.125 68.490 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 182.720 68.490 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 182.315 68.490 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 181.910 68.490 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 181.505 68.490 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 181.100 68.490 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 180.700 68.490 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 180.300 68.490 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 179.900 68.490 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 179.500 68.490 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 179.100 68.490 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 178.700 68.490 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 178.300 68.490 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 177.900 68.490 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 177.500 68.490 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 177.100 68.490 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 176.700 68.490 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 176.300 68.490 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 175.900 68.490 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 175.500 68.490 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 175.100 68.490 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 174.700 68.490 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 174.300 68.490 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.290 173.900 68.490 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 28.210 68.125 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 27.780 68.125 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 27.350 68.125 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 26.920 68.125 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 26.490 68.125 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 26.060 68.125 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 25.630 68.125 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 25.200 68.125 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 24.770 68.125 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 24.340 68.125 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 23.910 68.125 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 197.705 68.080 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 197.300 68.080 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 196.895 68.080 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 196.490 68.080 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 196.085 68.080 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 195.680 68.080 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 195.275 68.080 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 194.870 68.080 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 194.465 68.080 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 194.060 68.080 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 193.655 68.080 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 193.250 68.080 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 192.845 68.080 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 192.440 68.080 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 192.035 68.080 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 191.630 68.080 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 191.225 68.080 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 190.820 68.080 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 190.415 68.080 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 190.010 68.080 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 189.605 68.080 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 189.200 68.080 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 188.795 68.080 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 188.390 68.080 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 187.985 68.080 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 187.580 68.080 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 187.175 68.080 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 186.770 68.080 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 186.365 68.080 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 185.960 68.080 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 185.555 68.080 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 185.150 68.080 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 184.745 68.080 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 184.340 68.080 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 183.935 68.080 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 183.530 68.080 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 183.125 68.080 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 182.720 68.080 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 182.315 68.080 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 181.910 68.080 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 181.505 68.080 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 181.100 68.080 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 180.700 68.080 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 180.300 68.080 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 179.900 68.080 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 179.500 68.080 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 179.100 68.080 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 178.700 68.080 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 178.300 68.080 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 177.900 68.080 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 177.500 68.080 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 177.100 68.080 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 176.700 68.080 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 176.300 68.080 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 175.900 68.080 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 175.500 68.080 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 175.100 68.080 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 174.700 68.080 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 174.300 68.080 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.880 173.900 68.080 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 28.210 67.720 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 27.780 67.720 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 27.350 67.720 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 26.920 67.720 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 26.490 67.720 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 26.060 67.720 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 25.630 67.720 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 25.200 67.720 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 24.770 67.720 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 24.340 67.720 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 23.910 67.720 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 197.705 67.670 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 197.300 67.670 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 196.895 67.670 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 196.490 67.670 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 196.085 67.670 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 195.680 67.670 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 195.275 67.670 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 194.870 67.670 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 194.465 67.670 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 194.060 67.670 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 193.655 67.670 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 193.250 67.670 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 192.845 67.670 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 192.440 67.670 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 192.035 67.670 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 191.630 67.670 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 191.225 67.670 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 190.820 67.670 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 190.415 67.670 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 190.010 67.670 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 189.605 67.670 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 189.200 67.670 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 188.795 67.670 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 188.390 67.670 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 187.985 67.670 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 187.580 67.670 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 187.175 67.670 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 186.770 67.670 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 186.365 67.670 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 185.960 67.670 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 185.555 67.670 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 185.150 67.670 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 184.745 67.670 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 184.340 67.670 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 183.935 67.670 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 183.530 67.670 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 183.125 67.670 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 182.720 67.670 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 182.315 67.670 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 181.910 67.670 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 181.505 67.670 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 181.100 67.670 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 180.700 67.670 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 180.300 67.670 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 179.900 67.670 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 179.500 67.670 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 179.100 67.670 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 178.700 67.670 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 178.300 67.670 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 177.900 67.670 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 177.500 67.670 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 177.100 67.670 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 176.700 67.670 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 176.300 67.670 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 175.900 67.670 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 175.500 67.670 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 175.100 67.670 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 174.700 67.670 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 174.300 67.670 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.470 173.900 67.670 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 28.210 67.315 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 27.780 67.315 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 27.350 67.315 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 26.920 67.315 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 26.490 67.315 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 26.060 67.315 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 25.630 67.315 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 25.200 67.315 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 24.770 67.315 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 24.340 67.315 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 23.910 67.315 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 197.705 67.260 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 197.300 67.260 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 196.895 67.260 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 196.490 67.260 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 196.085 67.260 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 195.680 67.260 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 195.275 67.260 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 194.870 67.260 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 194.465 67.260 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 194.060 67.260 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 193.655 67.260 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 193.250 67.260 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 192.845 67.260 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 192.440 67.260 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 192.035 67.260 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 191.630 67.260 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 191.225 67.260 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 190.820 67.260 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 190.415 67.260 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 190.010 67.260 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 189.605 67.260 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 189.200 67.260 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 188.795 67.260 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 188.390 67.260 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 187.985 67.260 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 187.580 67.260 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 187.175 67.260 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 186.770 67.260 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 186.365 67.260 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 185.960 67.260 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 185.555 67.260 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 185.150 67.260 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 184.745 67.260 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 184.340 67.260 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 183.935 67.260 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 183.530 67.260 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 183.125 67.260 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 182.720 67.260 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 182.315 67.260 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 181.910 67.260 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 181.505 67.260 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 181.100 67.260 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 180.700 67.260 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 180.300 67.260 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 179.900 67.260 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 179.500 67.260 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 179.100 67.260 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 178.700 67.260 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 178.300 67.260 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 177.900 67.260 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 177.500 67.260 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 177.100 67.260 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 176.700 67.260 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 176.300 67.260 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 175.900 67.260 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 175.500 67.260 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 175.100 67.260 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 174.700 67.260 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 174.300 67.260 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.060 173.900 67.260 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 28.210 66.910 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 27.780 66.910 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 27.350 66.910 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 26.920 66.910 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 26.490 66.910 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 26.060 66.910 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 25.630 66.910 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 25.200 66.910 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 24.770 66.910 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 24.340 66.910 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 23.910 66.910 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 197.705 66.850 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 197.300 66.850 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 196.895 66.850 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 196.490 66.850 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 196.085 66.850 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 195.680 66.850 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 195.275 66.850 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 194.870 66.850 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 194.465 66.850 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 194.060 66.850 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 193.655 66.850 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 193.250 66.850 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 192.845 66.850 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 192.440 66.850 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 192.035 66.850 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 191.630 66.850 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 191.225 66.850 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 190.820 66.850 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 190.415 66.850 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 190.010 66.850 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 189.605 66.850 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 189.200 66.850 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 188.795 66.850 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 188.390 66.850 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 187.985 66.850 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 187.580 66.850 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 187.175 66.850 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 186.770 66.850 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 186.365 66.850 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 185.960 66.850 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 185.555 66.850 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 185.150 66.850 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 184.745 66.850 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 184.340 66.850 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 183.935 66.850 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 183.530 66.850 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 183.125 66.850 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 182.720 66.850 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 182.315 66.850 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 181.910 66.850 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 181.505 66.850 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 181.100 66.850 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 180.700 66.850 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 180.300 66.850 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 179.900 66.850 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 179.500 66.850 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 179.100 66.850 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 178.700 66.850 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 178.300 66.850 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 177.900 66.850 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 177.500 66.850 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 177.100 66.850 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 176.700 66.850 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 176.300 66.850 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 175.900 66.850 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 175.500 66.850 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 175.100 66.850 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 174.700 66.850 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 174.300 66.850 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.650 173.900 66.850 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 28.210 66.505 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 27.780 66.505 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 27.350 66.505 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 26.920 66.505 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 26.490 66.505 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 26.060 66.505 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 25.630 66.505 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 25.200 66.505 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 24.770 66.505 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 24.340 66.505 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 23.910 66.505 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 197.705 66.440 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 197.300 66.440 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 196.895 66.440 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 196.490 66.440 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 196.085 66.440 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 195.680 66.440 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 195.275 66.440 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 194.870 66.440 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 194.465 66.440 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 194.060 66.440 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 193.655 66.440 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 193.250 66.440 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 192.845 66.440 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 192.440 66.440 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 192.035 66.440 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 191.630 66.440 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 191.225 66.440 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 190.820 66.440 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 190.415 66.440 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 190.010 66.440 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 189.605 66.440 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 189.200 66.440 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 188.795 66.440 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 188.390 66.440 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 187.985 66.440 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 187.580 66.440 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 187.175 66.440 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 186.770 66.440 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 186.365 66.440 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 185.960 66.440 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 185.555 66.440 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 185.150 66.440 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 184.745 66.440 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 184.340 66.440 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 183.935 66.440 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 183.530 66.440 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 183.125 66.440 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 182.720 66.440 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 182.315 66.440 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 181.910 66.440 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 181.505 66.440 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 181.100 66.440 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 180.700 66.440 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 180.300 66.440 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 179.900 66.440 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 179.500 66.440 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 179.100 66.440 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 178.700 66.440 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 178.300 66.440 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 177.900 66.440 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 177.500 66.440 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 177.100 66.440 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 176.700 66.440 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 176.300 66.440 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 175.900 66.440 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 175.500 66.440 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 175.100 66.440 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 174.700 66.440 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 174.300 66.440 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.240 173.900 66.440 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 28.210 66.100 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 27.780 66.100 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 27.350 66.100 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 26.920 66.100 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 26.490 66.100 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 26.060 66.100 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 25.630 66.100 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 25.200 66.100 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 24.770 66.100 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 24.340 66.100 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 23.910 66.100 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 197.705 66.030 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 197.300 66.030 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 196.895 66.030 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 196.490 66.030 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 196.085 66.030 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 195.680 66.030 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 195.275 66.030 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 194.870 66.030 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 194.465 66.030 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 194.060 66.030 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 193.655 66.030 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 193.250 66.030 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 192.845 66.030 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 192.440 66.030 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 192.035 66.030 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 191.630 66.030 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 191.225 66.030 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 190.820 66.030 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 190.415 66.030 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 190.010 66.030 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 189.605 66.030 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 189.200 66.030 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 188.795 66.030 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 188.390 66.030 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 187.985 66.030 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 187.580 66.030 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 187.175 66.030 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 186.770 66.030 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 186.365 66.030 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 185.960 66.030 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 185.555 66.030 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 185.150 66.030 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 184.745 66.030 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 184.340 66.030 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 183.935 66.030 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 183.530 66.030 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 183.125 66.030 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 182.720 66.030 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 182.315 66.030 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 181.910 66.030 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 181.505 66.030 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 181.100 66.030 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 180.700 66.030 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 180.300 66.030 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 179.900 66.030 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 179.500 66.030 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 179.100 66.030 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 178.700 66.030 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 178.300 66.030 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 177.900 66.030 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 177.500 66.030 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 177.100 66.030 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 176.700 66.030 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 176.300 66.030 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 175.900 66.030 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 175.500 66.030 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 175.100 66.030 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 174.700 66.030 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 174.300 66.030 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.830 173.900 66.030 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 28.210 65.695 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 27.780 65.695 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 27.350 65.695 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 26.920 65.695 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 26.490 65.695 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 26.060 65.695 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 25.630 65.695 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 25.200 65.695 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 24.770 65.695 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 24.340 65.695 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 23.910 65.695 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 197.705 65.620 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 197.300 65.620 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 196.895 65.620 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 196.490 65.620 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 196.085 65.620 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 195.680 65.620 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 195.275 65.620 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 194.870 65.620 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 194.465 65.620 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 194.060 65.620 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 193.655 65.620 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 193.250 65.620 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 192.845 65.620 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 192.440 65.620 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 192.035 65.620 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 191.630 65.620 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 191.225 65.620 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 190.820 65.620 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 190.415 65.620 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 190.010 65.620 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 189.605 65.620 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 189.200 65.620 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 188.795 65.620 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 188.390 65.620 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 187.985 65.620 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 187.580 65.620 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 187.175 65.620 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 186.770 65.620 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 186.365 65.620 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 185.960 65.620 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 185.555 65.620 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 185.150 65.620 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 184.745 65.620 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 184.340 65.620 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 183.935 65.620 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 183.530 65.620 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 183.125 65.620 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 182.720 65.620 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 182.315 65.620 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 181.910 65.620 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 181.505 65.620 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 181.100 65.620 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 180.700 65.620 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 180.300 65.620 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 179.900 65.620 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 179.500 65.620 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 179.100 65.620 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 178.700 65.620 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 178.300 65.620 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 177.900 65.620 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 177.500 65.620 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 177.100 65.620 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 176.700 65.620 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 176.300 65.620 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 175.900 65.620 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 175.500 65.620 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 175.100 65.620 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 174.700 65.620 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 174.300 65.620 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.420 173.900 65.620 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 28.210 65.290 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 27.780 65.290 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 27.350 65.290 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 26.920 65.290 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 26.490 65.290 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 26.060 65.290 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 25.630 65.290 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 25.200 65.290 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 24.770 65.290 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 24.340 65.290 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 23.910 65.290 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 197.705 65.210 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 197.300 65.210 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 196.895 65.210 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 196.490 65.210 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 196.085 65.210 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 195.680 65.210 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 195.275 65.210 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 194.870 65.210 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 194.465 65.210 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 194.060 65.210 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 193.655 65.210 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 193.250 65.210 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 192.845 65.210 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 192.440 65.210 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 192.035 65.210 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 191.630 65.210 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 191.225 65.210 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 190.820 65.210 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 190.415 65.210 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 190.010 65.210 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 189.605 65.210 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 189.200 65.210 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 188.795 65.210 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 188.390 65.210 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 187.985 65.210 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 187.580 65.210 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 187.175 65.210 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 186.770 65.210 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 186.365 65.210 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 185.960 65.210 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 185.555 65.210 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 185.150 65.210 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 184.745 65.210 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 184.340 65.210 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 183.935 65.210 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 183.530 65.210 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 183.125 65.210 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 182.720 65.210 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 182.315 65.210 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 181.910 65.210 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 181.505 65.210 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 181.100 65.210 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 180.700 65.210 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 180.300 65.210 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 179.900 65.210 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 179.500 65.210 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 179.100 65.210 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 178.700 65.210 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 178.300 65.210 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 177.900 65.210 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 177.500 65.210 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 177.100 65.210 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 176.700 65.210 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 176.300 65.210 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 175.900 65.210 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 175.500 65.210 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 175.100 65.210 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 174.700 65.210 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 174.300 65.210 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.010 173.900 65.210 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 28.210 64.885 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 27.780 64.885 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 27.350 64.885 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 26.920 64.885 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 26.490 64.885 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 26.060 64.885 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 25.630 64.885 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 25.200 64.885 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 24.770 64.885 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 24.340 64.885 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 23.910 64.885 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 197.705 64.800 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 197.300 64.800 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 196.895 64.800 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 196.490 64.800 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 196.085 64.800 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 195.680 64.800 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 195.275 64.800 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 194.870 64.800 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 194.465 64.800 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 194.060 64.800 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 193.655 64.800 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 193.250 64.800 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 192.845 64.800 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 192.440 64.800 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 192.035 64.800 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 191.630 64.800 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 191.225 64.800 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 190.820 64.800 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 190.415 64.800 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 190.010 64.800 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 189.605 64.800 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 189.200 64.800 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 188.795 64.800 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 188.390 64.800 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 187.985 64.800 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 187.580 64.800 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 187.175 64.800 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 186.770 64.800 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 186.365 64.800 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 185.960 64.800 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 185.555 64.800 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 185.150 64.800 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 184.745 64.800 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 184.340 64.800 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 183.935 64.800 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 183.530 64.800 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 183.125 64.800 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 182.720 64.800 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 182.315 64.800 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 181.910 64.800 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 181.505 64.800 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 181.100 64.800 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 180.700 64.800 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 180.300 64.800 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 179.900 64.800 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 179.500 64.800 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 179.100 64.800 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 178.700 64.800 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 178.300 64.800 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 177.900 64.800 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 177.500 64.800 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 177.100 64.800 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 176.700 64.800 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 176.300 64.800 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 175.900 64.800 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 175.500 64.800 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 175.100 64.800 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 174.700 64.800 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 174.300 64.800 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.600 173.900 64.800 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 28.210 64.480 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 27.780 64.480 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 27.350 64.480 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 26.920 64.480 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 26.490 64.480 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 26.060 64.480 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 25.630 64.480 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 25.200 64.480 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 24.770 64.480 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 24.340 64.480 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 23.910 64.480 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 197.705 64.390 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 197.300 64.390 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 196.895 64.390 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 196.490 64.390 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 196.085 64.390 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 195.680 64.390 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 195.275 64.390 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 194.870 64.390 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 194.465 64.390 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 194.060 64.390 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 193.655 64.390 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 193.250 64.390 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 192.845 64.390 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 192.440 64.390 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 192.035 64.390 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 191.630 64.390 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 191.225 64.390 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 190.820 64.390 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 190.415 64.390 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 190.010 64.390 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 189.605 64.390 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 189.200 64.390 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 188.795 64.390 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 188.390 64.390 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 187.985 64.390 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 187.580 64.390 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 187.175 64.390 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 186.770 64.390 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 186.365 64.390 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 185.960 64.390 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 185.555 64.390 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 185.150 64.390 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 184.745 64.390 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 184.340 64.390 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 183.935 64.390 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 183.530 64.390 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 183.125 64.390 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 182.720 64.390 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 182.315 64.390 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 181.910 64.390 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 181.505 64.390 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 181.100 64.390 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 180.700 64.390 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 180.300 64.390 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 179.900 64.390 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 179.500 64.390 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 179.100 64.390 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 178.700 64.390 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 178.300 64.390 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 177.900 64.390 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 177.500 64.390 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 177.100 64.390 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 176.700 64.390 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 176.300 64.390 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 175.900 64.390 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 175.500 64.390 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 175.100 64.390 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 174.700 64.390 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 174.300 64.390 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.190 173.900 64.390 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 28.210 64.075 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 27.780 64.075 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 27.350 64.075 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 26.920 64.075 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 26.490 64.075 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 26.060 64.075 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 25.630 64.075 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 25.200 64.075 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 24.770 64.075 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 24.340 64.075 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 23.910 64.075 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 197.705 63.980 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 197.300 63.980 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 196.895 63.980 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 196.490 63.980 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 196.085 63.980 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 195.680 63.980 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 195.275 63.980 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 194.870 63.980 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 194.465 63.980 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 194.060 63.980 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 193.655 63.980 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 193.250 63.980 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 192.845 63.980 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 192.440 63.980 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 192.035 63.980 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 191.630 63.980 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 191.225 63.980 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 190.820 63.980 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 190.415 63.980 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 190.010 63.980 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 189.605 63.980 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 189.200 63.980 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 188.795 63.980 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 188.390 63.980 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 187.985 63.980 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 187.580 63.980 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 187.175 63.980 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 186.770 63.980 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 186.365 63.980 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 185.960 63.980 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 185.555 63.980 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 185.150 63.980 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 184.745 63.980 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 184.340 63.980 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 183.935 63.980 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 183.530 63.980 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 183.125 63.980 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 182.720 63.980 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 182.315 63.980 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 181.910 63.980 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 181.505 63.980 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 181.100 63.980 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 180.700 63.980 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 180.300 63.980 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 179.900 63.980 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 179.500 63.980 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 179.100 63.980 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 178.700 63.980 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 178.300 63.980 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 177.900 63.980 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 177.500 63.980 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 177.100 63.980 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 176.700 63.980 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 176.300 63.980 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 175.900 63.980 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 175.500 63.980 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 175.100 63.980 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 174.700 63.980 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 174.300 63.980 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.780 173.900 63.980 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 28.210 63.670 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 27.780 63.670 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 27.350 63.670 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 26.920 63.670 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 26.490 63.670 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 26.060 63.670 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 25.630 63.670 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 25.200 63.670 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 24.770 63.670 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 24.340 63.670 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 23.910 63.670 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 197.705 63.570 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 197.300 63.570 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 196.895 63.570 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 196.490 63.570 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 196.085 63.570 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 195.680 63.570 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 195.275 63.570 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 194.870 63.570 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 194.465 63.570 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 194.060 63.570 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 193.655 63.570 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 193.250 63.570 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 192.845 63.570 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 192.440 63.570 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 192.035 63.570 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 191.630 63.570 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 191.225 63.570 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 190.820 63.570 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 190.415 63.570 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 190.010 63.570 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 189.605 63.570 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 189.200 63.570 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 188.795 63.570 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 188.390 63.570 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 187.985 63.570 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 187.580 63.570 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 187.175 63.570 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 186.770 63.570 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 186.365 63.570 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 185.960 63.570 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 185.555 63.570 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 185.150 63.570 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 184.745 63.570 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 184.340 63.570 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 183.935 63.570 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 183.530 63.570 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 183.125 63.570 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 182.720 63.570 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 182.315 63.570 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 181.910 63.570 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 181.505 63.570 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 181.100 63.570 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 180.700 63.570 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 180.300 63.570 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 179.900 63.570 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 179.500 63.570 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 179.100 63.570 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 178.700 63.570 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 178.300 63.570 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 177.900 63.570 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 177.500 63.570 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 177.100 63.570 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 176.700 63.570 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 176.300 63.570 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 175.900 63.570 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 175.500 63.570 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 175.100 63.570 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 174.700 63.570 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 174.300 63.570 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.370 173.900 63.570 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 28.210 63.265 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 27.780 63.265 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 27.350 63.265 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 26.920 63.265 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 26.490 63.265 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 26.060 63.265 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 25.630 63.265 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 25.200 63.265 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 24.770 63.265 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 24.340 63.265 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 23.910 63.265 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 197.705 63.160 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 197.300 63.160 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 196.895 63.160 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 196.490 63.160 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 196.085 63.160 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 195.680 63.160 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 195.275 63.160 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 194.870 63.160 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 194.465 63.160 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 194.060 63.160 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 193.655 63.160 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 193.250 63.160 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 192.845 63.160 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 192.440 63.160 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 192.035 63.160 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 191.630 63.160 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 191.225 63.160 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 190.820 63.160 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 190.415 63.160 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 190.010 63.160 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 189.605 63.160 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 189.200 63.160 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 188.795 63.160 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 188.390 63.160 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 187.985 63.160 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 187.580 63.160 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 187.175 63.160 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 186.770 63.160 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 186.365 63.160 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 185.960 63.160 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 185.555 63.160 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 185.150 63.160 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 184.745 63.160 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 184.340 63.160 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 183.935 63.160 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 183.530 63.160 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 183.125 63.160 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 182.720 63.160 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 182.315 63.160 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 181.910 63.160 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 181.505 63.160 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 181.100 63.160 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 180.700 63.160 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 180.300 63.160 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 179.900 63.160 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 179.500 63.160 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 179.100 63.160 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 178.700 63.160 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 178.300 63.160 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 177.900 63.160 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 177.500 63.160 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 177.100 63.160 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 176.700 63.160 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 176.300 63.160 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 175.900 63.160 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 175.500 63.160 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 175.100 63.160 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 174.700 63.160 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 174.300 63.160 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.960 173.900 63.160 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 28.210 62.860 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 27.780 62.860 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 27.350 62.860 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 26.920 62.860 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 26.490 62.860 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 26.060 62.860 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 25.630 62.860 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 25.200 62.860 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 24.770 62.860 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 24.340 62.860 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 23.910 62.860 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 197.705 62.750 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 197.300 62.750 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 196.895 62.750 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 196.490 62.750 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 196.085 62.750 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 195.680 62.750 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 195.275 62.750 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 194.870 62.750 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 194.465 62.750 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 194.060 62.750 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 193.655 62.750 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 193.250 62.750 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 192.845 62.750 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 192.440 62.750 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 192.035 62.750 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 191.630 62.750 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 191.225 62.750 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 190.820 62.750 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 190.415 62.750 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 190.010 62.750 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 189.605 62.750 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 189.200 62.750 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 188.795 62.750 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 188.390 62.750 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 187.985 62.750 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 187.580 62.750 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 187.175 62.750 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 186.770 62.750 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 186.365 62.750 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 185.960 62.750 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 185.555 62.750 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 185.150 62.750 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 184.745 62.750 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 184.340 62.750 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 183.935 62.750 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 183.530 62.750 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 183.125 62.750 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 182.720 62.750 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 182.315 62.750 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 181.910 62.750 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 181.505 62.750 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 181.100 62.750 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 180.700 62.750 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 180.300 62.750 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 179.900 62.750 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 179.500 62.750 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 179.100 62.750 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 178.700 62.750 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 178.300 62.750 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 177.900 62.750 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 177.500 62.750 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 177.100 62.750 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 176.700 62.750 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 176.300 62.750 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 175.900 62.750 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 175.500 62.750 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 175.100 62.750 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 174.700 62.750 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 174.300 62.750 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.550 173.900 62.750 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 28.210 62.455 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 27.780 62.455 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 27.350 62.455 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 26.920 62.455 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 26.490 62.455 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 26.060 62.455 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 25.630 62.455 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 25.200 62.455 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 24.770 62.455 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 24.340 62.455 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 23.910 62.455 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 197.705 62.340 197.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 197.300 62.340 197.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 196.895 62.340 197.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 196.490 62.340 196.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 196.085 62.340 196.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 195.680 62.340 195.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 195.275 62.340 195.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 194.870 62.340 195.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 194.465 62.340 194.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 194.060 62.340 194.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 193.655 62.340 193.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 193.250 62.340 193.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 192.845 62.340 193.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 192.440 62.340 192.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 192.035 62.340 192.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 191.630 62.340 191.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 191.225 62.340 191.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 190.820 62.340 191.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 190.415 62.340 190.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 190.010 62.340 190.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 189.605 62.340 189.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 189.200 62.340 189.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 188.795 62.340 188.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 188.390 62.340 188.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 187.985 62.340 188.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 187.580 62.340 187.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 187.175 62.340 187.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 186.770 62.340 186.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 186.365 62.340 186.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 185.960 62.340 186.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 185.555 62.340 185.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 185.150 62.340 185.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 184.745 62.340 184.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 184.340 62.340 184.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 183.935 62.340 184.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 183.530 62.340 183.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 183.125 62.340 183.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 182.720 62.340 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 182.315 62.340 182.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 181.910 62.340 182.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 181.505 62.340 181.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 181.100 62.340 181.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 180.700 62.340 180.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 180.300 62.340 180.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 179.900 62.340 180.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 179.500 62.340 179.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 179.100 62.340 179.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 178.700 62.340 178.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 178.300 62.340 178.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 177.900 62.340 178.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 177.500 62.340 177.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 177.100 62.340 177.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 176.700 62.340 176.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 176.300 62.340 176.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 175.900 62.340 176.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 175.500 62.340 175.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 175.100 62.340 175.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 174.700 62.340 174.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 174.300 62.340 174.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.140 173.900 62.340 174.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 28.210 62.050 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 27.780 62.050 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 27.350 62.050 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 26.920 62.050 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 26.490 62.050 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 26.060 62.050 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 25.630 62.050 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 25.200 62.050 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 24.770 62.050 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 24.340 62.050 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 23.910 62.050 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 28.210 61.645 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 27.780 61.645 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 27.350 61.645 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 26.920 61.645 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 26.490 61.645 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 26.060 61.645 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 25.630 61.645 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 25.200 61.645 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 24.770 61.645 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 24.340 61.645 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 23.910 61.645 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 28.210 61.240 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 27.780 61.240 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 27.350 61.240 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 26.920 61.240 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 26.490 61.240 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 26.060 61.240 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 25.630 61.240 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 25.200 61.240 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 24.770 61.240 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 24.340 61.240 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 23.910 61.240 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 28.210 60.835 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 27.780 60.835 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 27.350 60.835 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 26.920 60.835 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 26.490 60.835 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 26.060 60.835 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 25.630 60.835 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 25.200 60.835 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 24.770 60.835 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 24.340 60.835 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 23.910 60.835 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 28.210 60.430 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 27.780 60.430 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 27.350 60.430 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 26.920 60.430 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 26.490 60.430 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 26.060 60.430 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 25.630 60.430 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 25.200 60.430 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 24.770 60.430 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 24.340 60.430 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 23.910 60.430 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 28.210 60.025 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 27.780 60.025 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 27.350 60.025 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 26.920 60.025 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 26.490 60.025 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 26.060 60.025 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 25.630 60.025 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 25.200 60.025 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 24.770 60.025 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 24.340 60.025 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 23.910 60.025 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 28.210 59.620 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 27.780 59.620 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 27.350 59.620 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 26.920 59.620 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 26.490 59.620 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 26.060 59.620 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 25.630 59.620 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 25.200 59.620 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 24.770 59.620 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 24.340 59.620 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 23.910 59.620 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 28.210 59.215 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 27.780 59.215 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 27.350 59.215 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 26.920 59.215 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 26.490 59.215 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 26.060 59.215 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 25.630 59.215 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 25.200 59.215 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 24.770 59.215 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 24.340 59.215 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 23.910 59.215 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 28.210 58.810 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 27.780 58.810 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 27.350 58.810 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 26.920 58.810 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 26.490 58.810 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 26.060 58.810 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 25.630 58.810 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 25.200 58.810 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 24.770 58.810 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 24.340 58.810 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 23.910 58.810 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 28.210 58.405 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 27.780 58.405 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 27.350 58.405 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 26.920 58.405 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 26.490 58.405 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 26.060 58.405 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 25.630 58.405 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 25.200 58.405 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 24.770 58.405 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 24.340 58.405 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 23.910 58.405 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 28.210 58.000 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 27.780 58.000 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 27.350 58.000 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 26.920 58.000 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 26.490 58.000 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 26.060 58.000 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 25.630 58.000 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 25.200 58.000 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 24.770 58.000 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 24.340 58.000 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 23.910 58.000 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 28.210 57.595 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 27.780 57.595 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 27.350 57.595 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 26.920 57.595 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 26.490 57.595 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 26.060 57.595 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 25.630 57.595 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 25.200 57.595 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 24.770 57.595 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 24.340 57.595 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 23.910 57.595 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 28.210 57.190 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 27.780 57.190 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 27.350 57.190 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 26.920 57.190 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 26.490 57.190 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 26.060 57.190 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 25.630 57.190 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 25.200 57.190 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 24.770 57.190 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 24.340 57.190 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 23.910 57.190 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 28.210 56.785 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 27.780 56.785 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 27.350 56.785 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 26.920 56.785 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 26.490 56.785 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 26.060 56.785 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 25.630 56.785 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 25.200 56.785 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 24.770 56.785 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 24.340 56.785 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 23.910 56.785 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 28.210 56.375 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 27.780 56.375 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 27.350 56.375 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 26.920 56.375 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 26.490 56.375 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 26.060 56.375 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 25.630 56.375 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 25.200 56.375 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 24.770 56.375 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 24.340 56.375 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 23.910 56.375 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 28.210 55.965 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 27.780 55.965 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 27.350 55.965 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 26.920 55.965 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 26.490 55.965 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 26.060 55.965 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 25.630 55.965 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 25.200 55.965 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 24.770 55.965 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 24.340 55.965 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 23.910 55.965 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 28.210 55.555 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 27.780 55.555 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 27.350 55.555 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 26.920 55.555 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 26.490 55.555 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 26.060 55.555 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 25.630 55.555 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 25.200 55.555 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 24.770 55.555 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 24.340 55.555 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 23.910 55.555 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 28.210 55.145 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 27.780 55.145 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 27.350 55.145 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 26.920 55.145 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 26.490 55.145 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 26.060 55.145 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 25.630 55.145 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 25.200 55.145 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 24.770 55.145 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 24.340 55.145 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 23.910 55.145 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 28.210 54.735 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 27.780 54.735 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 27.350 54.735 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 26.920 54.735 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 26.490 54.735 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 26.060 54.735 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 25.630 54.735 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 25.200 54.735 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 24.770 54.735 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 24.340 54.735 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 23.910 54.735 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 28.210 54.325 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 27.780 54.325 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 27.350 54.325 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 26.920 54.325 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 26.490 54.325 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 26.060 54.325 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 25.630 54.325 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 25.200 54.325 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 24.770 54.325 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 24.340 54.325 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 23.910 54.325 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 28.210 53.915 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 27.780 53.915 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 27.350 53.915 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 26.920 53.915 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 26.490 53.915 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 26.060 53.915 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 25.630 53.915 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 25.200 53.915 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 24.770 53.915 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 24.340 53.915 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 23.910 53.915 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 28.210 53.505 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 27.780 53.505 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 27.350 53.505 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 26.920 53.505 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 26.490 53.505 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 26.060 53.505 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 25.630 53.505 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 25.200 53.505 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 24.770 53.505 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 24.340 53.505 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 23.910 53.505 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 28.210 53.095 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 27.780 53.095 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 27.350 53.095 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 26.920 53.095 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 26.490 53.095 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 26.060 53.095 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 25.630 53.095 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 25.200 53.095 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 24.770 53.095 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 24.340 53.095 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 23.910 53.095 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 28.210 52.685 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 27.780 52.685 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 27.350 52.685 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 26.920 52.685 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 26.490 52.685 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 26.060 52.685 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 25.630 52.685 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 25.200 52.685 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 24.770 52.685 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 24.340 52.685 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 23.910 52.685 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 28.210 52.275 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 27.780 52.275 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 27.350 52.275 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 26.920 52.275 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 26.490 52.275 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 26.060 52.275 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 25.630 52.275 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 25.200 52.275 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 24.770 52.275 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 24.340 52.275 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 23.910 52.275 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 28.210 51.865 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 27.780 51.865 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 27.350 51.865 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 26.920 51.865 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 26.490 51.865 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 26.060 51.865 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 25.630 51.865 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 25.200 51.865 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 24.770 51.865 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 24.340 51.865 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 23.910 51.865 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 28.210 51.455 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 27.780 51.455 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 27.350 51.455 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 26.920 51.455 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 26.490 51.455 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 26.060 51.455 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 25.630 51.455 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 25.200 51.455 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 24.770 51.455 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 24.340 51.455 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 23.910 51.455 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 28.210 51.045 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 27.780 51.045 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 27.350 51.045 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 26.920 51.045 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 26.490 51.045 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 26.060 51.045 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 25.630 51.045 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 25.200 51.045 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 24.770 51.045 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 24.340 51.045 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 23.910 51.045 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 28.210 24.310 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 27.780 24.310 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 27.350 24.310 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 26.920 24.310 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 26.490 24.310 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 26.060 24.310 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 25.630 24.310 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 25.200 24.310 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 24.770 24.310 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 24.340 24.310 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.110 23.910 24.310 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 28.210 23.905 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 27.780 23.905 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 27.350 23.905 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 26.920 23.905 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 26.490 23.905 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 26.060 23.905 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 25.630 23.905 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 25.200 23.905 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 24.770 23.905 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 24.340 23.905 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.705 23.910 23.905 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 28.210 23.500 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 27.780 23.500 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 27.350 23.500 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 26.920 23.500 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 26.490 23.500 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 26.060 23.500 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 25.630 23.500 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 25.200 23.500 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 24.770 23.500 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 24.340 23.500 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.300 23.910 23.500 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 28.210 23.095 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 27.780 23.095 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 27.350 23.095 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 26.920 23.095 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 26.490 23.095 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 26.060 23.095 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 25.630 23.095 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 25.200 23.095 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 24.770 23.095 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 24.340 23.095 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.895 23.910 23.095 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 28.210 22.690 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 27.780 22.690 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 27.350 22.690 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 26.920 22.690 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 26.490 22.690 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 26.060 22.690 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 25.630 22.690 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 25.200 22.690 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 24.770 22.690 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 24.340 22.690 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.490 23.910 22.690 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 28.210 22.285 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 27.780 22.285 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 27.350 22.285 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 26.920 22.285 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 26.490 22.285 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 26.060 22.285 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 25.630 22.285 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 25.200 22.285 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 24.770 22.285 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 24.340 22.285 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.085 23.910 22.285 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 28.210 21.880 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 27.780 21.880 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 27.350 21.880 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 26.920 21.880 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 26.490 21.880 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 26.060 21.880 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 25.630 21.880 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 25.200 21.880 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 24.770 21.880 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 24.340 21.880 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.680 23.910 21.880 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 28.210 21.475 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 27.780 21.475 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 27.350 21.475 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 26.920 21.475 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 26.490 21.475 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 26.060 21.475 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 25.630 21.475 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 25.200 21.475 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 24.770 21.475 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 24.340 21.475 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.275 23.910 21.475 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 28.210 21.070 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 27.780 21.070 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 27.350 21.070 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 26.920 21.070 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 26.490 21.070 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 26.060 21.070 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 25.630 21.070 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 25.200 21.070 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 24.770 21.070 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 24.340 21.070 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.870 23.910 21.070 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 28.210 20.665 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 27.780 20.665 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 27.350 20.665 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 26.920 20.665 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 26.490 20.665 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 26.060 20.665 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 25.630 20.665 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 25.200 20.665 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 24.770 20.665 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 24.340 20.665 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.465 23.910 20.665 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 28.210 20.260 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 27.780 20.260 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 27.350 20.260 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 26.920 20.260 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 26.490 20.260 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 26.060 20.260 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 25.630 20.260 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 25.200 20.260 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 24.770 20.260 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 24.340 20.260 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.060 23.910 20.260 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 28.210 19.855 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 27.780 19.855 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 27.350 19.855 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 26.920 19.855 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 26.490 19.855 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 26.060 19.855 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 25.630 19.855 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 25.200 19.855 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 24.770 19.855 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 24.340 19.855 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.655 23.910 19.855 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 28.210 19.450 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 27.780 19.450 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 27.350 19.450 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 26.920 19.450 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 26.490 19.450 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 26.060 19.450 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 25.630 19.450 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 25.200 19.450 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 24.770 19.450 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 24.340 19.450 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.250 23.910 19.450 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 28.210 19.045 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 27.780 19.045 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 27.350 19.045 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 26.920 19.045 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 26.490 19.045 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 26.060 19.045 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 25.630 19.045 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 25.200 19.045 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 24.770 19.045 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 24.340 19.045 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.845 23.910 19.045 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 28.210 18.640 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 27.780 18.640 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 27.350 18.640 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 26.920 18.640 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 26.490 18.640 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 26.060 18.640 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 25.630 18.640 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 25.200 18.640 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 24.770 18.640 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 24.340 18.640 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.440 23.910 18.640 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 28.210 18.235 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 27.780 18.235 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 27.350 18.235 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 26.920 18.235 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 26.490 18.235 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 26.060 18.235 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 25.630 18.235 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 25.200 18.235 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 24.770 18.235 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 24.340 18.235 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.035 23.910 18.235 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 28.210 17.830 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 27.780 17.830 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 27.350 17.830 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 26.920 17.830 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 26.490 17.830 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 26.060 17.830 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 25.630 17.830 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 25.200 17.830 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 24.770 17.830 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 24.340 17.830 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.630 23.910 17.830 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 28.210 17.425 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 27.780 17.425 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 27.350 17.425 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 26.920 17.425 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 26.490 17.425 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 26.060 17.425 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 25.630 17.425 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 25.200 17.425 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 24.770 17.425 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 24.340 17.425 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.225 23.910 17.425 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 28.210 17.020 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 27.780 17.020 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 27.350 17.020 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 26.920 17.020 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 26.490 17.020 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 26.060 17.020 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 25.630 17.020 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 25.200 17.020 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 24.770 17.020 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 24.340 17.020 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.820 23.910 17.020 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 28.210 16.615 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 27.780 16.615 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 27.350 16.615 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 26.920 16.615 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 26.490 16.615 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 26.060 16.615 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 25.630 16.615 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 25.200 16.615 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 24.770 16.615 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 24.340 16.615 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.415 23.910 16.615 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 28.210 16.210 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 27.780 16.210 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 27.350 16.210 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 26.920 16.210 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 26.490 16.210 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 26.060 16.210 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 25.630 16.210 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 25.200 16.210 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 24.770 16.210 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 24.340 16.210 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.010 23.910 16.210 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 28.210 15.805 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 27.780 15.805 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 27.350 15.805 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 26.920 15.805 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 26.490 15.805 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 26.060 15.805 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 25.630 15.805 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 25.200 15.805 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 24.770 15.805 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 24.340 15.805 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.605 23.910 15.805 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 28.210 15.400 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 27.780 15.400 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 27.350 15.400 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 26.920 15.400 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 26.490 15.400 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 26.060 15.400 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 25.630 15.400 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 25.200 15.400 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 24.770 15.400 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 24.340 15.400 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.200 23.910 15.400 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 28.210 14.995 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 27.780 14.995 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 27.350 14.995 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 26.920 14.995 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 26.490 14.995 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 26.060 14.995 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 25.630 14.995 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 25.200 14.995 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 24.770 14.995 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 24.340 14.995 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 23.910 14.995 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 28.210 14.590 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 27.780 14.590 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 27.350 14.590 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 26.920 14.590 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 26.490 14.590 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 26.060 14.590 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 25.630 14.590 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 25.200 14.590 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 24.770 14.590 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 24.340 14.590 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.390 23.910 14.590 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 28.210 14.185 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 27.780 14.185 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 27.350 14.185 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 26.920 14.185 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 26.490 14.185 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 26.060 14.185 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 25.630 14.185 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 25.200 14.185 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 24.770 14.185 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 24.340 14.185 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.985 23.910 14.185 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 28.210 13.780 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 27.780 13.780 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 27.350 13.780 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 26.920 13.780 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 26.490 13.780 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 26.060 13.780 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 25.630 13.780 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 25.200 13.780 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 24.770 13.780 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 24.340 13.780 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.580 23.910 13.780 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 28.210 13.375 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 27.780 13.375 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 27.350 13.375 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 26.920 13.375 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 26.490 13.375 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 26.060 13.375 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 25.630 13.375 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 25.200 13.375 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 24.770 13.375 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 24.340 13.375 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.175 23.910 13.375 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 28.210 12.970 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 27.780 12.970 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 27.350 12.970 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 26.920 12.970 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 26.490 12.970 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 26.060 12.970 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 25.630 12.970 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 25.200 12.970 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 24.770 12.970 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 24.340 12.970 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.770 23.910 12.970 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 197.645 12.875 197.965 ;
      LAYER met4 ;
        RECT 12.555 197.645 12.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 197.240 12.875 197.560 ;
      LAYER met4 ;
        RECT 12.555 197.240 12.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 196.835 12.875 197.155 ;
      LAYER met4 ;
        RECT 12.555 196.835 12.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 196.430 12.875 196.750 ;
      LAYER met4 ;
        RECT 12.555 196.430 12.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 196.025 12.875 196.345 ;
      LAYER met4 ;
        RECT 12.555 196.025 12.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 195.620 12.875 195.940 ;
      LAYER met4 ;
        RECT 12.555 195.620 12.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 195.215 12.875 195.535 ;
      LAYER met4 ;
        RECT 12.555 195.215 12.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 194.810 12.875 195.130 ;
      LAYER met4 ;
        RECT 12.555 194.810 12.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 194.405 12.875 194.725 ;
      LAYER met4 ;
        RECT 12.555 194.405 12.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 194.000 12.875 194.320 ;
      LAYER met4 ;
        RECT 12.555 194.000 12.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 193.595 12.875 193.915 ;
      LAYER met4 ;
        RECT 12.555 193.595 12.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 193.190 12.875 193.510 ;
      LAYER met4 ;
        RECT 12.555 193.190 12.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 192.785 12.875 193.105 ;
      LAYER met4 ;
        RECT 12.555 192.785 12.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 192.380 12.875 192.700 ;
      LAYER met4 ;
        RECT 12.555 192.380 12.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 191.975 12.875 192.295 ;
      LAYER met4 ;
        RECT 12.555 191.975 12.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 191.570 12.875 191.890 ;
      LAYER met4 ;
        RECT 12.555 191.570 12.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 191.165 12.875 191.485 ;
      LAYER met4 ;
        RECT 12.555 191.165 12.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 190.760 12.875 191.080 ;
      LAYER met4 ;
        RECT 12.555 190.760 12.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 190.355 12.875 190.675 ;
      LAYER met4 ;
        RECT 12.555 190.355 12.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 189.950 12.875 190.270 ;
      LAYER met4 ;
        RECT 12.555 189.950 12.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 189.545 12.875 189.865 ;
      LAYER met4 ;
        RECT 12.555 189.545 12.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 189.140 12.875 189.460 ;
      LAYER met4 ;
        RECT 12.555 189.140 12.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 188.735 12.875 189.055 ;
      LAYER met4 ;
        RECT 12.555 188.735 12.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 188.330 12.875 188.650 ;
      LAYER met4 ;
        RECT 12.555 188.330 12.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 187.925 12.875 188.245 ;
      LAYER met4 ;
        RECT 12.555 187.925 12.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 187.520 12.875 187.840 ;
      LAYER met4 ;
        RECT 12.555 187.520 12.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 187.115 12.875 187.435 ;
      LAYER met4 ;
        RECT 12.555 187.115 12.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 186.710 12.875 187.030 ;
      LAYER met4 ;
        RECT 12.555 186.710 12.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 186.305 12.875 186.625 ;
      LAYER met4 ;
        RECT 12.555 186.305 12.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 185.900 12.875 186.220 ;
      LAYER met4 ;
        RECT 12.555 185.900 12.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 185.495 12.875 185.815 ;
      LAYER met4 ;
        RECT 12.555 185.495 12.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 185.090 12.875 185.410 ;
      LAYER met4 ;
        RECT 12.555 185.090 12.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 184.685 12.875 185.005 ;
      LAYER met4 ;
        RECT 12.555 184.685 12.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 184.280 12.875 184.600 ;
      LAYER met4 ;
        RECT 12.555 184.280 12.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 183.875 12.875 184.195 ;
      LAYER met4 ;
        RECT 12.555 183.875 12.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 183.470 12.875 183.790 ;
      LAYER met4 ;
        RECT 12.555 183.470 12.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 183.065 12.875 183.385 ;
      LAYER met4 ;
        RECT 12.555 183.065 12.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 182.660 12.875 182.980 ;
      LAYER met4 ;
        RECT 12.555 182.660 12.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 182.255 12.875 182.575 ;
      LAYER met4 ;
        RECT 12.555 182.255 12.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 181.850 12.875 182.170 ;
      LAYER met4 ;
        RECT 12.555 181.850 12.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.555 181.445 12.875 181.765 ;
      LAYER met4 ;
        RECT 12.555 181.445 12.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 173.840 12.875 181.360 ;
      LAYER met4 ;
        RECT 1.270 173.840 12.875 181.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 28.210 12.565 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 27.780 12.565 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 27.350 12.565 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 26.920 12.565 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 26.490 12.565 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 26.060 12.565 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 25.630 12.565 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 25.200 12.565 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 24.770 12.565 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 24.340 12.565 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.365 23.910 12.565 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 197.645 12.475 197.965 ;
      LAYER met4 ;
        RECT 12.155 197.645 12.475 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 197.240 12.475 197.560 ;
      LAYER met4 ;
        RECT 12.155 197.240 12.475 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 196.835 12.475 197.155 ;
      LAYER met4 ;
        RECT 12.155 196.835 12.475 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 196.430 12.475 196.750 ;
      LAYER met4 ;
        RECT 12.155 196.430 12.475 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 196.025 12.475 196.345 ;
      LAYER met4 ;
        RECT 12.155 196.025 12.475 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 195.620 12.475 195.940 ;
      LAYER met4 ;
        RECT 12.155 195.620 12.475 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 195.215 12.475 195.535 ;
      LAYER met4 ;
        RECT 12.155 195.215 12.475 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 194.810 12.475 195.130 ;
      LAYER met4 ;
        RECT 12.155 194.810 12.475 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 194.405 12.475 194.725 ;
      LAYER met4 ;
        RECT 12.155 194.405 12.475 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 194.000 12.475 194.320 ;
      LAYER met4 ;
        RECT 12.155 194.000 12.475 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 193.595 12.475 193.915 ;
      LAYER met4 ;
        RECT 12.155 193.595 12.475 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 193.190 12.475 193.510 ;
      LAYER met4 ;
        RECT 12.155 193.190 12.475 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 192.785 12.475 193.105 ;
      LAYER met4 ;
        RECT 12.155 192.785 12.475 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 192.380 12.475 192.700 ;
      LAYER met4 ;
        RECT 12.155 192.380 12.475 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 191.975 12.475 192.295 ;
      LAYER met4 ;
        RECT 12.155 191.975 12.475 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 191.570 12.475 191.890 ;
      LAYER met4 ;
        RECT 12.155 191.570 12.475 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 191.165 12.475 191.485 ;
      LAYER met4 ;
        RECT 12.155 191.165 12.475 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 190.760 12.475 191.080 ;
      LAYER met4 ;
        RECT 12.155 190.760 12.475 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 190.355 12.475 190.675 ;
      LAYER met4 ;
        RECT 12.155 190.355 12.475 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 189.950 12.475 190.270 ;
      LAYER met4 ;
        RECT 12.155 189.950 12.475 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 189.545 12.475 189.865 ;
      LAYER met4 ;
        RECT 12.155 189.545 12.475 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 189.140 12.475 189.460 ;
      LAYER met4 ;
        RECT 12.155 189.140 12.475 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 188.735 12.475 189.055 ;
      LAYER met4 ;
        RECT 12.155 188.735 12.475 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 188.330 12.475 188.650 ;
      LAYER met4 ;
        RECT 12.155 188.330 12.475 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 187.925 12.475 188.245 ;
      LAYER met4 ;
        RECT 12.155 187.925 12.475 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 187.520 12.475 187.840 ;
      LAYER met4 ;
        RECT 12.155 187.520 12.475 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 187.115 12.475 187.435 ;
      LAYER met4 ;
        RECT 12.155 187.115 12.475 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 186.710 12.475 187.030 ;
      LAYER met4 ;
        RECT 12.155 186.710 12.475 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 186.305 12.475 186.625 ;
      LAYER met4 ;
        RECT 12.155 186.305 12.475 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 185.900 12.475 186.220 ;
      LAYER met4 ;
        RECT 12.155 185.900 12.475 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 185.495 12.475 185.815 ;
      LAYER met4 ;
        RECT 12.155 185.495 12.475 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 185.090 12.475 185.410 ;
      LAYER met4 ;
        RECT 12.155 185.090 12.475 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 184.685 12.475 185.005 ;
      LAYER met4 ;
        RECT 12.155 184.685 12.475 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 184.280 12.475 184.600 ;
      LAYER met4 ;
        RECT 12.155 184.280 12.475 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 183.875 12.475 184.195 ;
      LAYER met4 ;
        RECT 12.155 183.875 12.475 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 183.470 12.475 183.790 ;
      LAYER met4 ;
        RECT 12.155 183.470 12.475 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 183.065 12.475 183.385 ;
      LAYER met4 ;
        RECT 12.155 183.065 12.475 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 182.660 12.475 182.980 ;
      LAYER met4 ;
        RECT 12.155 182.660 12.475 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 182.255 12.475 182.575 ;
      LAYER met4 ;
        RECT 12.155 182.255 12.475 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 181.850 12.475 182.170 ;
      LAYER met4 ;
        RECT 12.155 181.850 12.475 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.155 181.445 12.475 181.765 ;
      LAYER met4 ;
        RECT 12.155 181.445 12.475 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 28.210 12.160 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 27.780 12.160 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 27.350 12.160 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 26.920 12.160 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 26.490 12.160 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 26.060 12.160 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 25.630 12.160 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 25.200 12.160 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 24.770 12.160 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 24.340 12.160 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.960 23.910 12.160 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 197.645 12.075 197.965 ;
      LAYER met4 ;
        RECT 11.755 197.645 12.075 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 197.240 12.075 197.560 ;
      LAYER met4 ;
        RECT 11.755 197.240 12.075 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 196.835 12.075 197.155 ;
      LAYER met4 ;
        RECT 11.755 196.835 12.075 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 196.430 12.075 196.750 ;
      LAYER met4 ;
        RECT 11.755 196.430 12.075 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 196.025 12.075 196.345 ;
      LAYER met4 ;
        RECT 11.755 196.025 12.075 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 195.620 12.075 195.940 ;
      LAYER met4 ;
        RECT 11.755 195.620 12.075 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 195.215 12.075 195.535 ;
      LAYER met4 ;
        RECT 11.755 195.215 12.075 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 194.810 12.075 195.130 ;
      LAYER met4 ;
        RECT 11.755 194.810 12.075 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 194.405 12.075 194.725 ;
      LAYER met4 ;
        RECT 11.755 194.405 12.075 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 194.000 12.075 194.320 ;
      LAYER met4 ;
        RECT 11.755 194.000 12.075 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 193.595 12.075 193.915 ;
      LAYER met4 ;
        RECT 11.755 193.595 12.075 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 193.190 12.075 193.510 ;
      LAYER met4 ;
        RECT 11.755 193.190 12.075 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 192.785 12.075 193.105 ;
      LAYER met4 ;
        RECT 11.755 192.785 12.075 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 192.380 12.075 192.700 ;
      LAYER met4 ;
        RECT 11.755 192.380 12.075 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 191.975 12.075 192.295 ;
      LAYER met4 ;
        RECT 11.755 191.975 12.075 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 191.570 12.075 191.890 ;
      LAYER met4 ;
        RECT 11.755 191.570 12.075 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 191.165 12.075 191.485 ;
      LAYER met4 ;
        RECT 11.755 191.165 12.075 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 190.760 12.075 191.080 ;
      LAYER met4 ;
        RECT 11.755 190.760 12.075 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 190.355 12.075 190.675 ;
      LAYER met4 ;
        RECT 11.755 190.355 12.075 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 189.950 12.075 190.270 ;
      LAYER met4 ;
        RECT 11.755 189.950 12.075 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 189.545 12.075 189.865 ;
      LAYER met4 ;
        RECT 11.755 189.545 12.075 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 189.140 12.075 189.460 ;
      LAYER met4 ;
        RECT 11.755 189.140 12.075 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 188.735 12.075 189.055 ;
      LAYER met4 ;
        RECT 11.755 188.735 12.075 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 188.330 12.075 188.650 ;
      LAYER met4 ;
        RECT 11.755 188.330 12.075 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 187.925 12.075 188.245 ;
      LAYER met4 ;
        RECT 11.755 187.925 12.075 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 187.520 12.075 187.840 ;
      LAYER met4 ;
        RECT 11.755 187.520 12.075 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 187.115 12.075 187.435 ;
      LAYER met4 ;
        RECT 11.755 187.115 12.075 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 186.710 12.075 187.030 ;
      LAYER met4 ;
        RECT 11.755 186.710 12.075 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 186.305 12.075 186.625 ;
      LAYER met4 ;
        RECT 11.755 186.305 12.075 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 185.900 12.075 186.220 ;
      LAYER met4 ;
        RECT 11.755 185.900 12.075 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 185.495 12.075 185.815 ;
      LAYER met4 ;
        RECT 11.755 185.495 12.075 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 185.090 12.075 185.410 ;
      LAYER met4 ;
        RECT 11.755 185.090 12.075 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 184.685 12.075 185.005 ;
      LAYER met4 ;
        RECT 11.755 184.685 12.075 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 184.280 12.075 184.600 ;
      LAYER met4 ;
        RECT 11.755 184.280 12.075 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 183.875 12.075 184.195 ;
      LAYER met4 ;
        RECT 11.755 183.875 12.075 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 183.470 12.075 183.790 ;
      LAYER met4 ;
        RECT 11.755 183.470 12.075 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 183.065 12.075 183.385 ;
      LAYER met4 ;
        RECT 11.755 183.065 12.075 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 182.660 12.075 182.980 ;
      LAYER met4 ;
        RECT 11.755 182.660 12.075 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 182.255 12.075 182.575 ;
      LAYER met4 ;
        RECT 11.755 182.255 12.075 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 181.850 12.075 182.170 ;
      LAYER met4 ;
        RECT 11.755 181.850 12.075 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.755 181.445 12.075 181.765 ;
      LAYER met4 ;
        RECT 11.755 181.445 12.075 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 28.210 11.755 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 27.780 11.755 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 27.350 11.755 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 26.920 11.755 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 26.490 11.755 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 26.060 11.755 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 25.630 11.755 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 25.200 11.755 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 24.770 11.755 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 24.340 11.755 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.555 23.910 11.755 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 197.645 11.675 197.965 ;
      LAYER met4 ;
        RECT 11.355 197.645 11.675 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 197.240 11.675 197.560 ;
      LAYER met4 ;
        RECT 11.355 197.240 11.675 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 196.835 11.675 197.155 ;
      LAYER met4 ;
        RECT 11.355 196.835 11.675 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 196.430 11.675 196.750 ;
      LAYER met4 ;
        RECT 11.355 196.430 11.675 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 196.025 11.675 196.345 ;
      LAYER met4 ;
        RECT 11.355 196.025 11.675 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 195.620 11.675 195.940 ;
      LAYER met4 ;
        RECT 11.355 195.620 11.675 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 195.215 11.675 195.535 ;
      LAYER met4 ;
        RECT 11.355 195.215 11.675 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 194.810 11.675 195.130 ;
      LAYER met4 ;
        RECT 11.355 194.810 11.675 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 194.405 11.675 194.725 ;
      LAYER met4 ;
        RECT 11.355 194.405 11.675 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 194.000 11.675 194.320 ;
      LAYER met4 ;
        RECT 11.355 194.000 11.675 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 193.595 11.675 193.915 ;
      LAYER met4 ;
        RECT 11.355 193.595 11.675 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 193.190 11.675 193.510 ;
      LAYER met4 ;
        RECT 11.355 193.190 11.675 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 192.785 11.675 193.105 ;
      LAYER met4 ;
        RECT 11.355 192.785 11.675 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 192.380 11.675 192.700 ;
      LAYER met4 ;
        RECT 11.355 192.380 11.675 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 191.975 11.675 192.295 ;
      LAYER met4 ;
        RECT 11.355 191.975 11.675 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 191.570 11.675 191.890 ;
      LAYER met4 ;
        RECT 11.355 191.570 11.675 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 191.165 11.675 191.485 ;
      LAYER met4 ;
        RECT 11.355 191.165 11.675 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 190.760 11.675 191.080 ;
      LAYER met4 ;
        RECT 11.355 190.760 11.675 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 190.355 11.675 190.675 ;
      LAYER met4 ;
        RECT 11.355 190.355 11.675 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 189.950 11.675 190.270 ;
      LAYER met4 ;
        RECT 11.355 189.950 11.675 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 189.545 11.675 189.865 ;
      LAYER met4 ;
        RECT 11.355 189.545 11.675 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 189.140 11.675 189.460 ;
      LAYER met4 ;
        RECT 11.355 189.140 11.675 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 188.735 11.675 189.055 ;
      LAYER met4 ;
        RECT 11.355 188.735 11.675 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 188.330 11.675 188.650 ;
      LAYER met4 ;
        RECT 11.355 188.330 11.675 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 187.925 11.675 188.245 ;
      LAYER met4 ;
        RECT 11.355 187.925 11.675 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 187.520 11.675 187.840 ;
      LAYER met4 ;
        RECT 11.355 187.520 11.675 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 187.115 11.675 187.435 ;
      LAYER met4 ;
        RECT 11.355 187.115 11.675 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 186.710 11.675 187.030 ;
      LAYER met4 ;
        RECT 11.355 186.710 11.675 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 186.305 11.675 186.625 ;
      LAYER met4 ;
        RECT 11.355 186.305 11.675 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 185.900 11.675 186.220 ;
      LAYER met4 ;
        RECT 11.355 185.900 11.675 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 185.495 11.675 185.815 ;
      LAYER met4 ;
        RECT 11.355 185.495 11.675 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 185.090 11.675 185.410 ;
      LAYER met4 ;
        RECT 11.355 185.090 11.675 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 184.685 11.675 185.005 ;
      LAYER met4 ;
        RECT 11.355 184.685 11.675 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 184.280 11.675 184.600 ;
      LAYER met4 ;
        RECT 11.355 184.280 11.675 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 183.875 11.675 184.195 ;
      LAYER met4 ;
        RECT 11.355 183.875 11.675 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 183.470 11.675 183.790 ;
      LAYER met4 ;
        RECT 11.355 183.470 11.675 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 183.065 11.675 183.385 ;
      LAYER met4 ;
        RECT 11.355 183.065 11.675 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 182.660 11.675 182.980 ;
      LAYER met4 ;
        RECT 11.355 182.660 11.675 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 182.255 11.675 182.575 ;
      LAYER met4 ;
        RECT 11.355 182.255 11.675 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 181.850 11.675 182.170 ;
      LAYER met4 ;
        RECT 11.355 181.850 11.675 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.355 181.445 11.675 181.765 ;
      LAYER met4 ;
        RECT 11.355 181.445 11.675 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 28.210 11.350 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 27.780 11.350 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 27.350 11.350 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 26.920 11.350 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 26.490 11.350 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 26.060 11.350 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 25.630 11.350 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 25.200 11.350 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 24.770 11.350 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 24.340 11.350 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.150 23.910 11.350 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 197.645 11.275 197.965 ;
      LAYER met4 ;
        RECT 10.955 197.645 11.275 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 197.240 11.275 197.560 ;
      LAYER met4 ;
        RECT 10.955 197.240 11.275 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 196.835 11.275 197.155 ;
      LAYER met4 ;
        RECT 10.955 196.835 11.275 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 196.430 11.275 196.750 ;
      LAYER met4 ;
        RECT 10.955 196.430 11.275 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 196.025 11.275 196.345 ;
      LAYER met4 ;
        RECT 10.955 196.025 11.275 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 195.620 11.275 195.940 ;
      LAYER met4 ;
        RECT 10.955 195.620 11.275 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 195.215 11.275 195.535 ;
      LAYER met4 ;
        RECT 10.955 195.215 11.275 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 194.810 11.275 195.130 ;
      LAYER met4 ;
        RECT 10.955 194.810 11.275 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 194.405 11.275 194.725 ;
      LAYER met4 ;
        RECT 10.955 194.405 11.275 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 194.000 11.275 194.320 ;
      LAYER met4 ;
        RECT 10.955 194.000 11.275 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 193.595 11.275 193.915 ;
      LAYER met4 ;
        RECT 10.955 193.595 11.275 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 193.190 11.275 193.510 ;
      LAYER met4 ;
        RECT 10.955 193.190 11.275 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 192.785 11.275 193.105 ;
      LAYER met4 ;
        RECT 10.955 192.785 11.275 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 192.380 11.275 192.700 ;
      LAYER met4 ;
        RECT 10.955 192.380 11.275 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 191.975 11.275 192.295 ;
      LAYER met4 ;
        RECT 10.955 191.975 11.275 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 191.570 11.275 191.890 ;
      LAYER met4 ;
        RECT 10.955 191.570 11.275 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 191.165 11.275 191.485 ;
      LAYER met4 ;
        RECT 10.955 191.165 11.275 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 190.760 11.275 191.080 ;
      LAYER met4 ;
        RECT 10.955 190.760 11.275 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 190.355 11.275 190.675 ;
      LAYER met4 ;
        RECT 10.955 190.355 11.275 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 189.950 11.275 190.270 ;
      LAYER met4 ;
        RECT 10.955 189.950 11.275 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 189.545 11.275 189.865 ;
      LAYER met4 ;
        RECT 10.955 189.545 11.275 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 189.140 11.275 189.460 ;
      LAYER met4 ;
        RECT 10.955 189.140 11.275 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 188.735 11.275 189.055 ;
      LAYER met4 ;
        RECT 10.955 188.735 11.275 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 188.330 11.275 188.650 ;
      LAYER met4 ;
        RECT 10.955 188.330 11.275 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 187.925 11.275 188.245 ;
      LAYER met4 ;
        RECT 10.955 187.925 11.275 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 187.520 11.275 187.840 ;
      LAYER met4 ;
        RECT 10.955 187.520 11.275 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 187.115 11.275 187.435 ;
      LAYER met4 ;
        RECT 10.955 187.115 11.275 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 186.710 11.275 187.030 ;
      LAYER met4 ;
        RECT 10.955 186.710 11.275 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 186.305 11.275 186.625 ;
      LAYER met4 ;
        RECT 10.955 186.305 11.275 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 185.900 11.275 186.220 ;
      LAYER met4 ;
        RECT 10.955 185.900 11.275 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 185.495 11.275 185.815 ;
      LAYER met4 ;
        RECT 10.955 185.495 11.275 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 185.090 11.275 185.410 ;
      LAYER met4 ;
        RECT 10.955 185.090 11.275 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 184.685 11.275 185.005 ;
      LAYER met4 ;
        RECT 10.955 184.685 11.275 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 184.280 11.275 184.600 ;
      LAYER met4 ;
        RECT 10.955 184.280 11.275 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 183.875 11.275 184.195 ;
      LAYER met4 ;
        RECT 10.955 183.875 11.275 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 183.470 11.275 183.790 ;
      LAYER met4 ;
        RECT 10.955 183.470 11.275 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 183.065 11.275 183.385 ;
      LAYER met4 ;
        RECT 10.955 183.065 11.275 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 182.660 11.275 182.980 ;
      LAYER met4 ;
        RECT 10.955 182.660 11.275 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 182.255 11.275 182.575 ;
      LAYER met4 ;
        RECT 10.955 182.255 11.275 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 181.850 11.275 182.170 ;
      LAYER met4 ;
        RECT 10.955 181.850 11.275 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.955 181.445 11.275 181.765 ;
      LAYER met4 ;
        RECT 10.955 181.445 11.275 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 28.210 10.945 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 27.780 10.945 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 27.350 10.945 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 26.920 10.945 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 26.490 10.945 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 26.060 10.945 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 25.630 10.945 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 25.200 10.945 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 24.770 10.945 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 24.340 10.945 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.745 23.910 10.945 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 197.645 10.875 197.965 ;
      LAYER met4 ;
        RECT 10.555 197.645 10.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 197.240 10.875 197.560 ;
      LAYER met4 ;
        RECT 10.555 197.240 10.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 196.835 10.875 197.155 ;
      LAYER met4 ;
        RECT 10.555 196.835 10.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 196.430 10.875 196.750 ;
      LAYER met4 ;
        RECT 10.555 196.430 10.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 196.025 10.875 196.345 ;
      LAYER met4 ;
        RECT 10.555 196.025 10.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 195.620 10.875 195.940 ;
      LAYER met4 ;
        RECT 10.555 195.620 10.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 195.215 10.875 195.535 ;
      LAYER met4 ;
        RECT 10.555 195.215 10.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 194.810 10.875 195.130 ;
      LAYER met4 ;
        RECT 10.555 194.810 10.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 194.405 10.875 194.725 ;
      LAYER met4 ;
        RECT 10.555 194.405 10.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 194.000 10.875 194.320 ;
      LAYER met4 ;
        RECT 10.555 194.000 10.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 193.595 10.875 193.915 ;
      LAYER met4 ;
        RECT 10.555 193.595 10.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 193.190 10.875 193.510 ;
      LAYER met4 ;
        RECT 10.555 193.190 10.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 192.785 10.875 193.105 ;
      LAYER met4 ;
        RECT 10.555 192.785 10.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 192.380 10.875 192.700 ;
      LAYER met4 ;
        RECT 10.555 192.380 10.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 191.975 10.875 192.295 ;
      LAYER met4 ;
        RECT 10.555 191.975 10.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 191.570 10.875 191.890 ;
      LAYER met4 ;
        RECT 10.555 191.570 10.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 191.165 10.875 191.485 ;
      LAYER met4 ;
        RECT 10.555 191.165 10.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 190.760 10.875 191.080 ;
      LAYER met4 ;
        RECT 10.555 190.760 10.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 190.355 10.875 190.675 ;
      LAYER met4 ;
        RECT 10.555 190.355 10.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 189.950 10.875 190.270 ;
      LAYER met4 ;
        RECT 10.555 189.950 10.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 189.545 10.875 189.865 ;
      LAYER met4 ;
        RECT 10.555 189.545 10.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 189.140 10.875 189.460 ;
      LAYER met4 ;
        RECT 10.555 189.140 10.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 188.735 10.875 189.055 ;
      LAYER met4 ;
        RECT 10.555 188.735 10.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 188.330 10.875 188.650 ;
      LAYER met4 ;
        RECT 10.555 188.330 10.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 187.925 10.875 188.245 ;
      LAYER met4 ;
        RECT 10.555 187.925 10.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 187.520 10.875 187.840 ;
      LAYER met4 ;
        RECT 10.555 187.520 10.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 187.115 10.875 187.435 ;
      LAYER met4 ;
        RECT 10.555 187.115 10.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 186.710 10.875 187.030 ;
      LAYER met4 ;
        RECT 10.555 186.710 10.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 186.305 10.875 186.625 ;
      LAYER met4 ;
        RECT 10.555 186.305 10.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 185.900 10.875 186.220 ;
      LAYER met4 ;
        RECT 10.555 185.900 10.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 185.495 10.875 185.815 ;
      LAYER met4 ;
        RECT 10.555 185.495 10.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 185.090 10.875 185.410 ;
      LAYER met4 ;
        RECT 10.555 185.090 10.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 184.685 10.875 185.005 ;
      LAYER met4 ;
        RECT 10.555 184.685 10.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 184.280 10.875 184.600 ;
      LAYER met4 ;
        RECT 10.555 184.280 10.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 183.875 10.875 184.195 ;
      LAYER met4 ;
        RECT 10.555 183.875 10.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 183.470 10.875 183.790 ;
      LAYER met4 ;
        RECT 10.555 183.470 10.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 183.065 10.875 183.385 ;
      LAYER met4 ;
        RECT 10.555 183.065 10.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 182.660 10.875 182.980 ;
      LAYER met4 ;
        RECT 10.555 182.660 10.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 182.255 10.875 182.575 ;
      LAYER met4 ;
        RECT 10.555 182.255 10.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 181.850 10.875 182.170 ;
      LAYER met4 ;
        RECT 10.555 181.850 10.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.555 181.445 10.875 181.765 ;
      LAYER met4 ;
        RECT 10.555 181.445 10.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 28.210 10.540 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 27.780 10.540 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 27.350 10.540 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 26.920 10.540 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 26.490 10.540 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 26.060 10.540 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 25.630 10.540 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 25.200 10.540 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 24.770 10.540 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 24.340 10.540 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.340 23.910 10.540 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 197.645 10.475 197.965 ;
      LAYER met4 ;
        RECT 10.155 197.645 10.475 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 197.240 10.475 197.560 ;
      LAYER met4 ;
        RECT 10.155 197.240 10.475 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 196.835 10.475 197.155 ;
      LAYER met4 ;
        RECT 10.155 196.835 10.475 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 196.430 10.475 196.750 ;
      LAYER met4 ;
        RECT 10.155 196.430 10.475 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 196.025 10.475 196.345 ;
      LAYER met4 ;
        RECT 10.155 196.025 10.475 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 195.620 10.475 195.940 ;
      LAYER met4 ;
        RECT 10.155 195.620 10.475 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 195.215 10.475 195.535 ;
      LAYER met4 ;
        RECT 10.155 195.215 10.475 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 194.810 10.475 195.130 ;
      LAYER met4 ;
        RECT 10.155 194.810 10.475 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 194.405 10.475 194.725 ;
      LAYER met4 ;
        RECT 10.155 194.405 10.475 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 194.000 10.475 194.320 ;
      LAYER met4 ;
        RECT 10.155 194.000 10.475 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 193.595 10.475 193.915 ;
      LAYER met4 ;
        RECT 10.155 193.595 10.475 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 193.190 10.475 193.510 ;
      LAYER met4 ;
        RECT 10.155 193.190 10.475 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 192.785 10.475 193.105 ;
      LAYER met4 ;
        RECT 10.155 192.785 10.475 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 192.380 10.475 192.700 ;
      LAYER met4 ;
        RECT 10.155 192.380 10.475 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 191.975 10.475 192.295 ;
      LAYER met4 ;
        RECT 10.155 191.975 10.475 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 191.570 10.475 191.890 ;
      LAYER met4 ;
        RECT 10.155 191.570 10.475 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 191.165 10.475 191.485 ;
      LAYER met4 ;
        RECT 10.155 191.165 10.475 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 190.760 10.475 191.080 ;
      LAYER met4 ;
        RECT 10.155 190.760 10.475 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 190.355 10.475 190.675 ;
      LAYER met4 ;
        RECT 10.155 190.355 10.475 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 189.950 10.475 190.270 ;
      LAYER met4 ;
        RECT 10.155 189.950 10.475 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 189.545 10.475 189.865 ;
      LAYER met4 ;
        RECT 10.155 189.545 10.475 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 189.140 10.475 189.460 ;
      LAYER met4 ;
        RECT 10.155 189.140 10.475 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 188.735 10.475 189.055 ;
      LAYER met4 ;
        RECT 10.155 188.735 10.475 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 188.330 10.475 188.650 ;
      LAYER met4 ;
        RECT 10.155 188.330 10.475 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 187.925 10.475 188.245 ;
      LAYER met4 ;
        RECT 10.155 187.925 10.475 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 187.520 10.475 187.840 ;
      LAYER met4 ;
        RECT 10.155 187.520 10.475 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 187.115 10.475 187.435 ;
      LAYER met4 ;
        RECT 10.155 187.115 10.475 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 186.710 10.475 187.030 ;
      LAYER met4 ;
        RECT 10.155 186.710 10.475 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 186.305 10.475 186.625 ;
      LAYER met4 ;
        RECT 10.155 186.305 10.475 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 185.900 10.475 186.220 ;
      LAYER met4 ;
        RECT 10.155 185.900 10.475 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 185.495 10.475 185.815 ;
      LAYER met4 ;
        RECT 10.155 185.495 10.475 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 185.090 10.475 185.410 ;
      LAYER met4 ;
        RECT 10.155 185.090 10.475 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 184.685 10.475 185.005 ;
      LAYER met4 ;
        RECT 10.155 184.685 10.475 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 184.280 10.475 184.600 ;
      LAYER met4 ;
        RECT 10.155 184.280 10.475 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 183.875 10.475 184.195 ;
      LAYER met4 ;
        RECT 10.155 183.875 10.475 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 183.470 10.475 183.790 ;
      LAYER met4 ;
        RECT 10.155 183.470 10.475 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 183.065 10.475 183.385 ;
      LAYER met4 ;
        RECT 10.155 183.065 10.475 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 182.660 10.475 182.980 ;
      LAYER met4 ;
        RECT 10.155 182.660 10.475 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 182.255 10.475 182.575 ;
      LAYER met4 ;
        RECT 10.155 182.255 10.475 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 181.850 10.475 182.170 ;
      LAYER met4 ;
        RECT 10.155 181.850 10.475 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.155 181.445 10.475 181.765 ;
      LAYER met4 ;
        RECT 10.155 181.445 10.475 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 28.210 10.135 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 27.780 10.135 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 27.350 10.135 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 26.920 10.135 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 26.490 10.135 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 26.060 10.135 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 25.630 10.135 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 25.200 10.135 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 24.770 10.135 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 24.340 10.135 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.935 23.910 10.135 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 197.645 10.075 197.965 ;
      LAYER met4 ;
        RECT 9.755 197.645 10.075 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 197.240 10.075 197.560 ;
      LAYER met4 ;
        RECT 9.755 197.240 10.075 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 196.835 10.075 197.155 ;
      LAYER met4 ;
        RECT 9.755 196.835 10.075 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 196.430 10.075 196.750 ;
      LAYER met4 ;
        RECT 9.755 196.430 10.075 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 196.025 10.075 196.345 ;
      LAYER met4 ;
        RECT 9.755 196.025 10.075 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 195.620 10.075 195.940 ;
      LAYER met4 ;
        RECT 9.755 195.620 10.075 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 195.215 10.075 195.535 ;
      LAYER met4 ;
        RECT 9.755 195.215 10.075 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 194.810 10.075 195.130 ;
      LAYER met4 ;
        RECT 9.755 194.810 10.075 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 194.405 10.075 194.725 ;
      LAYER met4 ;
        RECT 9.755 194.405 10.075 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 194.000 10.075 194.320 ;
      LAYER met4 ;
        RECT 9.755 194.000 10.075 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 193.595 10.075 193.915 ;
      LAYER met4 ;
        RECT 9.755 193.595 10.075 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 193.190 10.075 193.510 ;
      LAYER met4 ;
        RECT 9.755 193.190 10.075 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 192.785 10.075 193.105 ;
      LAYER met4 ;
        RECT 9.755 192.785 10.075 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 192.380 10.075 192.700 ;
      LAYER met4 ;
        RECT 9.755 192.380 10.075 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 191.975 10.075 192.295 ;
      LAYER met4 ;
        RECT 9.755 191.975 10.075 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 191.570 10.075 191.890 ;
      LAYER met4 ;
        RECT 9.755 191.570 10.075 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 191.165 10.075 191.485 ;
      LAYER met4 ;
        RECT 9.755 191.165 10.075 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 190.760 10.075 191.080 ;
      LAYER met4 ;
        RECT 9.755 190.760 10.075 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 190.355 10.075 190.675 ;
      LAYER met4 ;
        RECT 9.755 190.355 10.075 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 189.950 10.075 190.270 ;
      LAYER met4 ;
        RECT 9.755 189.950 10.075 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 189.545 10.075 189.865 ;
      LAYER met4 ;
        RECT 9.755 189.545 10.075 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 189.140 10.075 189.460 ;
      LAYER met4 ;
        RECT 9.755 189.140 10.075 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 188.735 10.075 189.055 ;
      LAYER met4 ;
        RECT 9.755 188.735 10.075 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 188.330 10.075 188.650 ;
      LAYER met4 ;
        RECT 9.755 188.330 10.075 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 187.925 10.075 188.245 ;
      LAYER met4 ;
        RECT 9.755 187.925 10.075 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 187.520 10.075 187.840 ;
      LAYER met4 ;
        RECT 9.755 187.520 10.075 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 187.115 10.075 187.435 ;
      LAYER met4 ;
        RECT 9.755 187.115 10.075 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 186.710 10.075 187.030 ;
      LAYER met4 ;
        RECT 9.755 186.710 10.075 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 186.305 10.075 186.625 ;
      LAYER met4 ;
        RECT 9.755 186.305 10.075 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 185.900 10.075 186.220 ;
      LAYER met4 ;
        RECT 9.755 185.900 10.075 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 185.495 10.075 185.815 ;
      LAYER met4 ;
        RECT 9.755 185.495 10.075 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 185.090 10.075 185.410 ;
      LAYER met4 ;
        RECT 9.755 185.090 10.075 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 184.685 10.075 185.005 ;
      LAYER met4 ;
        RECT 9.755 184.685 10.075 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 184.280 10.075 184.600 ;
      LAYER met4 ;
        RECT 9.755 184.280 10.075 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 183.875 10.075 184.195 ;
      LAYER met4 ;
        RECT 9.755 183.875 10.075 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 183.470 10.075 183.790 ;
      LAYER met4 ;
        RECT 9.755 183.470 10.075 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 183.065 10.075 183.385 ;
      LAYER met4 ;
        RECT 9.755 183.065 10.075 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 182.660 10.075 182.980 ;
      LAYER met4 ;
        RECT 9.755 182.660 10.075 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 182.255 10.075 182.575 ;
      LAYER met4 ;
        RECT 9.755 182.255 10.075 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 181.850 10.075 182.170 ;
      LAYER met4 ;
        RECT 9.755 181.850 10.075 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.755 181.445 10.075 181.765 ;
      LAYER met4 ;
        RECT 9.755 181.445 10.075 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 28.210 9.730 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 27.780 9.730 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 27.350 9.730 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 26.920 9.730 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 26.490 9.730 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 26.060 9.730 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 25.630 9.730 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 25.200 9.730 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 24.770 9.730 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 24.340 9.730 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.530 23.910 9.730 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 197.645 9.675 197.965 ;
      LAYER met4 ;
        RECT 9.355 197.645 9.675 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 197.240 9.675 197.560 ;
      LAYER met4 ;
        RECT 9.355 197.240 9.675 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 196.835 9.675 197.155 ;
      LAYER met4 ;
        RECT 9.355 196.835 9.675 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 196.430 9.675 196.750 ;
      LAYER met4 ;
        RECT 9.355 196.430 9.675 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 196.025 9.675 196.345 ;
      LAYER met4 ;
        RECT 9.355 196.025 9.675 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 195.620 9.675 195.940 ;
      LAYER met4 ;
        RECT 9.355 195.620 9.675 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 195.215 9.675 195.535 ;
      LAYER met4 ;
        RECT 9.355 195.215 9.675 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 194.810 9.675 195.130 ;
      LAYER met4 ;
        RECT 9.355 194.810 9.675 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 194.405 9.675 194.725 ;
      LAYER met4 ;
        RECT 9.355 194.405 9.675 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 194.000 9.675 194.320 ;
      LAYER met4 ;
        RECT 9.355 194.000 9.675 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 193.595 9.675 193.915 ;
      LAYER met4 ;
        RECT 9.355 193.595 9.675 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 193.190 9.675 193.510 ;
      LAYER met4 ;
        RECT 9.355 193.190 9.675 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 192.785 9.675 193.105 ;
      LAYER met4 ;
        RECT 9.355 192.785 9.675 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 192.380 9.675 192.700 ;
      LAYER met4 ;
        RECT 9.355 192.380 9.675 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 191.975 9.675 192.295 ;
      LAYER met4 ;
        RECT 9.355 191.975 9.675 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 191.570 9.675 191.890 ;
      LAYER met4 ;
        RECT 9.355 191.570 9.675 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 191.165 9.675 191.485 ;
      LAYER met4 ;
        RECT 9.355 191.165 9.675 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 190.760 9.675 191.080 ;
      LAYER met4 ;
        RECT 9.355 190.760 9.675 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 190.355 9.675 190.675 ;
      LAYER met4 ;
        RECT 9.355 190.355 9.675 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 189.950 9.675 190.270 ;
      LAYER met4 ;
        RECT 9.355 189.950 9.675 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 189.545 9.675 189.865 ;
      LAYER met4 ;
        RECT 9.355 189.545 9.675 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 189.140 9.675 189.460 ;
      LAYER met4 ;
        RECT 9.355 189.140 9.675 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 188.735 9.675 189.055 ;
      LAYER met4 ;
        RECT 9.355 188.735 9.675 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 188.330 9.675 188.650 ;
      LAYER met4 ;
        RECT 9.355 188.330 9.675 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 187.925 9.675 188.245 ;
      LAYER met4 ;
        RECT 9.355 187.925 9.675 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 187.520 9.675 187.840 ;
      LAYER met4 ;
        RECT 9.355 187.520 9.675 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 187.115 9.675 187.435 ;
      LAYER met4 ;
        RECT 9.355 187.115 9.675 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 186.710 9.675 187.030 ;
      LAYER met4 ;
        RECT 9.355 186.710 9.675 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 186.305 9.675 186.625 ;
      LAYER met4 ;
        RECT 9.355 186.305 9.675 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 185.900 9.675 186.220 ;
      LAYER met4 ;
        RECT 9.355 185.900 9.675 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 185.495 9.675 185.815 ;
      LAYER met4 ;
        RECT 9.355 185.495 9.675 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 185.090 9.675 185.410 ;
      LAYER met4 ;
        RECT 9.355 185.090 9.675 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 184.685 9.675 185.005 ;
      LAYER met4 ;
        RECT 9.355 184.685 9.675 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 184.280 9.675 184.600 ;
      LAYER met4 ;
        RECT 9.355 184.280 9.675 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 183.875 9.675 184.195 ;
      LAYER met4 ;
        RECT 9.355 183.875 9.675 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 183.470 9.675 183.790 ;
      LAYER met4 ;
        RECT 9.355 183.470 9.675 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 183.065 9.675 183.385 ;
      LAYER met4 ;
        RECT 9.355 183.065 9.675 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 182.660 9.675 182.980 ;
      LAYER met4 ;
        RECT 9.355 182.660 9.675 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 182.255 9.675 182.575 ;
      LAYER met4 ;
        RECT 9.355 182.255 9.675 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 181.850 9.675 182.170 ;
      LAYER met4 ;
        RECT 9.355 181.850 9.675 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 181.445 9.675 181.765 ;
      LAYER met4 ;
        RECT 9.355 181.445 9.675 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 28.210 9.325 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 27.780 9.325 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 27.350 9.325 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 26.920 9.325 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 26.490 9.325 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 26.060 9.325 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 25.630 9.325 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 25.200 9.325 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 24.770 9.325 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 24.340 9.325 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.125 23.910 9.325 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 197.645 9.275 197.965 ;
      LAYER met4 ;
        RECT 8.955 197.645 9.275 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 197.240 9.275 197.560 ;
      LAYER met4 ;
        RECT 8.955 197.240 9.275 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 196.835 9.275 197.155 ;
      LAYER met4 ;
        RECT 8.955 196.835 9.275 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 196.430 9.275 196.750 ;
      LAYER met4 ;
        RECT 8.955 196.430 9.275 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 196.025 9.275 196.345 ;
      LAYER met4 ;
        RECT 8.955 196.025 9.275 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 195.620 9.275 195.940 ;
      LAYER met4 ;
        RECT 8.955 195.620 9.275 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 195.215 9.275 195.535 ;
      LAYER met4 ;
        RECT 8.955 195.215 9.275 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 194.810 9.275 195.130 ;
      LAYER met4 ;
        RECT 8.955 194.810 9.275 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 194.405 9.275 194.725 ;
      LAYER met4 ;
        RECT 8.955 194.405 9.275 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 194.000 9.275 194.320 ;
      LAYER met4 ;
        RECT 8.955 194.000 9.275 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 193.595 9.275 193.915 ;
      LAYER met4 ;
        RECT 8.955 193.595 9.275 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 193.190 9.275 193.510 ;
      LAYER met4 ;
        RECT 8.955 193.190 9.275 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 192.785 9.275 193.105 ;
      LAYER met4 ;
        RECT 8.955 192.785 9.275 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 192.380 9.275 192.700 ;
      LAYER met4 ;
        RECT 8.955 192.380 9.275 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 191.975 9.275 192.295 ;
      LAYER met4 ;
        RECT 8.955 191.975 9.275 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 191.570 9.275 191.890 ;
      LAYER met4 ;
        RECT 8.955 191.570 9.275 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 191.165 9.275 191.485 ;
      LAYER met4 ;
        RECT 8.955 191.165 9.275 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 190.760 9.275 191.080 ;
      LAYER met4 ;
        RECT 8.955 190.760 9.275 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 190.355 9.275 190.675 ;
      LAYER met4 ;
        RECT 8.955 190.355 9.275 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 189.950 9.275 190.270 ;
      LAYER met4 ;
        RECT 8.955 189.950 9.275 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 189.545 9.275 189.865 ;
      LAYER met4 ;
        RECT 8.955 189.545 9.275 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 189.140 9.275 189.460 ;
      LAYER met4 ;
        RECT 8.955 189.140 9.275 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 188.735 9.275 189.055 ;
      LAYER met4 ;
        RECT 8.955 188.735 9.275 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 188.330 9.275 188.650 ;
      LAYER met4 ;
        RECT 8.955 188.330 9.275 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 187.925 9.275 188.245 ;
      LAYER met4 ;
        RECT 8.955 187.925 9.275 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 187.520 9.275 187.840 ;
      LAYER met4 ;
        RECT 8.955 187.520 9.275 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 187.115 9.275 187.435 ;
      LAYER met4 ;
        RECT 8.955 187.115 9.275 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 186.710 9.275 187.030 ;
      LAYER met4 ;
        RECT 8.955 186.710 9.275 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 186.305 9.275 186.625 ;
      LAYER met4 ;
        RECT 8.955 186.305 9.275 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 185.900 9.275 186.220 ;
      LAYER met4 ;
        RECT 8.955 185.900 9.275 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 185.495 9.275 185.815 ;
      LAYER met4 ;
        RECT 8.955 185.495 9.275 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 185.090 9.275 185.410 ;
      LAYER met4 ;
        RECT 8.955 185.090 9.275 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 184.685 9.275 185.005 ;
      LAYER met4 ;
        RECT 8.955 184.685 9.275 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 184.280 9.275 184.600 ;
      LAYER met4 ;
        RECT 8.955 184.280 9.275 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 183.875 9.275 184.195 ;
      LAYER met4 ;
        RECT 8.955 183.875 9.275 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 183.470 9.275 183.790 ;
      LAYER met4 ;
        RECT 8.955 183.470 9.275 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 183.065 9.275 183.385 ;
      LAYER met4 ;
        RECT 8.955 183.065 9.275 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 182.660 9.275 182.980 ;
      LAYER met4 ;
        RECT 8.955 182.660 9.275 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 182.255 9.275 182.575 ;
      LAYER met4 ;
        RECT 8.955 182.255 9.275 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 181.850 9.275 182.170 ;
      LAYER met4 ;
        RECT 8.955 181.850 9.275 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.955 181.445 9.275 181.765 ;
      LAYER met4 ;
        RECT 8.955 181.445 9.275 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 28.210 8.920 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 27.780 8.920 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 27.350 8.920 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 26.920 8.920 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 26.490 8.920 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 26.060 8.920 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 25.630 8.920 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 25.200 8.920 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 24.770 8.920 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 24.340 8.920 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.720 23.910 8.920 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 197.645 8.875 197.965 ;
      LAYER met4 ;
        RECT 8.555 197.645 8.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 197.240 8.875 197.560 ;
      LAYER met4 ;
        RECT 8.555 197.240 8.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 196.835 8.875 197.155 ;
      LAYER met4 ;
        RECT 8.555 196.835 8.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 196.430 8.875 196.750 ;
      LAYER met4 ;
        RECT 8.555 196.430 8.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 196.025 8.875 196.345 ;
      LAYER met4 ;
        RECT 8.555 196.025 8.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 195.620 8.875 195.940 ;
      LAYER met4 ;
        RECT 8.555 195.620 8.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 195.215 8.875 195.535 ;
      LAYER met4 ;
        RECT 8.555 195.215 8.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 194.810 8.875 195.130 ;
      LAYER met4 ;
        RECT 8.555 194.810 8.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 194.405 8.875 194.725 ;
      LAYER met4 ;
        RECT 8.555 194.405 8.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 194.000 8.875 194.320 ;
      LAYER met4 ;
        RECT 8.555 194.000 8.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 193.595 8.875 193.915 ;
      LAYER met4 ;
        RECT 8.555 193.595 8.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 193.190 8.875 193.510 ;
      LAYER met4 ;
        RECT 8.555 193.190 8.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 192.785 8.875 193.105 ;
      LAYER met4 ;
        RECT 8.555 192.785 8.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 192.380 8.875 192.700 ;
      LAYER met4 ;
        RECT 8.555 192.380 8.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 191.975 8.875 192.295 ;
      LAYER met4 ;
        RECT 8.555 191.975 8.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 191.570 8.875 191.890 ;
      LAYER met4 ;
        RECT 8.555 191.570 8.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 191.165 8.875 191.485 ;
      LAYER met4 ;
        RECT 8.555 191.165 8.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 190.760 8.875 191.080 ;
      LAYER met4 ;
        RECT 8.555 190.760 8.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 190.355 8.875 190.675 ;
      LAYER met4 ;
        RECT 8.555 190.355 8.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 189.950 8.875 190.270 ;
      LAYER met4 ;
        RECT 8.555 189.950 8.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 189.545 8.875 189.865 ;
      LAYER met4 ;
        RECT 8.555 189.545 8.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 189.140 8.875 189.460 ;
      LAYER met4 ;
        RECT 8.555 189.140 8.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 188.735 8.875 189.055 ;
      LAYER met4 ;
        RECT 8.555 188.735 8.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 188.330 8.875 188.650 ;
      LAYER met4 ;
        RECT 8.555 188.330 8.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 187.925 8.875 188.245 ;
      LAYER met4 ;
        RECT 8.555 187.925 8.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 187.520 8.875 187.840 ;
      LAYER met4 ;
        RECT 8.555 187.520 8.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 187.115 8.875 187.435 ;
      LAYER met4 ;
        RECT 8.555 187.115 8.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 186.710 8.875 187.030 ;
      LAYER met4 ;
        RECT 8.555 186.710 8.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 186.305 8.875 186.625 ;
      LAYER met4 ;
        RECT 8.555 186.305 8.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 185.900 8.875 186.220 ;
      LAYER met4 ;
        RECT 8.555 185.900 8.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 185.495 8.875 185.815 ;
      LAYER met4 ;
        RECT 8.555 185.495 8.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 185.090 8.875 185.410 ;
      LAYER met4 ;
        RECT 8.555 185.090 8.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 184.685 8.875 185.005 ;
      LAYER met4 ;
        RECT 8.555 184.685 8.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 184.280 8.875 184.600 ;
      LAYER met4 ;
        RECT 8.555 184.280 8.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 183.875 8.875 184.195 ;
      LAYER met4 ;
        RECT 8.555 183.875 8.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 183.470 8.875 183.790 ;
      LAYER met4 ;
        RECT 8.555 183.470 8.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 183.065 8.875 183.385 ;
      LAYER met4 ;
        RECT 8.555 183.065 8.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 182.660 8.875 182.980 ;
      LAYER met4 ;
        RECT 8.555 182.660 8.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 182.255 8.875 182.575 ;
      LAYER met4 ;
        RECT 8.555 182.255 8.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 181.850 8.875 182.170 ;
      LAYER met4 ;
        RECT 8.555 181.850 8.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.555 181.445 8.875 181.765 ;
      LAYER met4 ;
        RECT 8.555 181.445 8.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 28.210 8.515 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 27.780 8.515 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 27.350 8.515 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 26.920 8.515 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 26.490 8.515 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 26.060 8.515 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 25.630 8.515 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 25.200 8.515 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 24.770 8.515 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 24.340 8.515 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.315 23.910 8.515 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 197.645 8.475 197.965 ;
      LAYER met4 ;
        RECT 8.155 197.645 8.475 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 197.240 8.475 197.560 ;
      LAYER met4 ;
        RECT 8.155 197.240 8.475 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 196.835 8.475 197.155 ;
      LAYER met4 ;
        RECT 8.155 196.835 8.475 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 196.430 8.475 196.750 ;
      LAYER met4 ;
        RECT 8.155 196.430 8.475 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 196.025 8.475 196.345 ;
      LAYER met4 ;
        RECT 8.155 196.025 8.475 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 195.620 8.475 195.940 ;
      LAYER met4 ;
        RECT 8.155 195.620 8.475 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 195.215 8.475 195.535 ;
      LAYER met4 ;
        RECT 8.155 195.215 8.475 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 194.810 8.475 195.130 ;
      LAYER met4 ;
        RECT 8.155 194.810 8.475 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 194.405 8.475 194.725 ;
      LAYER met4 ;
        RECT 8.155 194.405 8.475 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 194.000 8.475 194.320 ;
      LAYER met4 ;
        RECT 8.155 194.000 8.475 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 193.595 8.475 193.915 ;
      LAYER met4 ;
        RECT 8.155 193.595 8.475 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 193.190 8.475 193.510 ;
      LAYER met4 ;
        RECT 8.155 193.190 8.475 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 192.785 8.475 193.105 ;
      LAYER met4 ;
        RECT 8.155 192.785 8.475 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 192.380 8.475 192.700 ;
      LAYER met4 ;
        RECT 8.155 192.380 8.475 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 191.975 8.475 192.295 ;
      LAYER met4 ;
        RECT 8.155 191.975 8.475 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 191.570 8.475 191.890 ;
      LAYER met4 ;
        RECT 8.155 191.570 8.475 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 191.165 8.475 191.485 ;
      LAYER met4 ;
        RECT 8.155 191.165 8.475 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 190.760 8.475 191.080 ;
      LAYER met4 ;
        RECT 8.155 190.760 8.475 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 190.355 8.475 190.675 ;
      LAYER met4 ;
        RECT 8.155 190.355 8.475 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 189.950 8.475 190.270 ;
      LAYER met4 ;
        RECT 8.155 189.950 8.475 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 189.545 8.475 189.865 ;
      LAYER met4 ;
        RECT 8.155 189.545 8.475 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 189.140 8.475 189.460 ;
      LAYER met4 ;
        RECT 8.155 189.140 8.475 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 188.735 8.475 189.055 ;
      LAYER met4 ;
        RECT 8.155 188.735 8.475 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 188.330 8.475 188.650 ;
      LAYER met4 ;
        RECT 8.155 188.330 8.475 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 187.925 8.475 188.245 ;
      LAYER met4 ;
        RECT 8.155 187.925 8.475 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 187.520 8.475 187.840 ;
      LAYER met4 ;
        RECT 8.155 187.520 8.475 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 187.115 8.475 187.435 ;
      LAYER met4 ;
        RECT 8.155 187.115 8.475 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 186.710 8.475 187.030 ;
      LAYER met4 ;
        RECT 8.155 186.710 8.475 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 186.305 8.475 186.625 ;
      LAYER met4 ;
        RECT 8.155 186.305 8.475 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 185.900 8.475 186.220 ;
      LAYER met4 ;
        RECT 8.155 185.900 8.475 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 185.495 8.475 185.815 ;
      LAYER met4 ;
        RECT 8.155 185.495 8.475 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 185.090 8.475 185.410 ;
      LAYER met4 ;
        RECT 8.155 185.090 8.475 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 184.685 8.475 185.005 ;
      LAYER met4 ;
        RECT 8.155 184.685 8.475 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 184.280 8.475 184.600 ;
      LAYER met4 ;
        RECT 8.155 184.280 8.475 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 183.875 8.475 184.195 ;
      LAYER met4 ;
        RECT 8.155 183.875 8.475 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 183.470 8.475 183.790 ;
      LAYER met4 ;
        RECT 8.155 183.470 8.475 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 183.065 8.475 183.385 ;
      LAYER met4 ;
        RECT 8.155 183.065 8.475 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 182.660 8.475 182.980 ;
      LAYER met4 ;
        RECT 8.155 182.660 8.475 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 182.255 8.475 182.575 ;
      LAYER met4 ;
        RECT 8.155 182.255 8.475 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 181.850 8.475 182.170 ;
      LAYER met4 ;
        RECT 8.155 181.850 8.475 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.155 181.445 8.475 181.765 ;
      LAYER met4 ;
        RECT 8.155 181.445 8.475 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 28.210 8.110 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 27.780 8.110 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 27.350 8.110 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 26.920 8.110 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 26.490 8.110 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 26.060 8.110 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 25.630 8.110 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 25.200 8.110 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 24.770 8.110 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 24.340 8.110 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.910 23.910 8.110 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 197.645 8.075 197.965 ;
      LAYER met4 ;
        RECT 7.755 197.645 8.075 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 197.240 8.075 197.560 ;
      LAYER met4 ;
        RECT 7.755 197.240 8.075 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 196.835 8.075 197.155 ;
      LAYER met4 ;
        RECT 7.755 196.835 8.075 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 196.430 8.075 196.750 ;
      LAYER met4 ;
        RECT 7.755 196.430 8.075 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 196.025 8.075 196.345 ;
      LAYER met4 ;
        RECT 7.755 196.025 8.075 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 195.620 8.075 195.940 ;
      LAYER met4 ;
        RECT 7.755 195.620 8.075 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 195.215 8.075 195.535 ;
      LAYER met4 ;
        RECT 7.755 195.215 8.075 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 194.810 8.075 195.130 ;
      LAYER met4 ;
        RECT 7.755 194.810 8.075 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 194.405 8.075 194.725 ;
      LAYER met4 ;
        RECT 7.755 194.405 8.075 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 194.000 8.075 194.320 ;
      LAYER met4 ;
        RECT 7.755 194.000 8.075 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 193.595 8.075 193.915 ;
      LAYER met4 ;
        RECT 7.755 193.595 8.075 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 193.190 8.075 193.510 ;
      LAYER met4 ;
        RECT 7.755 193.190 8.075 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 192.785 8.075 193.105 ;
      LAYER met4 ;
        RECT 7.755 192.785 8.075 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 192.380 8.075 192.700 ;
      LAYER met4 ;
        RECT 7.755 192.380 8.075 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 191.975 8.075 192.295 ;
      LAYER met4 ;
        RECT 7.755 191.975 8.075 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 191.570 8.075 191.890 ;
      LAYER met4 ;
        RECT 7.755 191.570 8.075 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 191.165 8.075 191.485 ;
      LAYER met4 ;
        RECT 7.755 191.165 8.075 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 190.760 8.075 191.080 ;
      LAYER met4 ;
        RECT 7.755 190.760 8.075 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 190.355 8.075 190.675 ;
      LAYER met4 ;
        RECT 7.755 190.355 8.075 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 189.950 8.075 190.270 ;
      LAYER met4 ;
        RECT 7.755 189.950 8.075 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 189.545 8.075 189.865 ;
      LAYER met4 ;
        RECT 7.755 189.545 8.075 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 189.140 8.075 189.460 ;
      LAYER met4 ;
        RECT 7.755 189.140 8.075 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 188.735 8.075 189.055 ;
      LAYER met4 ;
        RECT 7.755 188.735 8.075 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 188.330 8.075 188.650 ;
      LAYER met4 ;
        RECT 7.755 188.330 8.075 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 187.925 8.075 188.245 ;
      LAYER met4 ;
        RECT 7.755 187.925 8.075 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 187.520 8.075 187.840 ;
      LAYER met4 ;
        RECT 7.755 187.520 8.075 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 187.115 8.075 187.435 ;
      LAYER met4 ;
        RECT 7.755 187.115 8.075 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 186.710 8.075 187.030 ;
      LAYER met4 ;
        RECT 7.755 186.710 8.075 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 186.305 8.075 186.625 ;
      LAYER met4 ;
        RECT 7.755 186.305 8.075 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 185.900 8.075 186.220 ;
      LAYER met4 ;
        RECT 7.755 185.900 8.075 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 185.495 8.075 185.815 ;
      LAYER met4 ;
        RECT 7.755 185.495 8.075 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 185.090 8.075 185.410 ;
      LAYER met4 ;
        RECT 7.755 185.090 8.075 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 184.685 8.075 185.005 ;
      LAYER met4 ;
        RECT 7.755 184.685 8.075 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 184.280 8.075 184.600 ;
      LAYER met4 ;
        RECT 7.755 184.280 8.075 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 183.875 8.075 184.195 ;
      LAYER met4 ;
        RECT 7.755 183.875 8.075 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 183.470 8.075 183.790 ;
      LAYER met4 ;
        RECT 7.755 183.470 8.075 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 183.065 8.075 183.385 ;
      LAYER met4 ;
        RECT 7.755 183.065 8.075 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 182.660 8.075 182.980 ;
      LAYER met4 ;
        RECT 7.755 182.660 8.075 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 182.255 8.075 182.575 ;
      LAYER met4 ;
        RECT 7.755 182.255 8.075 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 181.850 8.075 182.170 ;
      LAYER met4 ;
        RECT 7.755 181.850 8.075 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.755 181.445 8.075 181.765 ;
      LAYER met4 ;
        RECT 7.755 181.445 8.075 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 28.210 7.705 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 27.780 7.705 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 27.350 7.705 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 26.920 7.705 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 26.490 7.705 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 26.060 7.705 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 25.630 7.705 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 25.200 7.705 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 24.770 7.705 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 24.340 7.705 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.505 23.910 7.705 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 197.645 7.675 197.965 ;
      LAYER met4 ;
        RECT 7.355 197.645 7.675 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 197.240 7.675 197.560 ;
      LAYER met4 ;
        RECT 7.355 197.240 7.675 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 196.835 7.675 197.155 ;
      LAYER met4 ;
        RECT 7.355 196.835 7.675 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 196.430 7.675 196.750 ;
      LAYER met4 ;
        RECT 7.355 196.430 7.675 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 196.025 7.675 196.345 ;
      LAYER met4 ;
        RECT 7.355 196.025 7.675 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 195.620 7.675 195.940 ;
      LAYER met4 ;
        RECT 7.355 195.620 7.675 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 195.215 7.675 195.535 ;
      LAYER met4 ;
        RECT 7.355 195.215 7.675 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 194.810 7.675 195.130 ;
      LAYER met4 ;
        RECT 7.355 194.810 7.675 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 194.405 7.675 194.725 ;
      LAYER met4 ;
        RECT 7.355 194.405 7.675 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 194.000 7.675 194.320 ;
      LAYER met4 ;
        RECT 7.355 194.000 7.675 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 193.595 7.675 193.915 ;
      LAYER met4 ;
        RECT 7.355 193.595 7.675 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 193.190 7.675 193.510 ;
      LAYER met4 ;
        RECT 7.355 193.190 7.675 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 192.785 7.675 193.105 ;
      LAYER met4 ;
        RECT 7.355 192.785 7.675 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 192.380 7.675 192.700 ;
      LAYER met4 ;
        RECT 7.355 192.380 7.675 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 191.975 7.675 192.295 ;
      LAYER met4 ;
        RECT 7.355 191.975 7.675 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 191.570 7.675 191.890 ;
      LAYER met4 ;
        RECT 7.355 191.570 7.675 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 191.165 7.675 191.485 ;
      LAYER met4 ;
        RECT 7.355 191.165 7.675 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 190.760 7.675 191.080 ;
      LAYER met4 ;
        RECT 7.355 190.760 7.675 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 190.355 7.675 190.675 ;
      LAYER met4 ;
        RECT 7.355 190.355 7.675 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 189.950 7.675 190.270 ;
      LAYER met4 ;
        RECT 7.355 189.950 7.675 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 189.545 7.675 189.865 ;
      LAYER met4 ;
        RECT 7.355 189.545 7.675 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 189.140 7.675 189.460 ;
      LAYER met4 ;
        RECT 7.355 189.140 7.675 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 188.735 7.675 189.055 ;
      LAYER met4 ;
        RECT 7.355 188.735 7.675 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 188.330 7.675 188.650 ;
      LAYER met4 ;
        RECT 7.355 188.330 7.675 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 187.925 7.675 188.245 ;
      LAYER met4 ;
        RECT 7.355 187.925 7.675 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 187.520 7.675 187.840 ;
      LAYER met4 ;
        RECT 7.355 187.520 7.675 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 187.115 7.675 187.435 ;
      LAYER met4 ;
        RECT 7.355 187.115 7.675 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 186.710 7.675 187.030 ;
      LAYER met4 ;
        RECT 7.355 186.710 7.675 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 186.305 7.675 186.625 ;
      LAYER met4 ;
        RECT 7.355 186.305 7.675 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 185.900 7.675 186.220 ;
      LAYER met4 ;
        RECT 7.355 185.900 7.675 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 185.495 7.675 185.815 ;
      LAYER met4 ;
        RECT 7.355 185.495 7.675 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 185.090 7.675 185.410 ;
      LAYER met4 ;
        RECT 7.355 185.090 7.675 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 184.685 7.675 185.005 ;
      LAYER met4 ;
        RECT 7.355 184.685 7.675 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 184.280 7.675 184.600 ;
      LAYER met4 ;
        RECT 7.355 184.280 7.675 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 183.875 7.675 184.195 ;
      LAYER met4 ;
        RECT 7.355 183.875 7.675 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 183.470 7.675 183.790 ;
      LAYER met4 ;
        RECT 7.355 183.470 7.675 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 183.065 7.675 183.385 ;
      LAYER met4 ;
        RECT 7.355 183.065 7.675 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 182.660 7.675 182.980 ;
      LAYER met4 ;
        RECT 7.355 182.660 7.675 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 182.255 7.675 182.575 ;
      LAYER met4 ;
        RECT 7.355 182.255 7.675 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 181.850 7.675 182.170 ;
      LAYER met4 ;
        RECT 7.355 181.850 7.675 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.355 181.445 7.675 181.765 ;
      LAYER met4 ;
        RECT 7.355 181.445 7.675 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 28.210 7.300 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 27.780 7.300 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 27.350 7.300 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 26.920 7.300 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 26.490 7.300 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 26.060 7.300 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 25.630 7.300 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 25.200 7.300 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 24.770 7.300 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 24.340 7.300 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 23.910 7.300 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 197.645 7.275 197.965 ;
      LAYER met4 ;
        RECT 6.955 197.645 7.275 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 197.240 7.275 197.560 ;
      LAYER met4 ;
        RECT 6.955 197.240 7.275 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 196.835 7.275 197.155 ;
      LAYER met4 ;
        RECT 6.955 196.835 7.275 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 196.430 7.275 196.750 ;
      LAYER met4 ;
        RECT 6.955 196.430 7.275 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 196.025 7.275 196.345 ;
      LAYER met4 ;
        RECT 6.955 196.025 7.275 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 195.620 7.275 195.940 ;
      LAYER met4 ;
        RECT 6.955 195.620 7.275 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 195.215 7.275 195.535 ;
      LAYER met4 ;
        RECT 6.955 195.215 7.275 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 194.810 7.275 195.130 ;
      LAYER met4 ;
        RECT 6.955 194.810 7.275 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 194.405 7.275 194.725 ;
      LAYER met4 ;
        RECT 6.955 194.405 7.275 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 194.000 7.275 194.320 ;
      LAYER met4 ;
        RECT 6.955 194.000 7.275 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 193.595 7.275 193.915 ;
      LAYER met4 ;
        RECT 6.955 193.595 7.275 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 193.190 7.275 193.510 ;
      LAYER met4 ;
        RECT 6.955 193.190 7.275 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 192.785 7.275 193.105 ;
      LAYER met4 ;
        RECT 6.955 192.785 7.275 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 192.380 7.275 192.700 ;
      LAYER met4 ;
        RECT 6.955 192.380 7.275 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 191.975 7.275 192.295 ;
      LAYER met4 ;
        RECT 6.955 191.975 7.275 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 191.570 7.275 191.890 ;
      LAYER met4 ;
        RECT 6.955 191.570 7.275 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 191.165 7.275 191.485 ;
      LAYER met4 ;
        RECT 6.955 191.165 7.275 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 190.760 7.275 191.080 ;
      LAYER met4 ;
        RECT 6.955 190.760 7.275 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 190.355 7.275 190.675 ;
      LAYER met4 ;
        RECT 6.955 190.355 7.275 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 189.950 7.275 190.270 ;
      LAYER met4 ;
        RECT 6.955 189.950 7.275 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 189.545 7.275 189.865 ;
      LAYER met4 ;
        RECT 6.955 189.545 7.275 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 189.140 7.275 189.460 ;
      LAYER met4 ;
        RECT 6.955 189.140 7.275 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 188.735 7.275 189.055 ;
      LAYER met4 ;
        RECT 6.955 188.735 7.275 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 188.330 7.275 188.650 ;
      LAYER met4 ;
        RECT 6.955 188.330 7.275 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 187.925 7.275 188.245 ;
      LAYER met4 ;
        RECT 6.955 187.925 7.275 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 187.520 7.275 187.840 ;
      LAYER met4 ;
        RECT 6.955 187.520 7.275 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 187.115 7.275 187.435 ;
      LAYER met4 ;
        RECT 6.955 187.115 7.275 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 186.710 7.275 187.030 ;
      LAYER met4 ;
        RECT 6.955 186.710 7.275 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 186.305 7.275 186.625 ;
      LAYER met4 ;
        RECT 6.955 186.305 7.275 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 185.900 7.275 186.220 ;
      LAYER met4 ;
        RECT 6.955 185.900 7.275 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 185.495 7.275 185.815 ;
      LAYER met4 ;
        RECT 6.955 185.495 7.275 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 185.090 7.275 185.410 ;
      LAYER met4 ;
        RECT 6.955 185.090 7.275 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 184.685 7.275 185.005 ;
      LAYER met4 ;
        RECT 6.955 184.685 7.275 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 184.280 7.275 184.600 ;
      LAYER met4 ;
        RECT 6.955 184.280 7.275 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 183.875 7.275 184.195 ;
      LAYER met4 ;
        RECT 6.955 183.875 7.275 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 183.470 7.275 183.790 ;
      LAYER met4 ;
        RECT 6.955 183.470 7.275 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 183.065 7.275 183.385 ;
      LAYER met4 ;
        RECT 6.955 183.065 7.275 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 182.660 7.275 182.980 ;
      LAYER met4 ;
        RECT 6.955 182.660 7.275 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 182.255 7.275 182.575 ;
      LAYER met4 ;
        RECT 6.955 182.255 7.275 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 181.850 7.275 182.170 ;
      LAYER met4 ;
        RECT 6.955 181.850 7.275 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.955 181.445 7.275 181.765 ;
      LAYER met4 ;
        RECT 6.955 181.445 7.275 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 28.210 6.895 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 27.780 6.895 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 27.350 6.895 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 26.920 6.895 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 26.490 6.895 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 26.060 6.895 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 25.630 6.895 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 25.200 6.895 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 24.770 6.895 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 24.340 6.895 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.695 23.910 6.895 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 197.645 6.875 197.965 ;
      LAYER met4 ;
        RECT 6.555 197.645 6.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 197.240 6.875 197.560 ;
      LAYER met4 ;
        RECT 6.555 197.240 6.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 196.835 6.875 197.155 ;
      LAYER met4 ;
        RECT 6.555 196.835 6.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 196.430 6.875 196.750 ;
      LAYER met4 ;
        RECT 6.555 196.430 6.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 196.025 6.875 196.345 ;
      LAYER met4 ;
        RECT 6.555 196.025 6.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 195.620 6.875 195.940 ;
      LAYER met4 ;
        RECT 6.555 195.620 6.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 195.215 6.875 195.535 ;
      LAYER met4 ;
        RECT 6.555 195.215 6.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 194.810 6.875 195.130 ;
      LAYER met4 ;
        RECT 6.555 194.810 6.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 194.405 6.875 194.725 ;
      LAYER met4 ;
        RECT 6.555 194.405 6.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 194.000 6.875 194.320 ;
      LAYER met4 ;
        RECT 6.555 194.000 6.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 193.595 6.875 193.915 ;
      LAYER met4 ;
        RECT 6.555 193.595 6.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 193.190 6.875 193.510 ;
      LAYER met4 ;
        RECT 6.555 193.190 6.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 192.785 6.875 193.105 ;
      LAYER met4 ;
        RECT 6.555 192.785 6.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 192.380 6.875 192.700 ;
      LAYER met4 ;
        RECT 6.555 192.380 6.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 191.975 6.875 192.295 ;
      LAYER met4 ;
        RECT 6.555 191.975 6.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 191.570 6.875 191.890 ;
      LAYER met4 ;
        RECT 6.555 191.570 6.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 191.165 6.875 191.485 ;
      LAYER met4 ;
        RECT 6.555 191.165 6.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 190.760 6.875 191.080 ;
      LAYER met4 ;
        RECT 6.555 190.760 6.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 190.355 6.875 190.675 ;
      LAYER met4 ;
        RECT 6.555 190.355 6.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 189.950 6.875 190.270 ;
      LAYER met4 ;
        RECT 6.555 189.950 6.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 189.545 6.875 189.865 ;
      LAYER met4 ;
        RECT 6.555 189.545 6.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 189.140 6.875 189.460 ;
      LAYER met4 ;
        RECT 6.555 189.140 6.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 188.735 6.875 189.055 ;
      LAYER met4 ;
        RECT 6.555 188.735 6.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 188.330 6.875 188.650 ;
      LAYER met4 ;
        RECT 6.555 188.330 6.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 187.925 6.875 188.245 ;
      LAYER met4 ;
        RECT 6.555 187.925 6.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 187.520 6.875 187.840 ;
      LAYER met4 ;
        RECT 6.555 187.520 6.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 187.115 6.875 187.435 ;
      LAYER met4 ;
        RECT 6.555 187.115 6.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 186.710 6.875 187.030 ;
      LAYER met4 ;
        RECT 6.555 186.710 6.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 186.305 6.875 186.625 ;
      LAYER met4 ;
        RECT 6.555 186.305 6.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 185.900 6.875 186.220 ;
      LAYER met4 ;
        RECT 6.555 185.900 6.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 185.495 6.875 185.815 ;
      LAYER met4 ;
        RECT 6.555 185.495 6.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 185.090 6.875 185.410 ;
      LAYER met4 ;
        RECT 6.555 185.090 6.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 184.685 6.875 185.005 ;
      LAYER met4 ;
        RECT 6.555 184.685 6.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 184.280 6.875 184.600 ;
      LAYER met4 ;
        RECT 6.555 184.280 6.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 183.875 6.875 184.195 ;
      LAYER met4 ;
        RECT 6.555 183.875 6.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 183.470 6.875 183.790 ;
      LAYER met4 ;
        RECT 6.555 183.470 6.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 183.065 6.875 183.385 ;
      LAYER met4 ;
        RECT 6.555 183.065 6.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 182.660 6.875 182.980 ;
      LAYER met4 ;
        RECT 6.555 182.660 6.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 182.255 6.875 182.575 ;
      LAYER met4 ;
        RECT 6.555 182.255 6.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 181.850 6.875 182.170 ;
      LAYER met4 ;
        RECT 6.555 181.850 6.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.555 181.445 6.875 181.765 ;
      LAYER met4 ;
        RECT 6.555 181.445 6.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 28.210 6.490 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 27.780 6.490 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 27.350 6.490 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 26.920 6.490 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 26.490 6.490 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 26.060 6.490 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 25.630 6.490 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 25.200 6.490 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 24.770 6.490 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 24.340 6.490 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.290 23.910 6.490 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 197.645 6.475 197.965 ;
      LAYER met4 ;
        RECT 6.155 197.645 6.475 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 197.240 6.475 197.560 ;
      LAYER met4 ;
        RECT 6.155 197.240 6.475 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 196.835 6.475 197.155 ;
      LAYER met4 ;
        RECT 6.155 196.835 6.475 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 196.430 6.475 196.750 ;
      LAYER met4 ;
        RECT 6.155 196.430 6.475 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 196.025 6.475 196.345 ;
      LAYER met4 ;
        RECT 6.155 196.025 6.475 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 195.620 6.475 195.940 ;
      LAYER met4 ;
        RECT 6.155 195.620 6.475 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 195.215 6.475 195.535 ;
      LAYER met4 ;
        RECT 6.155 195.215 6.475 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 194.810 6.475 195.130 ;
      LAYER met4 ;
        RECT 6.155 194.810 6.475 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 194.405 6.475 194.725 ;
      LAYER met4 ;
        RECT 6.155 194.405 6.475 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 194.000 6.475 194.320 ;
      LAYER met4 ;
        RECT 6.155 194.000 6.475 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 193.595 6.475 193.915 ;
      LAYER met4 ;
        RECT 6.155 193.595 6.475 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 193.190 6.475 193.510 ;
      LAYER met4 ;
        RECT 6.155 193.190 6.475 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 192.785 6.475 193.105 ;
      LAYER met4 ;
        RECT 6.155 192.785 6.475 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 192.380 6.475 192.700 ;
      LAYER met4 ;
        RECT 6.155 192.380 6.475 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 191.975 6.475 192.295 ;
      LAYER met4 ;
        RECT 6.155 191.975 6.475 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 191.570 6.475 191.890 ;
      LAYER met4 ;
        RECT 6.155 191.570 6.475 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 191.165 6.475 191.485 ;
      LAYER met4 ;
        RECT 6.155 191.165 6.475 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 190.760 6.475 191.080 ;
      LAYER met4 ;
        RECT 6.155 190.760 6.475 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 190.355 6.475 190.675 ;
      LAYER met4 ;
        RECT 6.155 190.355 6.475 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 189.950 6.475 190.270 ;
      LAYER met4 ;
        RECT 6.155 189.950 6.475 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 189.545 6.475 189.865 ;
      LAYER met4 ;
        RECT 6.155 189.545 6.475 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 189.140 6.475 189.460 ;
      LAYER met4 ;
        RECT 6.155 189.140 6.475 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 188.735 6.475 189.055 ;
      LAYER met4 ;
        RECT 6.155 188.735 6.475 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 188.330 6.475 188.650 ;
      LAYER met4 ;
        RECT 6.155 188.330 6.475 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 187.925 6.475 188.245 ;
      LAYER met4 ;
        RECT 6.155 187.925 6.475 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 187.520 6.475 187.840 ;
      LAYER met4 ;
        RECT 6.155 187.520 6.475 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 187.115 6.475 187.435 ;
      LAYER met4 ;
        RECT 6.155 187.115 6.475 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 186.710 6.475 187.030 ;
      LAYER met4 ;
        RECT 6.155 186.710 6.475 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 186.305 6.475 186.625 ;
      LAYER met4 ;
        RECT 6.155 186.305 6.475 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 185.900 6.475 186.220 ;
      LAYER met4 ;
        RECT 6.155 185.900 6.475 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 185.495 6.475 185.815 ;
      LAYER met4 ;
        RECT 6.155 185.495 6.475 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 185.090 6.475 185.410 ;
      LAYER met4 ;
        RECT 6.155 185.090 6.475 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 184.685 6.475 185.005 ;
      LAYER met4 ;
        RECT 6.155 184.685 6.475 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 184.280 6.475 184.600 ;
      LAYER met4 ;
        RECT 6.155 184.280 6.475 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 183.875 6.475 184.195 ;
      LAYER met4 ;
        RECT 6.155 183.875 6.475 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 183.470 6.475 183.790 ;
      LAYER met4 ;
        RECT 6.155 183.470 6.475 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 183.065 6.475 183.385 ;
      LAYER met4 ;
        RECT 6.155 183.065 6.475 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 182.660 6.475 182.980 ;
      LAYER met4 ;
        RECT 6.155 182.660 6.475 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 182.255 6.475 182.575 ;
      LAYER met4 ;
        RECT 6.155 182.255 6.475 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 181.850 6.475 182.170 ;
      LAYER met4 ;
        RECT 6.155 181.850 6.475 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.155 181.445 6.475 181.765 ;
      LAYER met4 ;
        RECT 6.155 181.445 6.475 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 28.210 6.085 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 27.780 6.085 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 27.350 6.085 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 26.920 6.085 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 26.490 6.085 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 26.060 6.085 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 25.630 6.085 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 25.200 6.085 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 24.770 6.085 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 24.340 6.085 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.885 23.910 6.085 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 197.645 6.075 197.965 ;
      LAYER met4 ;
        RECT 5.755 197.645 6.075 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 197.240 6.075 197.560 ;
      LAYER met4 ;
        RECT 5.755 197.240 6.075 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 196.835 6.075 197.155 ;
      LAYER met4 ;
        RECT 5.755 196.835 6.075 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 196.430 6.075 196.750 ;
      LAYER met4 ;
        RECT 5.755 196.430 6.075 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 196.025 6.075 196.345 ;
      LAYER met4 ;
        RECT 5.755 196.025 6.075 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 195.620 6.075 195.940 ;
      LAYER met4 ;
        RECT 5.755 195.620 6.075 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 195.215 6.075 195.535 ;
      LAYER met4 ;
        RECT 5.755 195.215 6.075 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 194.810 6.075 195.130 ;
      LAYER met4 ;
        RECT 5.755 194.810 6.075 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 194.405 6.075 194.725 ;
      LAYER met4 ;
        RECT 5.755 194.405 6.075 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 194.000 6.075 194.320 ;
      LAYER met4 ;
        RECT 5.755 194.000 6.075 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 193.595 6.075 193.915 ;
      LAYER met4 ;
        RECT 5.755 193.595 6.075 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 193.190 6.075 193.510 ;
      LAYER met4 ;
        RECT 5.755 193.190 6.075 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 192.785 6.075 193.105 ;
      LAYER met4 ;
        RECT 5.755 192.785 6.075 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 192.380 6.075 192.700 ;
      LAYER met4 ;
        RECT 5.755 192.380 6.075 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 191.975 6.075 192.295 ;
      LAYER met4 ;
        RECT 5.755 191.975 6.075 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 191.570 6.075 191.890 ;
      LAYER met4 ;
        RECT 5.755 191.570 6.075 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 191.165 6.075 191.485 ;
      LAYER met4 ;
        RECT 5.755 191.165 6.075 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 190.760 6.075 191.080 ;
      LAYER met4 ;
        RECT 5.755 190.760 6.075 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 190.355 6.075 190.675 ;
      LAYER met4 ;
        RECT 5.755 190.355 6.075 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 189.950 6.075 190.270 ;
      LAYER met4 ;
        RECT 5.755 189.950 6.075 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 189.545 6.075 189.865 ;
      LAYER met4 ;
        RECT 5.755 189.545 6.075 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 189.140 6.075 189.460 ;
      LAYER met4 ;
        RECT 5.755 189.140 6.075 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 188.735 6.075 189.055 ;
      LAYER met4 ;
        RECT 5.755 188.735 6.075 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 188.330 6.075 188.650 ;
      LAYER met4 ;
        RECT 5.755 188.330 6.075 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 187.925 6.075 188.245 ;
      LAYER met4 ;
        RECT 5.755 187.925 6.075 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 187.520 6.075 187.840 ;
      LAYER met4 ;
        RECT 5.755 187.520 6.075 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 187.115 6.075 187.435 ;
      LAYER met4 ;
        RECT 5.755 187.115 6.075 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 186.710 6.075 187.030 ;
      LAYER met4 ;
        RECT 5.755 186.710 6.075 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 186.305 6.075 186.625 ;
      LAYER met4 ;
        RECT 5.755 186.305 6.075 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 185.900 6.075 186.220 ;
      LAYER met4 ;
        RECT 5.755 185.900 6.075 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 185.495 6.075 185.815 ;
      LAYER met4 ;
        RECT 5.755 185.495 6.075 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 185.090 6.075 185.410 ;
      LAYER met4 ;
        RECT 5.755 185.090 6.075 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 184.685 6.075 185.005 ;
      LAYER met4 ;
        RECT 5.755 184.685 6.075 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 184.280 6.075 184.600 ;
      LAYER met4 ;
        RECT 5.755 184.280 6.075 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 183.875 6.075 184.195 ;
      LAYER met4 ;
        RECT 5.755 183.875 6.075 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 183.470 6.075 183.790 ;
      LAYER met4 ;
        RECT 5.755 183.470 6.075 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 183.065 6.075 183.385 ;
      LAYER met4 ;
        RECT 5.755 183.065 6.075 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 182.660 6.075 182.980 ;
      LAYER met4 ;
        RECT 5.755 182.660 6.075 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 182.255 6.075 182.575 ;
      LAYER met4 ;
        RECT 5.755 182.255 6.075 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 181.850 6.075 182.170 ;
      LAYER met4 ;
        RECT 5.755 181.850 6.075 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.755 181.445 6.075 181.765 ;
      LAYER met4 ;
        RECT 5.755 181.445 6.075 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 28.210 5.680 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 27.780 5.680 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 27.350 5.680 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 26.920 5.680 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 26.490 5.680 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 26.060 5.680 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 25.630 5.680 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 25.200 5.680 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 24.770 5.680 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 24.340 5.680 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.480 23.910 5.680 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 197.645 5.675 197.965 ;
      LAYER met4 ;
        RECT 5.355 197.645 5.675 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 197.240 5.675 197.560 ;
      LAYER met4 ;
        RECT 5.355 197.240 5.675 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 196.835 5.675 197.155 ;
      LAYER met4 ;
        RECT 5.355 196.835 5.675 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 196.430 5.675 196.750 ;
      LAYER met4 ;
        RECT 5.355 196.430 5.675 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 196.025 5.675 196.345 ;
      LAYER met4 ;
        RECT 5.355 196.025 5.675 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 195.620 5.675 195.940 ;
      LAYER met4 ;
        RECT 5.355 195.620 5.675 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 195.215 5.675 195.535 ;
      LAYER met4 ;
        RECT 5.355 195.215 5.675 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 194.810 5.675 195.130 ;
      LAYER met4 ;
        RECT 5.355 194.810 5.675 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 194.405 5.675 194.725 ;
      LAYER met4 ;
        RECT 5.355 194.405 5.675 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 194.000 5.675 194.320 ;
      LAYER met4 ;
        RECT 5.355 194.000 5.675 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 193.595 5.675 193.915 ;
      LAYER met4 ;
        RECT 5.355 193.595 5.675 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 193.190 5.675 193.510 ;
      LAYER met4 ;
        RECT 5.355 193.190 5.675 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 192.785 5.675 193.105 ;
      LAYER met4 ;
        RECT 5.355 192.785 5.675 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 192.380 5.675 192.700 ;
      LAYER met4 ;
        RECT 5.355 192.380 5.675 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 191.975 5.675 192.295 ;
      LAYER met4 ;
        RECT 5.355 191.975 5.675 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 191.570 5.675 191.890 ;
      LAYER met4 ;
        RECT 5.355 191.570 5.675 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 191.165 5.675 191.485 ;
      LAYER met4 ;
        RECT 5.355 191.165 5.675 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 190.760 5.675 191.080 ;
      LAYER met4 ;
        RECT 5.355 190.760 5.675 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 190.355 5.675 190.675 ;
      LAYER met4 ;
        RECT 5.355 190.355 5.675 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 189.950 5.675 190.270 ;
      LAYER met4 ;
        RECT 5.355 189.950 5.675 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 189.545 5.675 189.865 ;
      LAYER met4 ;
        RECT 5.355 189.545 5.675 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 189.140 5.675 189.460 ;
      LAYER met4 ;
        RECT 5.355 189.140 5.675 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 188.735 5.675 189.055 ;
      LAYER met4 ;
        RECT 5.355 188.735 5.675 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 188.330 5.675 188.650 ;
      LAYER met4 ;
        RECT 5.355 188.330 5.675 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 187.925 5.675 188.245 ;
      LAYER met4 ;
        RECT 5.355 187.925 5.675 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 187.520 5.675 187.840 ;
      LAYER met4 ;
        RECT 5.355 187.520 5.675 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 187.115 5.675 187.435 ;
      LAYER met4 ;
        RECT 5.355 187.115 5.675 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 186.710 5.675 187.030 ;
      LAYER met4 ;
        RECT 5.355 186.710 5.675 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 186.305 5.675 186.625 ;
      LAYER met4 ;
        RECT 5.355 186.305 5.675 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 185.900 5.675 186.220 ;
      LAYER met4 ;
        RECT 5.355 185.900 5.675 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 185.495 5.675 185.815 ;
      LAYER met4 ;
        RECT 5.355 185.495 5.675 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 185.090 5.675 185.410 ;
      LAYER met4 ;
        RECT 5.355 185.090 5.675 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 184.685 5.675 185.005 ;
      LAYER met4 ;
        RECT 5.355 184.685 5.675 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 184.280 5.675 184.600 ;
      LAYER met4 ;
        RECT 5.355 184.280 5.675 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 183.875 5.675 184.195 ;
      LAYER met4 ;
        RECT 5.355 183.875 5.675 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 183.470 5.675 183.790 ;
      LAYER met4 ;
        RECT 5.355 183.470 5.675 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 183.065 5.675 183.385 ;
      LAYER met4 ;
        RECT 5.355 183.065 5.675 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 182.660 5.675 182.980 ;
      LAYER met4 ;
        RECT 5.355 182.660 5.675 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 182.255 5.675 182.575 ;
      LAYER met4 ;
        RECT 5.355 182.255 5.675 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 181.850 5.675 182.170 ;
      LAYER met4 ;
        RECT 5.355 181.850 5.675 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.355 181.445 5.675 181.765 ;
      LAYER met4 ;
        RECT 5.355 181.445 5.675 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 28.210 5.275 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 27.780 5.275 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 27.350 5.275 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 26.920 5.275 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 26.490 5.275 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 26.060 5.275 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 25.630 5.275 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 25.200 5.275 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 24.770 5.275 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 24.340 5.275 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.075 23.910 5.275 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 197.645 5.275 197.965 ;
      LAYER met4 ;
        RECT 4.955 197.645 5.275 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 197.240 5.275 197.560 ;
      LAYER met4 ;
        RECT 4.955 197.240 5.275 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 196.835 5.275 197.155 ;
      LAYER met4 ;
        RECT 4.955 196.835 5.275 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 196.430 5.275 196.750 ;
      LAYER met4 ;
        RECT 4.955 196.430 5.275 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 196.025 5.275 196.345 ;
      LAYER met4 ;
        RECT 4.955 196.025 5.275 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 195.620 5.275 195.940 ;
      LAYER met4 ;
        RECT 4.955 195.620 5.275 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 195.215 5.275 195.535 ;
      LAYER met4 ;
        RECT 4.955 195.215 5.275 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 194.810 5.275 195.130 ;
      LAYER met4 ;
        RECT 4.955 194.810 5.275 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 194.405 5.275 194.725 ;
      LAYER met4 ;
        RECT 4.955 194.405 5.275 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 194.000 5.275 194.320 ;
      LAYER met4 ;
        RECT 4.955 194.000 5.275 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 193.595 5.275 193.915 ;
      LAYER met4 ;
        RECT 4.955 193.595 5.275 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 193.190 5.275 193.510 ;
      LAYER met4 ;
        RECT 4.955 193.190 5.275 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 192.785 5.275 193.105 ;
      LAYER met4 ;
        RECT 4.955 192.785 5.275 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 192.380 5.275 192.700 ;
      LAYER met4 ;
        RECT 4.955 192.380 5.275 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 191.975 5.275 192.295 ;
      LAYER met4 ;
        RECT 4.955 191.975 5.275 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 191.570 5.275 191.890 ;
      LAYER met4 ;
        RECT 4.955 191.570 5.275 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 191.165 5.275 191.485 ;
      LAYER met4 ;
        RECT 4.955 191.165 5.275 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 190.760 5.275 191.080 ;
      LAYER met4 ;
        RECT 4.955 190.760 5.275 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 190.355 5.275 190.675 ;
      LAYER met4 ;
        RECT 4.955 190.355 5.275 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 189.950 5.275 190.270 ;
      LAYER met4 ;
        RECT 4.955 189.950 5.275 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 189.545 5.275 189.865 ;
      LAYER met4 ;
        RECT 4.955 189.545 5.275 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 189.140 5.275 189.460 ;
      LAYER met4 ;
        RECT 4.955 189.140 5.275 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 188.735 5.275 189.055 ;
      LAYER met4 ;
        RECT 4.955 188.735 5.275 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 188.330 5.275 188.650 ;
      LAYER met4 ;
        RECT 4.955 188.330 5.275 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 187.925 5.275 188.245 ;
      LAYER met4 ;
        RECT 4.955 187.925 5.275 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 187.520 5.275 187.840 ;
      LAYER met4 ;
        RECT 4.955 187.520 5.275 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 187.115 5.275 187.435 ;
      LAYER met4 ;
        RECT 4.955 187.115 5.275 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 186.710 5.275 187.030 ;
      LAYER met4 ;
        RECT 4.955 186.710 5.275 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 186.305 5.275 186.625 ;
      LAYER met4 ;
        RECT 4.955 186.305 5.275 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 185.900 5.275 186.220 ;
      LAYER met4 ;
        RECT 4.955 185.900 5.275 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 185.495 5.275 185.815 ;
      LAYER met4 ;
        RECT 4.955 185.495 5.275 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 185.090 5.275 185.410 ;
      LAYER met4 ;
        RECT 4.955 185.090 5.275 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 184.685 5.275 185.005 ;
      LAYER met4 ;
        RECT 4.955 184.685 5.275 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 184.280 5.275 184.600 ;
      LAYER met4 ;
        RECT 4.955 184.280 5.275 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 183.875 5.275 184.195 ;
      LAYER met4 ;
        RECT 4.955 183.875 5.275 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 183.470 5.275 183.790 ;
      LAYER met4 ;
        RECT 4.955 183.470 5.275 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 183.065 5.275 183.385 ;
      LAYER met4 ;
        RECT 4.955 183.065 5.275 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 182.660 5.275 182.980 ;
      LAYER met4 ;
        RECT 4.955 182.660 5.275 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 182.255 5.275 182.575 ;
      LAYER met4 ;
        RECT 4.955 182.255 5.275 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 181.850 5.275 182.170 ;
      LAYER met4 ;
        RECT 4.955 181.850 5.275 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.955 181.445 5.275 181.765 ;
      LAYER met4 ;
        RECT 4.955 181.445 5.275 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 28.210 4.870 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 27.780 4.870 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 27.350 4.870 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 26.920 4.870 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 26.490 4.870 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 26.060 4.870 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 25.630 4.870 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 25.200 4.870 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 24.770 4.870 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 24.340 4.870 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.670 23.910 4.870 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 197.645 4.875 197.965 ;
      LAYER met4 ;
        RECT 4.555 197.645 4.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 197.240 4.875 197.560 ;
      LAYER met4 ;
        RECT 4.555 197.240 4.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 196.835 4.875 197.155 ;
      LAYER met4 ;
        RECT 4.555 196.835 4.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 196.430 4.875 196.750 ;
      LAYER met4 ;
        RECT 4.555 196.430 4.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 196.025 4.875 196.345 ;
      LAYER met4 ;
        RECT 4.555 196.025 4.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 195.620 4.875 195.940 ;
      LAYER met4 ;
        RECT 4.555 195.620 4.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 195.215 4.875 195.535 ;
      LAYER met4 ;
        RECT 4.555 195.215 4.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 194.810 4.875 195.130 ;
      LAYER met4 ;
        RECT 4.555 194.810 4.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 194.405 4.875 194.725 ;
      LAYER met4 ;
        RECT 4.555 194.405 4.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 194.000 4.875 194.320 ;
      LAYER met4 ;
        RECT 4.555 194.000 4.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 193.595 4.875 193.915 ;
      LAYER met4 ;
        RECT 4.555 193.595 4.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 193.190 4.875 193.510 ;
      LAYER met4 ;
        RECT 4.555 193.190 4.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 192.785 4.875 193.105 ;
      LAYER met4 ;
        RECT 4.555 192.785 4.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 192.380 4.875 192.700 ;
      LAYER met4 ;
        RECT 4.555 192.380 4.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 191.975 4.875 192.295 ;
      LAYER met4 ;
        RECT 4.555 191.975 4.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 191.570 4.875 191.890 ;
      LAYER met4 ;
        RECT 4.555 191.570 4.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 191.165 4.875 191.485 ;
      LAYER met4 ;
        RECT 4.555 191.165 4.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 190.760 4.875 191.080 ;
      LAYER met4 ;
        RECT 4.555 190.760 4.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 190.355 4.875 190.675 ;
      LAYER met4 ;
        RECT 4.555 190.355 4.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 189.950 4.875 190.270 ;
      LAYER met4 ;
        RECT 4.555 189.950 4.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 189.545 4.875 189.865 ;
      LAYER met4 ;
        RECT 4.555 189.545 4.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 189.140 4.875 189.460 ;
      LAYER met4 ;
        RECT 4.555 189.140 4.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 188.735 4.875 189.055 ;
      LAYER met4 ;
        RECT 4.555 188.735 4.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 188.330 4.875 188.650 ;
      LAYER met4 ;
        RECT 4.555 188.330 4.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 187.925 4.875 188.245 ;
      LAYER met4 ;
        RECT 4.555 187.925 4.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 187.520 4.875 187.840 ;
      LAYER met4 ;
        RECT 4.555 187.520 4.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 187.115 4.875 187.435 ;
      LAYER met4 ;
        RECT 4.555 187.115 4.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 186.710 4.875 187.030 ;
      LAYER met4 ;
        RECT 4.555 186.710 4.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 186.305 4.875 186.625 ;
      LAYER met4 ;
        RECT 4.555 186.305 4.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 185.900 4.875 186.220 ;
      LAYER met4 ;
        RECT 4.555 185.900 4.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 185.495 4.875 185.815 ;
      LAYER met4 ;
        RECT 4.555 185.495 4.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 185.090 4.875 185.410 ;
      LAYER met4 ;
        RECT 4.555 185.090 4.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 184.685 4.875 185.005 ;
      LAYER met4 ;
        RECT 4.555 184.685 4.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 184.280 4.875 184.600 ;
      LAYER met4 ;
        RECT 4.555 184.280 4.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 183.875 4.875 184.195 ;
      LAYER met4 ;
        RECT 4.555 183.875 4.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 183.470 4.875 183.790 ;
      LAYER met4 ;
        RECT 4.555 183.470 4.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 183.065 4.875 183.385 ;
      LAYER met4 ;
        RECT 4.555 183.065 4.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 182.660 4.875 182.980 ;
      LAYER met4 ;
        RECT 4.555 182.660 4.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 182.255 4.875 182.575 ;
      LAYER met4 ;
        RECT 4.555 182.255 4.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 181.850 4.875 182.170 ;
      LAYER met4 ;
        RECT 4.555 181.850 4.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.555 181.445 4.875 181.765 ;
      LAYER met4 ;
        RECT 4.555 181.445 4.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 28.210 4.465 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 27.780 4.465 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 27.350 4.465 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 26.920 4.465 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 26.490 4.465 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 26.060 4.465 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 25.630 4.465 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 25.200 4.465 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 24.770 4.465 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 24.340 4.465 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.265 23.910 4.465 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 197.645 4.475 197.965 ;
      LAYER met4 ;
        RECT 4.155 197.645 4.475 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 197.240 4.475 197.560 ;
      LAYER met4 ;
        RECT 4.155 197.240 4.475 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 196.835 4.475 197.155 ;
      LAYER met4 ;
        RECT 4.155 196.835 4.475 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 196.430 4.475 196.750 ;
      LAYER met4 ;
        RECT 4.155 196.430 4.475 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 196.025 4.475 196.345 ;
      LAYER met4 ;
        RECT 4.155 196.025 4.475 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 195.620 4.475 195.940 ;
      LAYER met4 ;
        RECT 4.155 195.620 4.475 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 195.215 4.475 195.535 ;
      LAYER met4 ;
        RECT 4.155 195.215 4.475 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 194.810 4.475 195.130 ;
      LAYER met4 ;
        RECT 4.155 194.810 4.475 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 194.405 4.475 194.725 ;
      LAYER met4 ;
        RECT 4.155 194.405 4.475 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 194.000 4.475 194.320 ;
      LAYER met4 ;
        RECT 4.155 194.000 4.475 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 193.595 4.475 193.915 ;
      LAYER met4 ;
        RECT 4.155 193.595 4.475 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 193.190 4.475 193.510 ;
      LAYER met4 ;
        RECT 4.155 193.190 4.475 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 192.785 4.475 193.105 ;
      LAYER met4 ;
        RECT 4.155 192.785 4.475 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 192.380 4.475 192.700 ;
      LAYER met4 ;
        RECT 4.155 192.380 4.475 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 191.975 4.475 192.295 ;
      LAYER met4 ;
        RECT 4.155 191.975 4.475 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 191.570 4.475 191.890 ;
      LAYER met4 ;
        RECT 4.155 191.570 4.475 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 191.165 4.475 191.485 ;
      LAYER met4 ;
        RECT 4.155 191.165 4.475 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 190.760 4.475 191.080 ;
      LAYER met4 ;
        RECT 4.155 190.760 4.475 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 190.355 4.475 190.675 ;
      LAYER met4 ;
        RECT 4.155 190.355 4.475 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 189.950 4.475 190.270 ;
      LAYER met4 ;
        RECT 4.155 189.950 4.475 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 189.545 4.475 189.865 ;
      LAYER met4 ;
        RECT 4.155 189.545 4.475 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 189.140 4.475 189.460 ;
      LAYER met4 ;
        RECT 4.155 189.140 4.475 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 188.735 4.475 189.055 ;
      LAYER met4 ;
        RECT 4.155 188.735 4.475 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 188.330 4.475 188.650 ;
      LAYER met4 ;
        RECT 4.155 188.330 4.475 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 187.925 4.475 188.245 ;
      LAYER met4 ;
        RECT 4.155 187.925 4.475 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 187.520 4.475 187.840 ;
      LAYER met4 ;
        RECT 4.155 187.520 4.475 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 187.115 4.475 187.435 ;
      LAYER met4 ;
        RECT 4.155 187.115 4.475 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 186.710 4.475 187.030 ;
      LAYER met4 ;
        RECT 4.155 186.710 4.475 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 186.305 4.475 186.625 ;
      LAYER met4 ;
        RECT 4.155 186.305 4.475 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 185.900 4.475 186.220 ;
      LAYER met4 ;
        RECT 4.155 185.900 4.475 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 185.495 4.475 185.815 ;
      LAYER met4 ;
        RECT 4.155 185.495 4.475 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 185.090 4.475 185.410 ;
      LAYER met4 ;
        RECT 4.155 185.090 4.475 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 184.685 4.475 185.005 ;
      LAYER met4 ;
        RECT 4.155 184.685 4.475 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 184.280 4.475 184.600 ;
      LAYER met4 ;
        RECT 4.155 184.280 4.475 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 183.875 4.475 184.195 ;
      LAYER met4 ;
        RECT 4.155 183.875 4.475 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 183.470 4.475 183.790 ;
      LAYER met4 ;
        RECT 4.155 183.470 4.475 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 183.065 4.475 183.385 ;
      LAYER met4 ;
        RECT 4.155 183.065 4.475 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 182.660 4.475 182.980 ;
      LAYER met4 ;
        RECT 4.155 182.660 4.475 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 182.255 4.475 182.575 ;
      LAYER met4 ;
        RECT 4.155 182.255 4.475 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 181.850 4.475 182.170 ;
      LAYER met4 ;
        RECT 4.155 181.850 4.475 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.155 181.445 4.475 181.765 ;
      LAYER met4 ;
        RECT 4.155 181.445 4.475 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 28.210 4.060 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 27.780 4.060 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 27.350 4.060 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 26.920 4.060 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 26.490 4.060 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 26.060 4.060 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 25.630 4.060 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 25.200 4.060 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 24.770 4.060 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 24.340 4.060 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.860 23.910 4.060 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 197.645 4.075 197.965 ;
      LAYER met4 ;
        RECT 3.755 197.645 4.075 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 197.240 4.075 197.560 ;
      LAYER met4 ;
        RECT 3.755 197.240 4.075 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 196.835 4.075 197.155 ;
      LAYER met4 ;
        RECT 3.755 196.835 4.075 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 196.430 4.075 196.750 ;
      LAYER met4 ;
        RECT 3.755 196.430 4.075 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 196.025 4.075 196.345 ;
      LAYER met4 ;
        RECT 3.755 196.025 4.075 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 195.620 4.075 195.940 ;
      LAYER met4 ;
        RECT 3.755 195.620 4.075 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 195.215 4.075 195.535 ;
      LAYER met4 ;
        RECT 3.755 195.215 4.075 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 194.810 4.075 195.130 ;
      LAYER met4 ;
        RECT 3.755 194.810 4.075 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 194.405 4.075 194.725 ;
      LAYER met4 ;
        RECT 3.755 194.405 4.075 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 194.000 4.075 194.320 ;
      LAYER met4 ;
        RECT 3.755 194.000 4.075 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 193.595 4.075 193.915 ;
      LAYER met4 ;
        RECT 3.755 193.595 4.075 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 193.190 4.075 193.510 ;
      LAYER met4 ;
        RECT 3.755 193.190 4.075 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 192.785 4.075 193.105 ;
      LAYER met4 ;
        RECT 3.755 192.785 4.075 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 192.380 4.075 192.700 ;
      LAYER met4 ;
        RECT 3.755 192.380 4.075 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 191.975 4.075 192.295 ;
      LAYER met4 ;
        RECT 3.755 191.975 4.075 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 191.570 4.075 191.890 ;
      LAYER met4 ;
        RECT 3.755 191.570 4.075 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 191.165 4.075 191.485 ;
      LAYER met4 ;
        RECT 3.755 191.165 4.075 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 190.760 4.075 191.080 ;
      LAYER met4 ;
        RECT 3.755 190.760 4.075 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 190.355 4.075 190.675 ;
      LAYER met4 ;
        RECT 3.755 190.355 4.075 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 189.950 4.075 190.270 ;
      LAYER met4 ;
        RECT 3.755 189.950 4.075 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 189.545 4.075 189.865 ;
      LAYER met4 ;
        RECT 3.755 189.545 4.075 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 189.140 4.075 189.460 ;
      LAYER met4 ;
        RECT 3.755 189.140 4.075 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 188.735 4.075 189.055 ;
      LAYER met4 ;
        RECT 3.755 188.735 4.075 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 188.330 4.075 188.650 ;
      LAYER met4 ;
        RECT 3.755 188.330 4.075 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 187.925 4.075 188.245 ;
      LAYER met4 ;
        RECT 3.755 187.925 4.075 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 187.520 4.075 187.840 ;
      LAYER met4 ;
        RECT 3.755 187.520 4.075 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 187.115 4.075 187.435 ;
      LAYER met4 ;
        RECT 3.755 187.115 4.075 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 186.710 4.075 187.030 ;
      LAYER met4 ;
        RECT 3.755 186.710 4.075 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 186.305 4.075 186.625 ;
      LAYER met4 ;
        RECT 3.755 186.305 4.075 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 185.900 4.075 186.220 ;
      LAYER met4 ;
        RECT 3.755 185.900 4.075 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 185.495 4.075 185.815 ;
      LAYER met4 ;
        RECT 3.755 185.495 4.075 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 185.090 4.075 185.410 ;
      LAYER met4 ;
        RECT 3.755 185.090 4.075 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 184.685 4.075 185.005 ;
      LAYER met4 ;
        RECT 3.755 184.685 4.075 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 184.280 4.075 184.600 ;
      LAYER met4 ;
        RECT 3.755 184.280 4.075 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 183.875 4.075 184.195 ;
      LAYER met4 ;
        RECT 3.755 183.875 4.075 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 183.470 4.075 183.790 ;
      LAYER met4 ;
        RECT 3.755 183.470 4.075 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 183.065 4.075 183.385 ;
      LAYER met4 ;
        RECT 3.755 183.065 4.075 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 182.660 4.075 182.980 ;
      LAYER met4 ;
        RECT 3.755 182.660 4.075 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 182.255 4.075 182.575 ;
      LAYER met4 ;
        RECT 3.755 182.255 4.075 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 181.850 4.075 182.170 ;
      LAYER met4 ;
        RECT 3.755 181.850 4.075 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.755 181.445 4.075 181.765 ;
      LAYER met4 ;
        RECT 3.755 181.445 4.075 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 28.210 3.655 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 27.780 3.655 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 27.350 3.655 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 26.920 3.655 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 26.490 3.655 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 26.060 3.655 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 25.630 3.655 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 25.200 3.655 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 24.770 3.655 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 24.340 3.655 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.455 23.910 3.655 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 197.645 3.675 197.965 ;
      LAYER met4 ;
        RECT 3.355 197.645 3.675 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 197.240 3.675 197.560 ;
      LAYER met4 ;
        RECT 3.355 197.240 3.675 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 196.835 3.675 197.155 ;
      LAYER met4 ;
        RECT 3.355 196.835 3.675 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 196.430 3.675 196.750 ;
      LAYER met4 ;
        RECT 3.355 196.430 3.675 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 196.025 3.675 196.345 ;
      LAYER met4 ;
        RECT 3.355 196.025 3.675 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 195.620 3.675 195.940 ;
      LAYER met4 ;
        RECT 3.355 195.620 3.675 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 195.215 3.675 195.535 ;
      LAYER met4 ;
        RECT 3.355 195.215 3.675 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 194.810 3.675 195.130 ;
      LAYER met4 ;
        RECT 3.355 194.810 3.675 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 194.405 3.675 194.725 ;
      LAYER met4 ;
        RECT 3.355 194.405 3.675 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 194.000 3.675 194.320 ;
      LAYER met4 ;
        RECT 3.355 194.000 3.675 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 193.595 3.675 193.915 ;
      LAYER met4 ;
        RECT 3.355 193.595 3.675 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 193.190 3.675 193.510 ;
      LAYER met4 ;
        RECT 3.355 193.190 3.675 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 192.785 3.675 193.105 ;
      LAYER met4 ;
        RECT 3.355 192.785 3.675 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 192.380 3.675 192.700 ;
      LAYER met4 ;
        RECT 3.355 192.380 3.675 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 191.975 3.675 192.295 ;
      LAYER met4 ;
        RECT 3.355 191.975 3.675 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 191.570 3.675 191.890 ;
      LAYER met4 ;
        RECT 3.355 191.570 3.675 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 191.165 3.675 191.485 ;
      LAYER met4 ;
        RECT 3.355 191.165 3.675 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 190.760 3.675 191.080 ;
      LAYER met4 ;
        RECT 3.355 190.760 3.675 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 190.355 3.675 190.675 ;
      LAYER met4 ;
        RECT 3.355 190.355 3.675 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 189.950 3.675 190.270 ;
      LAYER met4 ;
        RECT 3.355 189.950 3.675 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 189.545 3.675 189.865 ;
      LAYER met4 ;
        RECT 3.355 189.545 3.675 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 189.140 3.675 189.460 ;
      LAYER met4 ;
        RECT 3.355 189.140 3.675 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 188.735 3.675 189.055 ;
      LAYER met4 ;
        RECT 3.355 188.735 3.675 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 188.330 3.675 188.650 ;
      LAYER met4 ;
        RECT 3.355 188.330 3.675 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 187.925 3.675 188.245 ;
      LAYER met4 ;
        RECT 3.355 187.925 3.675 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 187.520 3.675 187.840 ;
      LAYER met4 ;
        RECT 3.355 187.520 3.675 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 187.115 3.675 187.435 ;
      LAYER met4 ;
        RECT 3.355 187.115 3.675 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 186.710 3.675 187.030 ;
      LAYER met4 ;
        RECT 3.355 186.710 3.675 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 186.305 3.675 186.625 ;
      LAYER met4 ;
        RECT 3.355 186.305 3.675 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 185.900 3.675 186.220 ;
      LAYER met4 ;
        RECT 3.355 185.900 3.675 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 185.495 3.675 185.815 ;
      LAYER met4 ;
        RECT 3.355 185.495 3.675 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 185.090 3.675 185.410 ;
      LAYER met4 ;
        RECT 3.355 185.090 3.675 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 184.685 3.675 185.005 ;
      LAYER met4 ;
        RECT 3.355 184.685 3.675 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 184.280 3.675 184.600 ;
      LAYER met4 ;
        RECT 3.355 184.280 3.675 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 183.875 3.675 184.195 ;
      LAYER met4 ;
        RECT 3.355 183.875 3.675 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 183.470 3.675 183.790 ;
      LAYER met4 ;
        RECT 3.355 183.470 3.675 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 183.065 3.675 183.385 ;
      LAYER met4 ;
        RECT 3.355 183.065 3.675 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 182.660 3.675 182.980 ;
      LAYER met4 ;
        RECT 3.355 182.660 3.675 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 182.255 3.675 182.575 ;
      LAYER met4 ;
        RECT 3.355 182.255 3.675 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 181.850 3.675 182.170 ;
      LAYER met4 ;
        RECT 3.355 181.850 3.675 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.355 181.445 3.675 181.765 ;
      LAYER met4 ;
        RECT 3.355 181.445 3.675 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 28.210 3.250 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 27.780 3.250 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 27.350 3.250 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 26.920 3.250 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 26.490 3.250 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 26.060 3.250 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 25.630 3.250 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 25.200 3.250 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 24.770 3.250 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 24.340 3.250 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.050 23.910 3.250 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 197.645 3.275 197.965 ;
      LAYER met4 ;
        RECT 2.955 197.645 3.275 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 197.240 3.275 197.560 ;
      LAYER met4 ;
        RECT 2.955 197.240 3.275 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 196.835 3.275 197.155 ;
      LAYER met4 ;
        RECT 2.955 196.835 3.275 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 196.430 3.275 196.750 ;
      LAYER met4 ;
        RECT 2.955 196.430 3.275 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 196.025 3.275 196.345 ;
      LAYER met4 ;
        RECT 2.955 196.025 3.275 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 195.620 3.275 195.940 ;
      LAYER met4 ;
        RECT 2.955 195.620 3.275 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 195.215 3.275 195.535 ;
      LAYER met4 ;
        RECT 2.955 195.215 3.275 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 194.810 3.275 195.130 ;
      LAYER met4 ;
        RECT 2.955 194.810 3.275 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 194.405 3.275 194.725 ;
      LAYER met4 ;
        RECT 2.955 194.405 3.275 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 194.000 3.275 194.320 ;
      LAYER met4 ;
        RECT 2.955 194.000 3.275 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 193.595 3.275 193.915 ;
      LAYER met4 ;
        RECT 2.955 193.595 3.275 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 193.190 3.275 193.510 ;
      LAYER met4 ;
        RECT 2.955 193.190 3.275 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 192.785 3.275 193.105 ;
      LAYER met4 ;
        RECT 2.955 192.785 3.275 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 192.380 3.275 192.700 ;
      LAYER met4 ;
        RECT 2.955 192.380 3.275 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 191.975 3.275 192.295 ;
      LAYER met4 ;
        RECT 2.955 191.975 3.275 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 191.570 3.275 191.890 ;
      LAYER met4 ;
        RECT 2.955 191.570 3.275 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 191.165 3.275 191.485 ;
      LAYER met4 ;
        RECT 2.955 191.165 3.275 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 190.760 3.275 191.080 ;
      LAYER met4 ;
        RECT 2.955 190.760 3.275 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 190.355 3.275 190.675 ;
      LAYER met4 ;
        RECT 2.955 190.355 3.275 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 189.950 3.275 190.270 ;
      LAYER met4 ;
        RECT 2.955 189.950 3.275 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 189.545 3.275 189.865 ;
      LAYER met4 ;
        RECT 2.955 189.545 3.275 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 189.140 3.275 189.460 ;
      LAYER met4 ;
        RECT 2.955 189.140 3.275 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 188.735 3.275 189.055 ;
      LAYER met4 ;
        RECT 2.955 188.735 3.275 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 188.330 3.275 188.650 ;
      LAYER met4 ;
        RECT 2.955 188.330 3.275 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 187.925 3.275 188.245 ;
      LAYER met4 ;
        RECT 2.955 187.925 3.275 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 187.520 3.275 187.840 ;
      LAYER met4 ;
        RECT 2.955 187.520 3.275 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 187.115 3.275 187.435 ;
      LAYER met4 ;
        RECT 2.955 187.115 3.275 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 186.710 3.275 187.030 ;
      LAYER met4 ;
        RECT 2.955 186.710 3.275 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 186.305 3.275 186.625 ;
      LAYER met4 ;
        RECT 2.955 186.305 3.275 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 185.900 3.275 186.220 ;
      LAYER met4 ;
        RECT 2.955 185.900 3.275 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 185.495 3.275 185.815 ;
      LAYER met4 ;
        RECT 2.955 185.495 3.275 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 185.090 3.275 185.410 ;
      LAYER met4 ;
        RECT 2.955 185.090 3.275 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 184.685 3.275 185.005 ;
      LAYER met4 ;
        RECT 2.955 184.685 3.275 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 184.280 3.275 184.600 ;
      LAYER met4 ;
        RECT 2.955 184.280 3.275 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 183.875 3.275 184.195 ;
      LAYER met4 ;
        RECT 2.955 183.875 3.275 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 183.470 3.275 183.790 ;
      LAYER met4 ;
        RECT 2.955 183.470 3.275 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 183.065 3.275 183.385 ;
      LAYER met4 ;
        RECT 2.955 183.065 3.275 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 182.660 3.275 182.980 ;
      LAYER met4 ;
        RECT 2.955 182.660 3.275 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 182.255 3.275 182.575 ;
      LAYER met4 ;
        RECT 2.955 182.255 3.275 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 181.850 3.275 182.170 ;
      LAYER met4 ;
        RECT 2.955 181.850 3.275 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.955 181.445 3.275 181.765 ;
      LAYER met4 ;
        RECT 2.955 181.445 3.275 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 28.210 2.840 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 27.780 2.840 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 27.350 2.840 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 26.920 2.840 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 26.490 2.840 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 26.060 2.840 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 25.630 2.840 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 25.200 2.840 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 24.770 2.840 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 24.340 2.840 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.640 23.910 2.840 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 197.645 2.875 197.965 ;
      LAYER met4 ;
        RECT 2.555 197.645 2.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 197.240 2.875 197.560 ;
      LAYER met4 ;
        RECT 2.555 197.240 2.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 196.835 2.875 197.155 ;
      LAYER met4 ;
        RECT 2.555 196.835 2.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 196.430 2.875 196.750 ;
      LAYER met4 ;
        RECT 2.555 196.430 2.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 196.025 2.875 196.345 ;
      LAYER met4 ;
        RECT 2.555 196.025 2.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 195.620 2.875 195.940 ;
      LAYER met4 ;
        RECT 2.555 195.620 2.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 195.215 2.875 195.535 ;
      LAYER met4 ;
        RECT 2.555 195.215 2.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 194.810 2.875 195.130 ;
      LAYER met4 ;
        RECT 2.555 194.810 2.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 194.405 2.875 194.725 ;
      LAYER met4 ;
        RECT 2.555 194.405 2.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 194.000 2.875 194.320 ;
      LAYER met4 ;
        RECT 2.555 194.000 2.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 193.595 2.875 193.915 ;
      LAYER met4 ;
        RECT 2.555 193.595 2.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 193.190 2.875 193.510 ;
      LAYER met4 ;
        RECT 2.555 193.190 2.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 192.785 2.875 193.105 ;
      LAYER met4 ;
        RECT 2.555 192.785 2.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 192.380 2.875 192.700 ;
      LAYER met4 ;
        RECT 2.555 192.380 2.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 191.975 2.875 192.295 ;
      LAYER met4 ;
        RECT 2.555 191.975 2.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 191.570 2.875 191.890 ;
      LAYER met4 ;
        RECT 2.555 191.570 2.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 191.165 2.875 191.485 ;
      LAYER met4 ;
        RECT 2.555 191.165 2.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 190.760 2.875 191.080 ;
      LAYER met4 ;
        RECT 2.555 190.760 2.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 190.355 2.875 190.675 ;
      LAYER met4 ;
        RECT 2.555 190.355 2.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 189.950 2.875 190.270 ;
      LAYER met4 ;
        RECT 2.555 189.950 2.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 189.545 2.875 189.865 ;
      LAYER met4 ;
        RECT 2.555 189.545 2.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 189.140 2.875 189.460 ;
      LAYER met4 ;
        RECT 2.555 189.140 2.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 188.735 2.875 189.055 ;
      LAYER met4 ;
        RECT 2.555 188.735 2.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 188.330 2.875 188.650 ;
      LAYER met4 ;
        RECT 2.555 188.330 2.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 187.925 2.875 188.245 ;
      LAYER met4 ;
        RECT 2.555 187.925 2.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 187.520 2.875 187.840 ;
      LAYER met4 ;
        RECT 2.555 187.520 2.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 187.115 2.875 187.435 ;
      LAYER met4 ;
        RECT 2.555 187.115 2.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 186.710 2.875 187.030 ;
      LAYER met4 ;
        RECT 2.555 186.710 2.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 186.305 2.875 186.625 ;
      LAYER met4 ;
        RECT 2.555 186.305 2.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 185.900 2.875 186.220 ;
      LAYER met4 ;
        RECT 2.555 185.900 2.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 185.495 2.875 185.815 ;
      LAYER met4 ;
        RECT 2.555 185.495 2.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 185.090 2.875 185.410 ;
      LAYER met4 ;
        RECT 2.555 185.090 2.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 184.685 2.875 185.005 ;
      LAYER met4 ;
        RECT 2.555 184.685 2.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 184.280 2.875 184.600 ;
      LAYER met4 ;
        RECT 2.555 184.280 2.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 183.875 2.875 184.195 ;
      LAYER met4 ;
        RECT 2.555 183.875 2.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 183.470 2.875 183.790 ;
      LAYER met4 ;
        RECT 2.555 183.470 2.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 183.065 2.875 183.385 ;
      LAYER met4 ;
        RECT 2.555 183.065 2.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 182.660 2.875 182.980 ;
      LAYER met4 ;
        RECT 2.555 182.660 2.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 182.255 2.875 182.575 ;
      LAYER met4 ;
        RECT 2.555 182.255 2.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 181.850 2.875 182.170 ;
      LAYER met4 ;
        RECT 2.555 181.850 2.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 181.445 2.875 181.765 ;
      LAYER met4 ;
        RECT 2.555 181.445 2.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 28.210 2.430 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 27.780 2.430 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 27.350 2.430 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 26.920 2.430 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 26.490 2.430 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 26.060 2.430 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 25.630 2.430 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 25.200 2.430 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 24.770 2.430 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 24.340 2.430 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.230 23.910 2.430 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 197.645 2.475 197.965 ;
      LAYER met4 ;
        RECT 2.155 197.645 2.475 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 197.240 2.475 197.560 ;
      LAYER met4 ;
        RECT 2.155 197.240 2.475 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 196.835 2.475 197.155 ;
      LAYER met4 ;
        RECT 2.155 196.835 2.475 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 196.430 2.475 196.750 ;
      LAYER met4 ;
        RECT 2.155 196.430 2.475 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 196.025 2.475 196.345 ;
      LAYER met4 ;
        RECT 2.155 196.025 2.475 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 195.620 2.475 195.940 ;
      LAYER met4 ;
        RECT 2.155 195.620 2.475 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 195.215 2.475 195.535 ;
      LAYER met4 ;
        RECT 2.155 195.215 2.475 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 194.810 2.475 195.130 ;
      LAYER met4 ;
        RECT 2.155 194.810 2.475 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 194.405 2.475 194.725 ;
      LAYER met4 ;
        RECT 2.155 194.405 2.475 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 194.000 2.475 194.320 ;
      LAYER met4 ;
        RECT 2.155 194.000 2.475 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 193.595 2.475 193.915 ;
      LAYER met4 ;
        RECT 2.155 193.595 2.475 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 193.190 2.475 193.510 ;
      LAYER met4 ;
        RECT 2.155 193.190 2.475 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 192.785 2.475 193.105 ;
      LAYER met4 ;
        RECT 2.155 192.785 2.475 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 192.380 2.475 192.700 ;
      LAYER met4 ;
        RECT 2.155 192.380 2.475 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 191.975 2.475 192.295 ;
      LAYER met4 ;
        RECT 2.155 191.975 2.475 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 191.570 2.475 191.890 ;
      LAYER met4 ;
        RECT 2.155 191.570 2.475 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 191.165 2.475 191.485 ;
      LAYER met4 ;
        RECT 2.155 191.165 2.475 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 190.760 2.475 191.080 ;
      LAYER met4 ;
        RECT 2.155 190.760 2.475 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 190.355 2.475 190.675 ;
      LAYER met4 ;
        RECT 2.155 190.355 2.475 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 189.950 2.475 190.270 ;
      LAYER met4 ;
        RECT 2.155 189.950 2.475 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 189.545 2.475 189.865 ;
      LAYER met4 ;
        RECT 2.155 189.545 2.475 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 189.140 2.475 189.460 ;
      LAYER met4 ;
        RECT 2.155 189.140 2.475 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 188.735 2.475 189.055 ;
      LAYER met4 ;
        RECT 2.155 188.735 2.475 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 188.330 2.475 188.650 ;
      LAYER met4 ;
        RECT 2.155 188.330 2.475 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 187.925 2.475 188.245 ;
      LAYER met4 ;
        RECT 2.155 187.925 2.475 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 187.520 2.475 187.840 ;
      LAYER met4 ;
        RECT 2.155 187.520 2.475 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 187.115 2.475 187.435 ;
      LAYER met4 ;
        RECT 2.155 187.115 2.475 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 186.710 2.475 187.030 ;
      LAYER met4 ;
        RECT 2.155 186.710 2.475 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 186.305 2.475 186.625 ;
      LAYER met4 ;
        RECT 2.155 186.305 2.475 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 185.900 2.475 186.220 ;
      LAYER met4 ;
        RECT 2.155 185.900 2.475 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 185.495 2.475 185.815 ;
      LAYER met4 ;
        RECT 2.155 185.495 2.475 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 185.090 2.475 185.410 ;
      LAYER met4 ;
        RECT 2.155 185.090 2.475 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 184.685 2.475 185.005 ;
      LAYER met4 ;
        RECT 2.155 184.685 2.475 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 184.280 2.475 184.600 ;
      LAYER met4 ;
        RECT 2.155 184.280 2.475 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 183.875 2.475 184.195 ;
      LAYER met4 ;
        RECT 2.155 183.875 2.475 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 183.470 2.475 183.790 ;
      LAYER met4 ;
        RECT 2.155 183.470 2.475 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 183.065 2.475 183.385 ;
      LAYER met4 ;
        RECT 2.155 183.065 2.475 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 182.660 2.475 182.980 ;
      LAYER met4 ;
        RECT 2.155 182.660 2.475 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 182.255 2.475 182.575 ;
      LAYER met4 ;
        RECT 2.155 182.255 2.475 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 181.850 2.475 182.170 ;
      LAYER met4 ;
        RECT 2.155 181.850 2.475 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.155 181.445 2.475 181.765 ;
      LAYER met4 ;
        RECT 2.155 181.445 2.475 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 28.210 2.020 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 27.780 2.020 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 27.350 2.020 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 26.920 2.020 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 26.490 2.020 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 26.060 2.020 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 25.630 2.020 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 25.200 2.020 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 24.770 2.020 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 24.340 2.020 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.820 23.910 2.020 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 197.645 2.075 197.965 ;
      LAYER met4 ;
        RECT 1.755 197.645 2.075 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 197.240 2.075 197.560 ;
      LAYER met4 ;
        RECT 1.755 197.240 2.075 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 196.835 2.075 197.155 ;
      LAYER met4 ;
        RECT 1.755 196.835 2.075 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 196.430 2.075 196.750 ;
      LAYER met4 ;
        RECT 1.755 196.430 2.075 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 196.025 2.075 196.345 ;
      LAYER met4 ;
        RECT 1.755 196.025 2.075 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 195.620 2.075 195.940 ;
      LAYER met4 ;
        RECT 1.755 195.620 2.075 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 195.215 2.075 195.535 ;
      LAYER met4 ;
        RECT 1.755 195.215 2.075 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 194.810 2.075 195.130 ;
      LAYER met4 ;
        RECT 1.755 194.810 2.075 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 194.405 2.075 194.725 ;
      LAYER met4 ;
        RECT 1.755 194.405 2.075 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 194.000 2.075 194.320 ;
      LAYER met4 ;
        RECT 1.755 194.000 2.075 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 193.595 2.075 193.915 ;
      LAYER met4 ;
        RECT 1.755 193.595 2.075 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 193.190 2.075 193.510 ;
      LAYER met4 ;
        RECT 1.755 193.190 2.075 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 192.785 2.075 193.105 ;
      LAYER met4 ;
        RECT 1.755 192.785 2.075 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 192.380 2.075 192.700 ;
      LAYER met4 ;
        RECT 1.755 192.380 2.075 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 191.975 2.075 192.295 ;
      LAYER met4 ;
        RECT 1.755 191.975 2.075 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 191.570 2.075 191.890 ;
      LAYER met4 ;
        RECT 1.755 191.570 2.075 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 191.165 2.075 191.485 ;
      LAYER met4 ;
        RECT 1.755 191.165 2.075 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 190.760 2.075 191.080 ;
      LAYER met4 ;
        RECT 1.755 190.760 2.075 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 190.355 2.075 190.675 ;
      LAYER met4 ;
        RECT 1.755 190.355 2.075 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 189.950 2.075 190.270 ;
      LAYER met4 ;
        RECT 1.755 189.950 2.075 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 189.545 2.075 189.865 ;
      LAYER met4 ;
        RECT 1.755 189.545 2.075 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 189.140 2.075 189.460 ;
      LAYER met4 ;
        RECT 1.755 189.140 2.075 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 188.735 2.075 189.055 ;
      LAYER met4 ;
        RECT 1.755 188.735 2.075 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 188.330 2.075 188.650 ;
      LAYER met4 ;
        RECT 1.755 188.330 2.075 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 187.925 2.075 188.245 ;
      LAYER met4 ;
        RECT 1.755 187.925 2.075 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 187.520 2.075 187.840 ;
      LAYER met4 ;
        RECT 1.755 187.520 2.075 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 187.115 2.075 187.435 ;
      LAYER met4 ;
        RECT 1.755 187.115 2.075 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 186.710 2.075 187.030 ;
      LAYER met4 ;
        RECT 1.755 186.710 2.075 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 186.305 2.075 186.625 ;
      LAYER met4 ;
        RECT 1.755 186.305 2.075 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 185.900 2.075 186.220 ;
      LAYER met4 ;
        RECT 1.755 185.900 2.075 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 185.495 2.075 185.815 ;
      LAYER met4 ;
        RECT 1.755 185.495 2.075 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 185.090 2.075 185.410 ;
      LAYER met4 ;
        RECT 1.755 185.090 2.075 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 184.685 2.075 185.005 ;
      LAYER met4 ;
        RECT 1.755 184.685 2.075 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 184.280 2.075 184.600 ;
      LAYER met4 ;
        RECT 1.755 184.280 2.075 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 183.875 2.075 184.195 ;
      LAYER met4 ;
        RECT 1.755 183.875 2.075 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 183.470 2.075 183.790 ;
      LAYER met4 ;
        RECT 1.755 183.470 2.075 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 183.065 2.075 183.385 ;
      LAYER met4 ;
        RECT 1.755 183.065 2.075 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 182.660 2.075 182.980 ;
      LAYER met4 ;
        RECT 1.755 182.660 2.075 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 182.255 2.075 182.575 ;
      LAYER met4 ;
        RECT 1.755 182.255 2.075 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 181.850 2.075 182.170 ;
      LAYER met4 ;
        RECT 1.755 181.850 2.075 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.755 181.445 2.075 181.765 ;
      LAYER met4 ;
        RECT 1.755 181.445 2.075 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 197.645 1.675 197.965 ;
      LAYER met4 ;
        RECT 1.355 197.645 1.675 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 197.240 1.675 197.560 ;
      LAYER met4 ;
        RECT 1.355 197.240 1.675 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 196.835 1.675 197.155 ;
      LAYER met4 ;
        RECT 1.355 196.835 1.675 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 196.430 1.675 196.750 ;
      LAYER met4 ;
        RECT 1.355 196.430 1.675 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 196.025 1.675 196.345 ;
      LAYER met4 ;
        RECT 1.355 196.025 1.675 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 195.620 1.675 195.940 ;
      LAYER met4 ;
        RECT 1.355 195.620 1.675 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 195.215 1.675 195.535 ;
      LAYER met4 ;
        RECT 1.355 195.215 1.675 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 194.810 1.675 195.130 ;
      LAYER met4 ;
        RECT 1.355 194.810 1.675 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 194.405 1.675 194.725 ;
      LAYER met4 ;
        RECT 1.355 194.405 1.675 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 194.000 1.675 194.320 ;
      LAYER met4 ;
        RECT 1.355 194.000 1.675 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 193.595 1.675 193.915 ;
      LAYER met4 ;
        RECT 1.355 193.595 1.675 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 193.190 1.675 193.510 ;
      LAYER met4 ;
        RECT 1.355 193.190 1.675 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 192.785 1.675 193.105 ;
      LAYER met4 ;
        RECT 1.355 192.785 1.675 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 192.380 1.675 192.700 ;
      LAYER met4 ;
        RECT 1.355 192.380 1.675 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 191.975 1.675 192.295 ;
      LAYER met4 ;
        RECT 1.355 191.975 1.675 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 191.570 1.675 191.890 ;
      LAYER met4 ;
        RECT 1.355 191.570 1.675 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 191.165 1.675 191.485 ;
      LAYER met4 ;
        RECT 1.355 191.165 1.675 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 190.760 1.675 191.080 ;
      LAYER met4 ;
        RECT 1.355 190.760 1.675 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 190.355 1.675 190.675 ;
      LAYER met4 ;
        RECT 1.355 190.355 1.675 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 189.950 1.675 190.270 ;
      LAYER met4 ;
        RECT 1.355 189.950 1.675 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 189.545 1.675 189.865 ;
      LAYER met4 ;
        RECT 1.355 189.545 1.675 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 189.140 1.675 189.460 ;
      LAYER met4 ;
        RECT 1.355 189.140 1.675 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 188.735 1.675 189.055 ;
      LAYER met4 ;
        RECT 1.355 188.735 1.675 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 188.330 1.675 188.650 ;
      LAYER met4 ;
        RECT 1.355 188.330 1.675 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 187.925 1.675 188.245 ;
      LAYER met4 ;
        RECT 1.355 187.925 1.675 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 187.520 1.675 187.840 ;
      LAYER met4 ;
        RECT 1.355 187.520 1.675 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 187.115 1.675 187.435 ;
      LAYER met4 ;
        RECT 1.355 187.115 1.675 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 186.710 1.675 187.030 ;
      LAYER met4 ;
        RECT 1.355 186.710 1.675 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 186.305 1.675 186.625 ;
      LAYER met4 ;
        RECT 1.355 186.305 1.675 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 185.900 1.675 186.220 ;
      LAYER met4 ;
        RECT 1.355 185.900 1.675 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 185.495 1.675 185.815 ;
      LAYER met4 ;
        RECT 1.355 185.495 1.675 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 185.090 1.675 185.410 ;
      LAYER met4 ;
        RECT 1.355 185.090 1.675 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 184.685 1.675 185.005 ;
      LAYER met4 ;
        RECT 1.355 184.685 1.675 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 184.280 1.675 184.600 ;
      LAYER met4 ;
        RECT 1.355 184.280 1.675 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 183.875 1.675 184.195 ;
      LAYER met4 ;
        RECT 1.355 183.875 1.675 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 183.470 1.675 183.790 ;
      LAYER met4 ;
        RECT 1.355 183.470 1.675 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 183.065 1.675 183.385 ;
      LAYER met4 ;
        RECT 1.355 183.065 1.675 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 182.660 1.675 182.980 ;
      LAYER met4 ;
        RECT 1.355 182.660 1.675 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 182.255 1.675 182.575 ;
      LAYER met4 ;
        RECT 1.355 182.255 1.675 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 181.850 1.675 182.170 ;
      LAYER met4 ;
        RECT 1.355 181.850 1.675 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.355 181.445 1.675 181.765 ;
      LAYER met4 ;
        RECT 1.355 181.445 1.675 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 28.210 1.610 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 27.780 1.610 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 27.350 1.610 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 26.920 1.610 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 26.490 1.610 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 26.060 1.610 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 25.630 1.610 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 25.200 1.610 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 24.770 1.610 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 24.340 1.610 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.410 23.910 1.610 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 197.645 1.275 197.965 ;
      LAYER met4 ;
        RECT 1.270 197.645 1.275 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 197.240 1.275 197.560 ;
      LAYER met4 ;
        RECT 1.270 197.240 1.275 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 196.835 1.275 197.155 ;
      LAYER met4 ;
        RECT 1.270 196.835 1.275 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 196.430 1.275 196.750 ;
      LAYER met4 ;
        RECT 1.270 196.430 1.275 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 196.025 1.275 196.345 ;
      LAYER met4 ;
        RECT 1.270 196.025 1.275 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 195.620 1.275 195.940 ;
      LAYER met4 ;
        RECT 1.270 195.620 1.275 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 195.215 1.275 195.535 ;
      LAYER met4 ;
        RECT 1.270 195.215 1.275 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 194.810 1.275 195.130 ;
      LAYER met4 ;
        RECT 1.270 194.810 1.275 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 194.405 1.275 194.725 ;
      LAYER met4 ;
        RECT 1.270 194.405 1.275 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 194.000 1.275 194.320 ;
      LAYER met4 ;
        RECT 1.270 194.000 1.275 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 193.595 1.275 193.915 ;
      LAYER met4 ;
        RECT 1.270 193.595 1.275 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 193.190 1.275 193.510 ;
      LAYER met4 ;
        RECT 1.270 193.190 1.275 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 192.785 1.275 193.105 ;
      LAYER met4 ;
        RECT 1.270 192.785 1.275 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 192.380 1.275 192.700 ;
      LAYER met4 ;
        RECT 1.270 192.380 1.275 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 191.975 1.275 192.295 ;
      LAYER met4 ;
        RECT 1.270 191.975 1.275 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 191.570 1.275 191.890 ;
      LAYER met4 ;
        RECT 1.270 191.570 1.275 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 191.165 1.275 191.485 ;
      LAYER met4 ;
        RECT 1.270 191.165 1.275 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 190.760 1.275 191.080 ;
      LAYER met4 ;
        RECT 1.270 190.760 1.275 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 190.355 1.275 190.675 ;
      LAYER met4 ;
        RECT 1.270 190.355 1.275 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 189.950 1.275 190.270 ;
      LAYER met4 ;
        RECT 1.270 189.950 1.275 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 189.545 1.275 189.865 ;
      LAYER met4 ;
        RECT 1.270 189.545 1.275 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 189.140 1.275 189.460 ;
      LAYER met4 ;
        RECT 1.270 189.140 1.275 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 188.735 1.275 189.055 ;
      LAYER met4 ;
        RECT 1.270 188.735 1.275 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 188.330 1.275 188.650 ;
      LAYER met4 ;
        RECT 1.270 188.330 1.275 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 187.925 1.275 188.245 ;
      LAYER met4 ;
        RECT 1.270 187.925 1.275 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 187.520 1.275 187.840 ;
      LAYER met4 ;
        RECT 1.270 187.520 1.275 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 187.115 1.275 187.435 ;
      LAYER met4 ;
        RECT 1.270 187.115 1.275 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 186.710 1.275 187.030 ;
      LAYER met4 ;
        RECT 1.270 186.710 1.275 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 186.305 1.275 186.625 ;
      LAYER met4 ;
        RECT 1.270 186.305 1.275 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 185.900 1.275 186.220 ;
      LAYER met4 ;
        RECT 1.270 185.900 1.275 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 185.495 1.275 185.815 ;
      LAYER met4 ;
        RECT 1.270 185.495 1.275 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 185.090 1.275 185.410 ;
      LAYER met4 ;
        RECT 1.270 185.090 1.275 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 184.685 1.275 185.005 ;
      LAYER met4 ;
        RECT 1.270 184.685 1.275 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 184.280 1.275 184.600 ;
      LAYER met4 ;
        RECT 1.270 184.280 1.275 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 183.875 1.275 184.195 ;
      LAYER met4 ;
        RECT 1.270 183.875 1.275 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 183.470 1.275 183.790 ;
      LAYER met4 ;
        RECT 1.270 183.470 1.275 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 183.065 1.275 183.385 ;
      LAYER met4 ;
        RECT 1.270 183.065 1.275 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 182.660 1.275 182.980 ;
      LAYER met4 ;
        RECT 1.270 182.660 1.275 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 182.255 1.275 182.575 ;
      LAYER met4 ;
        RECT 1.270 182.255 1.275 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 181.850 1.275 182.170 ;
      LAYER met4 ;
        RECT 1.270 181.850 1.275 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.955 181.445 1.275 181.765 ;
      LAYER met4 ;
        RECT 1.270 181.445 1.275 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 28.210 1.200 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 27.780 1.200 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 27.350 1.200 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 26.920 1.200 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 26.490 1.200 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 26.060 1.200 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 25.630 1.200 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 25.200 1.200 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 24.770 1.200 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 24.340 1.200 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.000 23.910 1.200 24.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 197.645 0.875 197.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 197.240 0.875 197.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 196.835 0.875 197.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 196.430 0.875 196.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 196.025 0.875 196.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 195.620 0.875 195.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 195.215 0.875 195.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 194.810 0.875 195.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 194.405 0.875 194.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 194.000 0.875 194.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 193.595 0.875 193.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 193.190 0.875 193.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 192.785 0.875 193.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 192.380 0.875 192.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 191.975 0.875 192.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 191.570 0.875 191.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 191.165 0.875 191.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 190.760 0.875 191.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 190.355 0.875 190.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 189.950 0.875 190.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 189.545 0.875 189.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 189.140 0.875 189.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 188.735 0.875 189.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 188.330 0.875 188.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 187.925 0.875 188.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 187.520 0.875 187.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 187.115 0.875 187.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 186.710 0.875 187.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 186.305 0.875 186.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 185.900 0.875 186.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 185.495 0.875 185.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 185.090 0.875 185.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 184.685 0.875 185.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 184.280 0.875 184.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 183.875 0.875 184.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 183.470 0.875 183.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 183.065 0.875 183.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 182.660 0.875 182.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 182.255 0.875 182.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 181.850 0.875 182.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.555 181.445 0.875 181.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 28.210 0.790 28.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 27.780 0.790 27.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 27.350 0.790 27.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 26.920 0.790 27.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 26.490 0.790 26.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 26.060 0.790 26.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 25.630 0.790 25.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 25.200 0.790 25.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 24.770 0.790 24.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 24.340 0.790 24.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.590 23.910 0.790 24.110 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.755 56.240 74.290 60.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 60.410 74.200 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 60.000 74.200 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 59.590 74.200 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 59.180 74.200 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 58.770 74.200 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 58.360 74.200 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 57.950 74.200 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 57.540 74.200 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 57.130 74.200 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 56.720 74.200 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.000 56.310 74.200 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 60.410 73.795 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 60.000 73.795 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 59.590 73.795 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 59.180 73.795 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 58.770 73.795 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 58.360 73.795 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 57.950 73.795 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 57.540 73.795 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 57.130 73.795 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 56.720 73.795 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.595 56.310 73.795 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 60.410 73.390 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 60.000 73.390 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 59.590 73.390 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 59.180 73.390 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 58.770 73.390 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 58.360 73.390 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 57.950 73.390 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 57.540 73.390 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 57.130 73.390 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 56.720 73.390 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.190 56.310 73.390 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 60.410 72.985 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 60.000 72.985 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 59.590 72.985 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 59.180 72.985 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 58.770 72.985 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 58.360 72.985 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 57.950 72.985 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 57.540 72.985 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 57.130 72.985 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 56.720 72.985 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.785 56.310 72.985 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 60.410 72.580 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 60.000 72.580 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 59.590 72.580 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 59.180 72.580 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 58.770 72.580 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 58.360 72.580 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 57.950 72.580 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 57.540 72.580 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 57.130 72.580 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 56.720 72.580 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.380 56.310 72.580 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 60.410 72.175 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 60.000 72.175 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 59.590 72.175 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 59.180 72.175 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 58.770 72.175 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 58.360 72.175 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 57.950 72.175 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 57.540 72.175 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 57.130 72.175 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 56.720 72.175 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.975 56.310 72.175 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 60.410 71.770 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 60.000 71.770 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 59.590 71.770 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 59.180 71.770 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 58.770 71.770 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 58.360 71.770 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 57.950 71.770 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 57.540 71.770 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 57.130 71.770 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 56.720 71.770 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.570 56.310 71.770 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 60.410 71.365 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 60.000 71.365 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 59.590 71.365 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 59.180 71.365 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 58.770 71.365 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 58.360 71.365 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 57.950 71.365 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 57.540 71.365 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 57.130 71.365 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 56.720 71.365 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.165 56.310 71.365 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 60.410 70.960 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 60.000 70.960 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 59.590 70.960 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 59.180 70.960 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 58.770 70.960 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 58.360 70.960 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 57.950 70.960 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 57.540 70.960 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 57.130 70.960 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 56.720 70.960 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.760 56.310 70.960 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 60.410 70.555 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 60.000 70.555 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 59.590 70.555 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 59.180 70.555 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 58.770 70.555 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 58.360 70.555 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 57.950 70.555 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 57.540 70.555 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 57.130 70.555 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 56.720 70.555 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.355 56.310 70.555 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 60.410 70.150 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 60.000 70.150 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 59.590 70.150 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 59.180 70.150 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 58.770 70.150 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 58.360 70.150 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 57.950 70.150 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 57.540 70.150 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 57.130 70.150 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 56.720 70.150 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.950 56.310 70.150 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 60.410 69.745 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 60.000 69.745 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 59.590 69.745 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 59.180 69.745 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 58.770 69.745 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 58.360 69.745 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 57.950 69.745 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 57.540 69.745 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 57.130 69.745 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 56.720 69.745 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.545 56.310 69.745 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 60.410 69.340 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 60.000 69.340 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 59.590 69.340 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 59.180 69.340 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 58.770 69.340 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 58.360 69.340 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 57.950 69.340 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 57.540 69.340 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 57.130 69.340 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 56.720 69.340 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.140 56.310 69.340 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 60.410 68.935 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 60.000 68.935 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 59.590 68.935 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 59.180 68.935 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 58.770 68.935 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 58.360 68.935 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 57.950 68.935 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 57.540 68.935 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 57.130 68.935 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 56.720 68.935 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.735 56.310 68.935 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 60.410 68.530 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 60.000 68.530 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 59.590 68.530 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 59.180 68.530 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 58.770 68.530 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 58.360 68.530 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 57.950 68.530 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 57.540 68.530 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 57.130 68.530 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 56.720 68.530 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.330 56.310 68.530 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 60.410 68.125 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 60.000 68.125 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 59.590 68.125 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 59.180 68.125 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 58.770 68.125 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 58.360 68.125 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 57.950 68.125 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 57.540 68.125 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 57.130 68.125 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 56.720 68.125 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.925 56.310 68.125 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 60.410 67.720 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 60.000 67.720 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 59.590 67.720 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 59.180 67.720 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 58.770 67.720 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 58.360 67.720 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 57.950 67.720 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 57.540 67.720 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 57.130 67.720 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 56.720 67.720 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.520 56.310 67.720 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 60.410 67.315 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 60.000 67.315 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 59.590 67.315 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 59.180 67.315 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 58.770 67.315 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 58.360 67.315 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 57.950 67.315 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 57.540 67.315 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 57.130 67.315 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 56.720 67.315 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.115 56.310 67.315 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 60.410 66.910 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 60.000 66.910 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 59.590 66.910 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 59.180 66.910 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 58.770 66.910 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 58.360 66.910 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 57.950 66.910 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 57.540 66.910 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 57.130 66.910 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 56.720 66.910 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.710 56.310 66.910 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 60.410 66.505 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 60.000 66.505 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 59.590 66.505 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 59.180 66.505 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 58.770 66.505 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 58.360 66.505 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 57.950 66.505 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 57.540 66.505 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 57.130 66.505 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 56.720 66.505 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.305 56.310 66.505 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 60.410 66.100 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 60.000 66.100 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 59.590 66.100 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 59.180 66.100 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 58.770 66.100 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 58.360 66.100 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 57.950 66.100 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 57.540 66.100 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 57.130 66.100 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 56.720 66.100 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.900 56.310 66.100 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 60.410 65.695 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 60.000 65.695 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 59.590 65.695 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 59.180 65.695 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 58.770 65.695 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 58.360 65.695 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 57.950 65.695 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 57.540 65.695 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 57.130 65.695 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 56.720 65.695 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.495 56.310 65.695 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 60.410 65.290 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 60.000 65.290 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 59.590 65.290 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 59.180 65.290 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 58.770 65.290 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 58.360 65.290 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 57.950 65.290 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 57.540 65.290 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 57.130 65.290 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 56.720 65.290 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.090 56.310 65.290 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 60.410 64.885 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 60.000 64.885 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 59.590 64.885 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 59.180 64.885 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 58.770 64.885 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 58.360 64.885 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 57.950 64.885 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 57.540 64.885 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 57.130 64.885 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 56.720 64.885 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.685 56.310 64.885 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 60.410 64.480 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 60.000 64.480 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 59.590 64.480 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 59.180 64.480 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 58.770 64.480 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 58.360 64.480 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 57.950 64.480 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 57.540 64.480 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 57.130 64.480 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 56.720 64.480 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.280 56.310 64.480 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 60.410 64.075 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 60.000 64.075 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 59.590 64.075 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 59.180 64.075 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 58.770 64.075 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 58.360 64.075 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 57.950 64.075 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 57.540 64.075 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 57.130 64.075 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 56.720 64.075 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.875 56.310 64.075 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 60.410 63.670 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 60.000 63.670 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 59.590 63.670 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 59.180 63.670 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 58.770 63.670 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 58.360 63.670 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 57.950 63.670 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 57.540 63.670 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 57.130 63.670 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 56.720 63.670 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.470 56.310 63.670 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 60.410 63.265 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 60.000 63.265 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 59.590 63.265 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 59.180 63.265 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 58.770 63.265 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 58.360 63.265 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 57.950 63.265 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 57.540 63.265 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 57.130 63.265 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 56.720 63.265 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.065 56.310 63.265 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 60.410 62.860 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 60.000 62.860 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 59.590 62.860 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 59.180 62.860 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 58.770 62.860 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 58.360 62.860 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 57.950 62.860 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 57.540 62.860 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 57.130 62.860 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 56.720 62.860 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.660 56.310 62.860 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 60.410 62.455 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 60.000 62.455 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 59.590 62.455 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 59.180 62.455 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 58.770 62.455 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 58.360 62.455 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 57.950 62.455 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 57.540 62.455 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 57.130 62.455 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 56.720 62.455 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.255 56.310 62.455 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 60.410 62.050 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 60.000 62.050 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 59.590 62.050 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 59.180 62.050 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 58.770 62.050 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 58.360 62.050 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 57.950 62.050 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 57.540 62.050 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 57.130 62.050 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 56.720 62.050 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.850 56.310 62.050 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 60.410 61.645 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 60.000 61.645 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 59.590 61.645 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 59.180 61.645 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 58.770 61.645 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 58.360 61.645 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 57.950 61.645 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 57.540 61.645 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 57.130 61.645 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 56.720 61.645 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.445 56.310 61.645 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 60.410 61.240 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 60.000 61.240 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 59.590 61.240 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 59.180 61.240 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 58.770 61.240 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 58.360 61.240 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 57.950 61.240 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 57.540 61.240 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 57.130 61.240 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 56.720 61.240 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.040 56.310 61.240 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 60.410 60.835 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 60.000 60.835 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 59.590 60.835 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 59.180 60.835 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 58.770 60.835 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 58.360 60.835 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 57.950 60.835 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 57.540 60.835 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 57.130 60.835 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 56.720 60.835 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.635 56.310 60.835 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 60.410 60.430 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 60.000 60.430 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 59.590 60.430 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 59.180 60.430 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 58.770 60.430 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 58.360 60.430 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 57.950 60.430 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 57.540 60.430 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 57.130 60.430 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 56.720 60.430 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.230 56.310 60.430 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 60.410 60.025 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 60.000 60.025 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 59.590 60.025 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 59.180 60.025 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 58.770 60.025 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 58.360 60.025 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 57.950 60.025 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 57.540 60.025 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 57.130 60.025 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 56.720 60.025 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.825 56.310 60.025 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 60.410 59.620 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 60.000 59.620 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 59.590 59.620 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 59.180 59.620 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 58.770 59.620 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 58.360 59.620 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 57.950 59.620 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 57.540 59.620 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 57.130 59.620 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 56.720 59.620 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.420 56.310 59.620 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 60.410 59.215 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 60.000 59.215 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 59.590 59.215 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 59.180 59.215 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 58.770 59.215 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 58.360 59.215 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 57.950 59.215 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 57.540 59.215 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 57.130 59.215 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 56.720 59.215 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.015 56.310 59.215 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 60.410 58.810 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 60.000 58.810 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 59.590 58.810 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 59.180 58.810 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 58.770 58.810 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 58.360 58.810 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 57.950 58.810 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 57.540 58.810 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 57.130 58.810 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 56.720 58.810 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.610 56.310 58.810 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 60.410 58.405 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 60.000 58.405 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 59.590 58.405 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 59.180 58.405 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 58.770 58.405 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 58.360 58.405 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 57.950 58.405 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 57.540 58.405 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 57.130 58.405 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 56.720 58.405 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.205 56.310 58.405 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 60.410 58.000 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 60.000 58.000 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 59.590 58.000 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 59.180 58.000 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 58.770 58.000 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 58.360 58.000 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 57.950 58.000 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 57.540 58.000 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 57.130 58.000 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 56.720 58.000 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.800 56.310 58.000 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 60.410 57.595 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 60.000 57.595 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 59.590 57.595 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 59.180 57.595 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 58.770 57.595 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 58.360 57.595 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 57.950 57.595 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 57.540 57.595 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 57.130 57.595 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 56.720 57.595 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.395 56.310 57.595 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 60.410 57.190 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 60.000 57.190 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 59.590 57.190 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 59.180 57.190 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 58.770 57.190 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 58.360 57.190 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 57.950 57.190 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 57.540 57.190 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 57.130 57.190 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 56.720 57.190 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.990 56.310 57.190 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 60.410 56.785 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 60.000 56.785 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 59.590 56.785 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 59.180 56.785 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 58.770 56.785 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 58.360 56.785 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 57.950 56.785 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 57.540 56.785 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 57.130 56.785 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 56.720 56.785 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.585 56.310 56.785 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 60.410 56.375 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 60.000 56.375 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 59.590 56.375 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 59.180 56.375 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 58.770 56.375 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 58.360 56.375 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 57.950 56.375 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 57.540 56.375 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 57.130 56.375 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 56.720 56.375 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.175 56.310 56.375 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 60.410 55.965 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 60.000 55.965 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 59.590 55.965 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 59.180 55.965 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 58.770 55.965 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 58.360 55.965 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 57.950 55.965 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 57.540 55.965 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 57.130 55.965 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 56.720 55.965 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.765 56.310 55.965 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 60.410 55.555 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 60.000 55.555 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 59.590 55.555 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 59.180 55.555 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 58.770 55.555 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 58.360 55.555 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 57.950 55.555 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 57.540 55.555 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 57.130 55.555 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 56.720 55.555 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.355 56.310 55.555 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 60.410 55.145 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 60.000 55.145 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 59.590 55.145 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 59.180 55.145 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 58.770 55.145 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 58.360 55.145 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 57.950 55.145 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 57.540 55.145 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 57.130 55.145 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 56.720 55.145 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.945 56.310 55.145 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 60.410 54.735 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 60.000 54.735 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 59.590 54.735 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 59.180 54.735 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 58.770 54.735 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 58.360 54.735 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 57.950 54.735 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 57.540 54.735 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 57.130 54.735 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 56.720 54.735 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.535 56.310 54.735 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 60.410 54.325 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 60.000 54.325 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 59.590 54.325 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 59.180 54.325 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 58.770 54.325 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 58.360 54.325 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 57.950 54.325 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 57.540 54.325 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 57.130 54.325 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 56.720 54.325 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.125 56.310 54.325 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 60.410 53.915 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 60.000 53.915 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 59.590 53.915 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 59.180 53.915 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 58.770 53.915 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 58.360 53.915 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 57.950 53.915 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 57.540 53.915 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 57.130 53.915 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 56.720 53.915 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.715 56.310 53.915 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 60.410 53.505 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 60.000 53.505 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 59.590 53.505 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 59.180 53.505 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 58.770 53.505 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 58.360 53.505 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 57.950 53.505 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 57.540 53.505 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 57.130 53.505 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 56.720 53.505 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.305 56.310 53.505 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 60.410 53.095 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 60.000 53.095 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 59.590 53.095 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 59.180 53.095 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 58.770 53.095 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 58.360 53.095 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 57.950 53.095 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 57.540 53.095 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 57.130 53.095 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 56.720 53.095 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.895 56.310 53.095 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 60.410 52.685 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 60.000 52.685 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 59.590 52.685 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 59.180 52.685 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 58.770 52.685 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 58.360 52.685 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 57.950 52.685 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 57.540 52.685 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 57.130 52.685 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 56.720 52.685 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.485 56.310 52.685 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 60.410 52.275 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 60.000 52.275 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 59.590 52.275 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 59.180 52.275 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 58.770 52.275 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 58.360 52.275 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 57.950 52.275 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 57.540 52.275 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 57.130 52.275 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 56.720 52.275 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.075 56.310 52.275 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 60.410 51.865 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 60.000 51.865 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 59.590 51.865 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 59.180 51.865 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 58.770 51.865 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 58.360 51.865 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 57.950 51.865 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 57.540 51.865 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 57.130 51.865 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 56.720 51.865 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.665 56.310 51.865 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 60.410 51.455 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 60.000 51.455 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 59.590 51.455 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 59.180 51.455 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 58.770 51.455 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 58.360 51.455 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 57.950 51.455 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 57.540 51.455 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 57.130 51.455 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 56.720 51.455 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.255 56.310 51.455 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 60.410 51.045 60.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 60.000 51.045 60.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 59.590 51.045 59.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 59.180 51.045 59.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 58.770 51.045 58.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 58.360 51.045 58.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 57.950 51.045 58.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 57.540 51.045 57.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 57.130 51.045 57.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 56.720 51.045 56.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.845 56.310 51.045 56.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 60.350 24.370 60.670 ;
      LAYER met4 ;
        RECT 24.050 60.350 24.370 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 59.940 24.370 60.260 ;
      LAYER met4 ;
        RECT 24.050 59.940 24.370 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 59.530 24.370 59.850 ;
      LAYER met4 ;
        RECT 24.050 59.530 24.370 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 59.120 24.370 59.440 ;
      LAYER met4 ;
        RECT 24.050 59.120 24.370 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 58.710 24.370 59.030 ;
      LAYER met4 ;
        RECT 24.050 58.710 24.370 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 58.300 24.370 58.620 ;
      LAYER met4 ;
        RECT 24.050 58.300 24.370 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 57.890 24.370 58.210 ;
      LAYER met4 ;
        RECT 24.050 57.890 24.370 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 57.480 24.370 57.800 ;
      LAYER met4 ;
        RECT 24.050 57.480 24.370 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 57.070 24.370 57.390 ;
      LAYER met4 ;
        RECT 24.050 57.070 24.370 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 56.660 24.370 56.980 ;
      LAYER met4 ;
        RECT 24.050 56.660 24.370 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.050 56.250 24.370 56.570 ;
      LAYER met4 ;
        RECT 24.050 56.250 24.370 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 60.350 23.965 60.670 ;
      LAYER met4 ;
        RECT 23.645 60.350 23.965 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 59.940 23.965 60.260 ;
      LAYER met4 ;
        RECT 23.645 59.940 23.965 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 59.530 23.965 59.850 ;
      LAYER met4 ;
        RECT 23.645 59.530 23.965 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 59.120 23.965 59.440 ;
      LAYER met4 ;
        RECT 23.645 59.120 23.965 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 58.710 23.965 59.030 ;
      LAYER met4 ;
        RECT 23.645 58.710 23.965 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 58.300 23.965 58.620 ;
      LAYER met4 ;
        RECT 23.645 58.300 23.965 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 57.890 23.965 58.210 ;
      LAYER met4 ;
        RECT 23.645 57.890 23.965 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 57.480 23.965 57.800 ;
      LAYER met4 ;
        RECT 23.645 57.480 23.965 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 57.070 23.965 57.390 ;
      LAYER met4 ;
        RECT 23.645 57.070 23.965 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 56.660 23.965 56.980 ;
      LAYER met4 ;
        RECT 23.645 56.660 23.965 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.645 56.250 23.965 56.570 ;
      LAYER met4 ;
        RECT 23.645 56.250 23.965 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 60.350 23.560 60.670 ;
      LAYER met4 ;
        RECT 23.240 60.350 23.560 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 59.940 23.560 60.260 ;
      LAYER met4 ;
        RECT 23.240 59.940 23.560 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 59.530 23.560 59.850 ;
      LAYER met4 ;
        RECT 23.240 59.530 23.560 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 59.120 23.560 59.440 ;
      LAYER met4 ;
        RECT 23.240 59.120 23.560 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 58.710 23.560 59.030 ;
      LAYER met4 ;
        RECT 23.240 58.710 23.560 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 58.300 23.560 58.620 ;
      LAYER met4 ;
        RECT 23.240 58.300 23.560 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 57.890 23.560 58.210 ;
      LAYER met4 ;
        RECT 23.240 57.890 23.560 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 57.480 23.560 57.800 ;
      LAYER met4 ;
        RECT 23.240 57.480 23.560 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 57.070 23.560 57.390 ;
      LAYER met4 ;
        RECT 23.240 57.070 23.560 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 56.660 23.560 56.980 ;
      LAYER met4 ;
        RECT 23.240 56.660 23.560 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.240 56.250 23.560 56.570 ;
      LAYER met4 ;
        RECT 23.240 56.250 23.560 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 60.350 23.155 60.670 ;
      LAYER met4 ;
        RECT 22.835 60.350 23.155 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 59.940 23.155 60.260 ;
      LAYER met4 ;
        RECT 22.835 59.940 23.155 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 59.530 23.155 59.850 ;
      LAYER met4 ;
        RECT 22.835 59.530 23.155 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 59.120 23.155 59.440 ;
      LAYER met4 ;
        RECT 22.835 59.120 23.155 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 58.710 23.155 59.030 ;
      LAYER met4 ;
        RECT 22.835 58.710 23.155 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 58.300 23.155 58.620 ;
      LAYER met4 ;
        RECT 22.835 58.300 23.155 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 57.890 23.155 58.210 ;
      LAYER met4 ;
        RECT 22.835 57.890 23.155 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 57.480 23.155 57.800 ;
      LAYER met4 ;
        RECT 22.835 57.480 23.155 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 57.070 23.155 57.390 ;
      LAYER met4 ;
        RECT 22.835 57.070 23.155 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 56.660 23.155 56.980 ;
      LAYER met4 ;
        RECT 22.835 56.660 23.155 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.835 56.250 23.155 56.570 ;
      LAYER met4 ;
        RECT 22.835 56.250 23.155 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 60.350 22.750 60.670 ;
      LAYER met4 ;
        RECT 22.430 60.350 22.750 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 59.940 22.750 60.260 ;
      LAYER met4 ;
        RECT 22.430 59.940 22.750 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 59.530 22.750 59.850 ;
      LAYER met4 ;
        RECT 22.430 59.530 22.750 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 59.120 22.750 59.440 ;
      LAYER met4 ;
        RECT 22.430 59.120 22.750 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 58.710 22.750 59.030 ;
      LAYER met4 ;
        RECT 22.430 58.710 22.750 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 58.300 22.750 58.620 ;
      LAYER met4 ;
        RECT 22.430 58.300 22.750 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 57.890 22.750 58.210 ;
      LAYER met4 ;
        RECT 22.430 57.890 22.750 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 57.480 22.750 57.800 ;
      LAYER met4 ;
        RECT 22.430 57.480 22.750 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 57.070 22.750 57.390 ;
      LAYER met4 ;
        RECT 22.430 57.070 22.750 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 56.660 22.750 56.980 ;
      LAYER met4 ;
        RECT 22.430 56.660 22.750 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.430 56.250 22.750 56.570 ;
      LAYER met4 ;
        RECT 22.430 56.250 22.750 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 60.350 22.345 60.670 ;
      LAYER met4 ;
        RECT 22.025 60.350 22.345 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 59.940 22.345 60.260 ;
      LAYER met4 ;
        RECT 22.025 59.940 22.345 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 59.530 22.345 59.850 ;
      LAYER met4 ;
        RECT 22.025 59.530 22.345 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 59.120 22.345 59.440 ;
      LAYER met4 ;
        RECT 22.025 59.120 22.345 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 58.710 22.345 59.030 ;
      LAYER met4 ;
        RECT 22.025 58.710 22.345 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 58.300 22.345 58.620 ;
      LAYER met4 ;
        RECT 22.025 58.300 22.345 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 57.890 22.345 58.210 ;
      LAYER met4 ;
        RECT 22.025 57.890 22.345 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 57.480 22.345 57.800 ;
      LAYER met4 ;
        RECT 22.025 57.480 22.345 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 57.070 22.345 57.390 ;
      LAYER met4 ;
        RECT 22.025 57.070 22.345 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 56.660 22.345 56.980 ;
      LAYER met4 ;
        RECT 22.025 56.660 22.345 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.025 56.250 22.345 56.570 ;
      LAYER met4 ;
        RECT 22.025 56.250 22.345 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 60.350 21.940 60.670 ;
      LAYER met4 ;
        RECT 21.620 60.350 21.940 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 59.940 21.940 60.260 ;
      LAYER met4 ;
        RECT 21.620 59.940 21.940 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 59.530 21.940 59.850 ;
      LAYER met4 ;
        RECT 21.620 59.530 21.940 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 59.120 21.940 59.440 ;
      LAYER met4 ;
        RECT 21.620 59.120 21.940 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 58.710 21.940 59.030 ;
      LAYER met4 ;
        RECT 21.620 58.710 21.940 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 58.300 21.940 58.620 ;
      LAYER met4 ;
        RECT 21.620 58.300 21.940 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 57.890 21.940 58.210 ;
      LAYER met4 ;
        RECT 21.620 57.890 21.940 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 57.480 21.940 57.800 ;
      LAYER met4 ;
        RECT 21.620 57.480 21.940 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 57.070 21.940 57.390 ;
      LAYER met4 ;
        RECT 21.620 57.070 21.940 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 56.660 21.940 56.980 ;
      LAYER met4 ;
        RECT 21.620 56.660 21.940 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.620 56.250 21.940 56.570 ;
      LAYER met4 ;
        RECT 21.620 56.250 21.940 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 60.350 21.535 60.670 ;
      LAYER met4 ;
        RECT 21.215 60.350 21.535 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 59.940 21.535 60.260 ;
      LAYER met4 ;
        RECT 21.215 59.940 21.535 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 59.530 21.535 59.850 ;
      LAYER met4 ;
        RECT 21.215 59.530 21.535 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 59.120 21.535 59.440 ;
      LAYER met4 ;
        RECT 21.215 59.120 21.535 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 58.710 21.535 59.030 ;
      LAYER met4 ;
        RECT 21.215 58.710 21.535 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 58.300 21.535 58.620 ;
      LAYER met4 ;
        RECT 21.215 58.300 21.535 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 57.890 21.535 58.210 ;
      LAYER met4 ;
        RECT 21.215 57.890 21.535 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 57.480 21.535 57.800 ;
      LAYER met4 ;
        RECT 21.215 57.480 21.535 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 57.070 21.535 57.390 ;
      LAYER met4 ;
        RECT 21.215 57.070 21.535 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 56.660 21.535 56.980 ;
      LAYER met4 ;
        RECT 21.215 56.660 21.535 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.215 56.250 21.535 56.570 ;
      LAYER met4 ;
        RECT 21.215 56.250 21.535 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 60.350 21.130 60.670 ;
      LAYER met4 ;
        RECT 20.810 60.350 21.130 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 59.940 21.130 60.260 ;
      LAYER met4 ;
        RECT 20.810 59.940 21.130 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 59.530 21.130 59.850 ;
      LAYER met4 ;
        RECT 20.810 59.530 21.130 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 59.120 21.130 59.440 ;
      LAYER met4 ;
        RECT 20.810 59.120 21.130 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 58.710 21.130 59.030 ;
      LAYER met4 ;
        RECT 20.810 58.710 21.130 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 58.300 21.130 58.620 ;
      LAYER met4 ;
        RECT 20.810 58.300 21.130 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 57.890 21.130 58.210 ;
      LAYER met4 ;
        RECT 20.810 57.890 21.130 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 57.480 21.130 57.800 ;
      LAYER met4 ;
        RECT 20.810 57.480 21.130 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 57.070 21.130 57.390 ;
      LAYER met4 ;
        RECT 20.810 57.070 21.130 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 56.660 21.130 56.980 ;
      LAYER met4 ;
        RECT 20.810 56.660 21.130 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.810 56.250 21.130 56.570 ;
      LAYER met4 ;
        RECT 20.810 56.250 21.130 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 60.350 20.725 60.670 ;
      LAYER met4 ;
        RECT 20.405 60.350 20.725 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 59.940 20.725 60.260 ;
      LAYER met4 ;
        RECT 20.405 59.940 20.725 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 59.530 20.725 59.850 ;
      LAYER met4 ;
        RECT 20.405 59.530 20.725 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 59.120 20.725 59.440 ;
      LAYER met4 ;
        RECT 20.405 59.120 20.725 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 58.710 20.725 59.030 ;
      LAYER met4 ;
        RECT 20.405 58.710 20.725 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 58.300 20.725 58.620 ;
      LAYER met4 ;
        RECT 20.405 58.300 20.725 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 57.890 20.725 58.210 ;
      LAYER met4 ;
        RECT 20.405 57.890 20.725 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 57.480 20.725 57.800 ;
      LAYER met4 ;
        RECT 20.405 57.480 20.725 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 57.070 20.725 57.390 ;
      LAYER met4 ;
        RECT 20.405 57.070 20.725 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 56.660 20.725 56.980 ;
      LAYER met4 ;
        RECT 20.405 56.660 20.725 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.405 56.250 20.725 56.570 ;
      LAYER met4 ;
        RECT 20.405 56.250 20.725 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 60.350 20.320 60.670 ;
      LAYER met4 ;
        RECT 20.000 60.350 20.320 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 59.940 20.320 60.260 ;
      LAYER met4 ;
        RECT 20.000 59.940 20.320 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 59.530 20.320 59.850 ;
      LAYER met4 ;
        RECT 20.000 59.530 20.320 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 59.120 20.320 59.440 ;
      LAYER met4 ;
        RECT 20.000 59.120 20.320 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 58.710 20.320 59.030 ;
      LAYER met4 ;
        RECT 20.000 58.710 20.320 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 58.300 20.320 58.620 ;
      LAYER met4 ;
        RECT 20.000 58.300 20.320 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 57.890 20.320 58.210 ;
      LAYER met4 ;
        RECT 20.000 57.890 20.320 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 57.480 20.320 57.800 ;
      LAYER met4 ;
        RECT 20.000 57.480 20.320 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 57.070 20.320 57.390 ;
      LAYER met4 ;
        RECT 20.000 57.070 20.320 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 56.660 20.320 56.980 ;
      LAYER met4 ;
        RECT 20.000 56.660 20.320 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.000 56.250 20.320 56.570 ;
      LAYER met4 ;
        RECT 20.000 56.250 20.320 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 60.350 19.915 60.670 ;
      LAYER met4 ;
        RECT 19.595 60.350 19.915 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 59.940 19.915 60.260 ;
      LAYER met4 ;
        RECT 19.595 59.940 19.915 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 59.530 19.915 59.850 ;
      LAYER met4 ;
        RECT 19.595 59.530 19.915 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 59.120 19.915 59.440 ;
      LAYER met4 ;
        RECT 19.595 59.120 19.915 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 58.710 19.915 59.030 ;
      LAYER met4 ;
        RECT 19.595 58.710 19.915 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 58.300 19.915 58.620 ;
      LAYER met4 ;
        RECT 19.595 58.300 19.915 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 57.890 19.915 58.210 ;
      LAYER met4 ;
        RECT 19.595 57.890 19.915 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 57.480 19.915 57.800 ;
      LAYER met4 ;
        RECT 19.595 57.480 19.915 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 57.070 19.915 57.390 ;
      LAYER met4 ;
        RECT 19.595 57.070 19.915 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 56.660 19.915 56.980 ;
      LAYER met4 ;
        RECT 19.595 56.660 19.915 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.595 56.250 19.915 56.570 ;
      LAYER met4 ;
        RECT 19.595 56.250 19.915 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 60.350 19.510 60.670 ;
      LAYER met4 ;
        RECT 19.190 60.350 19.510 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 59.940 19.510 60.260 ;
      LAYER met4 ;
        RECT 19.190 59.940 19.510 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 59.530 19.510 59.850 ;
      LAYER met4 ;
        RECT 19.190 59.530 19.510 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 59.120 19.510 59.440 ;
      LAYER met4 ;
        RECT 19.190 59.120 19.510 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 58.710 19.510 59.030 ;
      LAYER met4 ;
        RECT 19.190 58.710 19.510 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 58.300 19.510 58.620 ;
      LAYER met4 ;
        RECT 19.190 58.300 19.510 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 57.890 19.510 58.210 ;
      LAYER met4 ;
        RECT 19.190 57.890 19.510 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 57.480 19.510 57.800 ;
      LAYER met4 ;
        RECT 19.190 57.480 19.510 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 57.070 19.510 57.390 ;
      LAYER met4 ;
        RECT 19.190 57.070 19.510 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 56.660 19.510 56.980 ;
      LAYER met4 ;
        RECT 19.190 56.660 19.510 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.190 56.250 19.510 56.570 ;
      LAYER met4 ;
        RECT 19.190 56.250 19.510 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 60.350 19.105 60.670 ;
      LAYER met4 ;
        RECT 18.785 60.350 19.105 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 59.940 19.105 60.260 ;
      LAYER met4 ;
        RECT 18.785 59.940 19.105 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 59.530 19.105 59.850 ;
      LAYER met4 ;
        RECT 18.785 59.530 19.105 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 59.120 19.105 59.440 ;
      LAYER met4 ;
        RECT 18.785 59.120 19.105 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 58.710 19.105 59.030 ;
      LAYER met4 ;
        RECT 18.785 58.710 19.105 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 58.300 19.105 58.620 ;
      LAYER met4 ;
        RECT 18.785 58.300 19.105 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 57.890 19.105 58.210 ;
      LAYER met4 ;
        RECT 18.785 57.890 19.105 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 57.480 19.105 57.800 ;
      LAYER met4 ;
        RECT 18.785 57.480 19.105 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 57.070 19.105 57.390 ;
      LAYER met4 ;
        RECT 18.785 57.070 19.105 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 56.660 19.105 56.980 ;
      LAYER met4 ;
        RECT 18.785 56.660 19.105 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.785 56.250 19.105 56.570 ;
      LAYER met4 ;
        RECT 18.785 56.250 19.105 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 60.350 18.700 60.670 ;
      LAYER met4 ;
        RECT 18.380 60.350 18.700 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 59.940 18.700 60.260 ;
      LAYER met4 ;
        RECT 18.380 59.940 18.700 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 59.530 18.700 59.850 ;
      LAYER met4 ;
        RECT 18.380 59.530 18.700 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 59.120 18.700 59.440 ;
      LAYER met4 ;
        RECT 18.380 59.120 18.700 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 58.710 18.700 59.030 ;
      LAYER met4 ;
        RECT 18.380 58.710 18.700 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 58.300 18.700 58.620 ;
      LAYER met4 ;
        RECT 18.380 58.300 18.700 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 57.890 18.700 58.210 ;
      LAYER met4 ;
        RECT 18.380 57.890 18.700 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 57.480 18.700 57.800 ;
      LAYER met4 ;
        RECT 18.380 57.480 18.700 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 57.070 18.700 57.390 ;
      LAYER met4 ;
        RECT 18.380 57.070 18.700 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 56.660 18.700 56.980 ;
      LAYER met4 ;
        RECT 18.380 56.660 18.700 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.380 56.250 18.700 56.570 ;
      LAYER met4 ;
        RECT 18.380 56.250 18.700 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 60.350 18.295 60.670 ;
      LAYER met4 ;
        RECT 17.975 60.350 18.295 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 59.940 18.295 60.260 ;
      LAYER met4 ;
        RECT 17.975 59.940 18.295 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 59.530 18.295 59.850 ;
      LAYER met4 ;
        RECT 17.975 59.530 18.295 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 59.120 18.295 59.440 ;
      LAYER met4 ;
        RECT 17.975 59.120 18.295 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 58.710 18.295 59.030 ;
      LAYER met4 ;
        RECT 17.975 58.710 18.295 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 58.300 18.295 58.620 ;
      LAYER met4 ;
        RECT 17.975 58.300 18.295 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 57.890 18.295 58.210 ;
      LAYER met4 ;
        RECT 17.975 57.890 18.295 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 57.480 18.295 57.800 ;
      LAYER met4 ;
        RECT 17.975 57.480 18.295 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 57.070 18.295 57.390 ;
      LAYER met4 ;
        RECT 17.975 57.070 18.295 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 56.660 18.295 56.980 ;
      LAYER met4 ;
        RECT 17.975 56.660 18.295 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.975 56.250 18.295 56.570 ;
      LAYER met4 ;
        RECT 17.975 56.250 18.295 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 60.350 17.890 60.670 ;
      LAYER met4 ;
        RECT 17.570 60.350 17.890 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 59.940 17.890 60.260 ;
      LAYER met4 ;
        RECT 17.570 59.940 17.890 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 59.530 17.890 59.850 ;
      LAYER met4 ;
        RECT 17.570 59.530 17.890 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 59.120 17.890 59.440 ;
      LAYER met4 ;
        RECT 17.570 59.120 17.890 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 58.710 17.890 59.030 ;
      LAYER met4 ;
        RECT 17.570 58.710 17.890 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 58.300 17.890 58.620 ;
      LAYER met4 ;
        RECT 17.570 58.300 17.890 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 57.890 17.890 58.210 ;
      LAYER met4 ;
        RECT 17.570 57.890 17.890 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 57.480 17.890 57.800 ;
      LAYER met4 ;
        RECT 17.570 57.480 17.890 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 57.070 17.890 57.390 ;
      LAYER met4 ;
        RECT 17.570 57.070 17.890 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 56.660 17.890 56.980 ;
      LAYER met4 ;
        RECT 17.570 56.660 17.890 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.570 56.250 17.890 56.570 ;
      LAYER met4 ;
        RECT 17.570 56.250 17.890 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 60.350 17.485 60.670 ;
      LAYER met4 ;
        RECT 17.165 60.350 17.485 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 59.940 17.485 60.260 ;
      LAYER met4 ;
        RECT 17.165 59.940 17.485 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 59.530 17.485 59.850 ;
      LAYER met4 ;
        RECT 17.165 59.530 17.485 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 59.120 17.485 59.440 ;
      LAYER met4 ;
        RECT 17.165 59.120 17.485 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 58.710 17.485 59.030 ;
      LAYER met4 ;
        RECT 17.165 58.710 17.485 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 58.300 17.485 58.620 ;
      LAYER met4 ;
        RECT 17.165 58.300 17.485 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 57.890 17.485 58.210 ;
      LAYER met4 ;
        RECT 17.165 57.890 17.485 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 57.480 17.485 57.800 ;
      LAYER met4 ;
        RECT 17.165 57.480 17.485 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 57.070 17.485 57.390 ;
      LAYER met4 ;
        RECT 17.165 57.070 17.485 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 56.660 17.485 56.980 ;
      LAYER met4 ;
        RECT 17.165 56.660 17.485 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.165 56.250 17.485 56.570 ;
      LAYER met4 ;
        RECT 17.165 56.250 17.485 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 60.350 17.080 60.670 ;
      LAYER met4 ;
        RECT 16.760 60.350 17.080 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 59.940 17.080 60.260 ;
      LAYER met4 ;
        RECT 16.760 59.940 17.080 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 59.530 17.080 59.850 ;
      LAYER met4 ;
        RECT 16.760 59.530 17.080 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 59.120 17.080 59.440 ;
      LAYER met4 ;
        RECT 16.760 59.120 17.080 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 58.710 17.080 59.030 ;
      LAYER met4 ;
        RECT 16.760 58.710 17.080 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 58.300 17.080 58.620 ;
      LAYER met4 ;
        RECT 16.760 58.300 17.080 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 57.890 17.080 58.210 ;
      LAYER met4 ;
        RECT 16.760 57.890 17.080 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 57.480 17.080 57.800 ;
      LAYER met4 ;
        RECT 16.760 57.480 17.080 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 57.070 17.080 57.390 ;
      LAYER met4 ;
        RECT 16.760 57.070 17.080 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 56.660 17.080 56.980 ;
      LAYER met4 ;
        RECT 16.760 56.660 17.080 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.760 56.250 17.080 56.570 ;
      LAYER met4 ;
        RECT 16.760 56.250 17.080 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 60.350 16.675 60.670 ;
      LAYER met4 ;
        RECT 16.355 60.350 16.675 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 59.940 16.675 60.260 ;
      LAYER met4 ;
        RECT 16.355 59.940 16.675 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 59.530 16.675 59.850 ;
      LAYER met4 ;
        RECT 16.355 59.530 16.675 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 59.120 16.675 59.440 ;
      LAYER met4 ;
        RECT 16.355 59.120 16.675 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 58.710 16.675 59.030 ;
      LAYER met4 ;
        RECT 16.355 58.710 16.675 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 58.300 16.675 58.620 ;
      LAYER met4 ;
        RECT 16.355 58.300 16.675 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 57.890 16.675 58.210 ;
      LAYER met4 ;
        RECT 16.355 57.890 16.675 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 57.480 16.675 57.800 ;
      LAYER met4 ;
        RECT 16.355 57.480 16.675 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 57.070 16.675 57.390 ;
      LAYER met4 ;
        RECT 16.355 57.070 16.675 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 56.660 16.675 56.980 ;
      LAYER met4 ;
        RECT 16.355 56.660 16.675 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.355 56.250 16.675 56.570 ;
      LAYER met4 ;
        RECT 16.355 56.250 16.675 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 60.350 16.270 60.670 ;
      LAYER met4 ;
        RECT 15.950 60.350 16.270 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 59.940 16.270 60.260 ;
      LAYER met4 ;
        RECT 15.950 59.940 16.270 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 59.530 16.270 59.850 ;
      LAYER met4 ;
        RECT 15.950 59.530 16.270 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 59.120 16.270 59.440 ;
      LAYER met4 ;
        RECT 15.950 59.120 16.270 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 58.710 16.270 59.030 ;
      LAYER met4 ;
        RECT 15.950 58.710 16.270 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 58.300 16.270 58.620 ;
      LAYER met4 ;
        RECT 15.950 58.300 16.270 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 57.890 16.270 58.210 ;
      LAYER met4 ;
        RECT 15.950 57.890 16.270 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 57.480 16.270 57.800 ;
      LAYER met4 ;
        RECT 15.950 57.480 16.270 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 57.070 16.270 57.390 ;
      LAYER met4 ;
        RECT 15.950 57.070 16.270 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 56.660 16.270 56.980 ;
      LAYER met4 ;
        RECT 15.950 56.660 16.270 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.950 56.250 16.270 56.570 ;
      LAYER met4 ;
        RECT 15.950 56.250 16.270 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 60.350 15.865 60.670 ;
      LAYER met4 ;
        RECT 15.545 60.350 15.865 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 59.940 15.865 60.260 ;
      LAYER met4 ;
        RECT 15.545 59.940 15.865 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 59.530 15.865 59.850 ;
      LAYER met4 ;
        RECT 15.545 59.530 15.865 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 59.120 15.865 59.440 ;
      LAYER met4 ;
        RECT 15.545 59.120 15.865 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 58.710 15.865 59.030 ;
      LAYER met4 ;
        RECT 15.545 58.710 15.865 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 58.300 15.865 58.620 ;
      LAYER met4 ;
        RECT 15.545 58.300 15.865 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 57.890 15.865 58.210 ;
      LAYER met4 ;
        RECT 15.545 57.890 15.865 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 57.480 15.865 57.800 ;
      LAYER met4 ;
        RECT 15.545 57.480 15.865 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 57.070 15.865 57.390 ;
      LAYER met4 ;
        RECT 15.545 57.070 15.865 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 56.660 15.865 56.980 ;
      LAYER met4 ;
        RECT 15.545 56.660 15.865 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.545 56.250 15.865 56.570 ;
      LAYER met4 ;
        RECT 15.545 56.250 15.865 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 60.350 15.460 60.670 ;
      LAYER met4 ;
        RECT 15.140 60.350 15.460 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 59.940 15.460 60.260 ;
      LAYER met4 ;
        RECT 15.140 59.940 15.460 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 59.530 15.460 59.850 ;
      LAYER met4 ;
        RECT 15.140 59.530 15.460 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 59.120 15.460 59.440 ;
      LAYER met4 ;
        RECT 15.140 59.120 15.460 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 58.710 15.460 59.030 ;
      LAYER met4 ;
        RECT 15.140 58.710 15.460 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 58.300 15.460 58.620 ;
      LAYER met4 ;
        RECT 15.140 58.300 15.460 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 57.890 15.460 58.210 ;
      LAYER met4 ;
        RECT 15.140 57.890 15.460 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 57.480 15.460 57.800 ;
      LAYER met4 ;
        RECT 15.140 57.480 15.460 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 57.070 15.460 57.390 ;
      LAYER met4 ;
        RECT 15.140 57.070 15.460 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 56.660 15.460 56.980 ;
      LAYER met4 ;
        RECT 15.140 56.660 15.460 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.140 56.250 15.460 56.570 ;
      LAYER met4 ;
        RECT 15.140 56.250 15.460 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 60.350 15.055 60.670 ;
      LAYER met4 ;
        RECT 14.735 60.350 15.055 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 59.940 15.055 60.260 ;
      LAYER met4 ;
        RECT 14.735 59.940 15.055 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 59.530 15.055 59.850 ;
      LAYER met4 ;
        RECT 14.735 59.530 15.055 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 59.120 15.055 59.440 ;
      LAYER met4 ;
        RECT 14.735 59.120 15.055 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 58.710 15.055 59.030 ;
      LAYER met4 ;
        RECT 14.735 58.710 15.055 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 58.300 15.055 58.620 ;
      LAYER met4 ;
        RECT 14.735 58.300 15.055 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 57.890 15.055 58.210 ;
      LAYER met4 ;
        RECT 14.735 57.890 15.055 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 57.480 15.055 57.800 ;
      LAYER met4 ;
        RECT 14.735 57.480 15.055 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 57.070 15.055 57.390 ;
      LAYER met4 ;
        RECT 14.735 57.070 15.055 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 56.660 15.055 56.980 ;
      LAYER met4 ;
        RECT 14.735 56.660 15.055 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.735 56.250 15.055 56.570 ;
      LAYER met4 ;
        RECT 14.735 56.250 15.055 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 60.350 14.650 60.670 ;
      LAYER met4 ;
        RECT 14.330 60.350 14.650 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 59.940 14.650 60.260 ;
      LAYER met4 ;
        RECT 14.330 59.940 14.650 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 59.530 14.650 59.850 ;
      LAYER met4 ;
        RECT 14.330 59.530 14.650 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 59.120 14.650 59.440 ;
      LAYER met4 ;
        RECT 14.330 59.120 14.650 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 58.710 14.650 59.030 ;
      LAYER met4 ;
        RECT 14.330 58.710 14.650 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 58.300 14.650 58.620 ;
      LAYER met4 ;
        RECT 14.330 58.300 14.650 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 57.890 14.650 58.210 ;
      LAYER met4 ;
        RECT 14.330 57.890 14.650 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 57.480 14.650 57.800 ;
      LAYER met4 ;
        RECT 14.330 57.480 14.650 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 57.070 14.650 57.390 ;
      LAYER met4 ;
        RECT 14.330 57.070 14.650 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 56.660 14.650 56.980 ;
      LAYER met4 ;
        RECT 14.330 56.660 14.650 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.330 56.250 14.650 56.570 ;
      LAYER met4 ;
        RECT 14.330 56.250 14.650 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 60.350 14.245 60.670 ;
      LAYER met4 ;
        RECT 13.925 60.350 14.245 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 59.940 14.245 60.260 ;
      LAYER met4 ;
        RECT 13.925 59.940 14.245 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 59.530 14.245 59.850 ;
      LAYER met4 ;
        RECT 13.925 59.530 14.245 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 59.120 14.245 59.440 ;
      LAYER met4 ;
        RECT 13.925 59.120 14.245 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 58.710 14.245 59.030 ;
      LAYER met4 ;
        RECT 13.925 58.710 14.245 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 58.300 14.245 58.620 ;
      LAYER met4 ;
        RECT 13.925 58.300 14.245 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 57.890 14.245 58.210 ;
      LAYER met4 ;
        RECT 13.925 57.890 14.245 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 57.480 14.245 57.800 ;
      LAYER met4 ;
        RECT 13.925 57.480 14.245 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 57.070 14.245 57.390 ;
      LAYER met4 ;
        RECT 13.925 57.070 14.245 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 56.660 14.245 56.980 ;
      LAYER met4 ;
        RECT 13.925 56.660 14.245 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.925 56.250 14.245 56.570 ;
      LAYER met4 ;
        RECT 13.925 56.250 14.245 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 60.350 13.840 60.670 ;
      LAYER met4 ;
        RECT 13.520 60.350 13.840 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 59.940 13.840 60.260 ;
      LAYER met4 ;
        RECT 13.520 59.940 13.840 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 59.530 13.840 59.850 ;
      LAYER met4 ;
        RECT 13.520 59.530 13.840 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 59.120 13.840 59.440 ;
      LAYER met4 ;
        RECT 13.520 59.120 13.840 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 58.710 13.840 59.030 ;
      LAYER met4 ;
        RECT 13.520 58.710 13.840 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 58.300 13.840 58.620 ;
      LAYER met4 ;
        RECT 13.520 58.300 13.840 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 57.890 13.840 58.210 ;
      LAYER met4 ;
        RECT 13.520 57.890 13.840 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 57.480 13.840 57.800 ;
      LAYER met4 ;
        RECT 13.520 57.480 13.840 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 57.070 13.840 57.390 ;
      LAYER met4 ;
        RECT 13.520 57.070 13.840 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 56.660 13.840 56.980 ;
      LAYER met4 ;
        RECT 13.520 56.660 13.840 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.520 56.250 13.840 56.570 ;
      LAYER met4 ;
        RECT 13.520 56.250 13.840 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 60.350 13.435 60.670 ;
      LAYER met4 ;
        RECT 13.115 60.350 13.435 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 59.940 13.435 60.260 ;
      LAYER met4 ;
        RECT 13.115 59.940 13.435 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 59.530 13.435 59.850 ;
      LAYER met4 ;
        RECT 13.115 59.530 13.435 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 59.120 13.435 59.440 ;
      LAYER met4 ;
        RECT 13.115 59.120 13.435 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 58.710 13.435 59.030 ;
      LAYER met4 ;
        RECT 13.115 58.710 13.435 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 58.300 13.435 58.620 ;
      LAYER met4 ;
        RECT 13.115 58.300 13.435 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 57.890 13.435 58.210 ;
      LAYER met4 ;
        RECT 13.115 57.890 13.435 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 57.480 13.435 57.800 ;
      LAYER met4 ;
        RECT 13.115 57.480 13.435 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 57.070 13.435 57.390 ;
      LAYER met4 ;
        RECT 13.115 57.070 13.435 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 56.660 13.435 56.980 ;
      LAYER met4 ;
        RECT 13.115 56.660 13.435 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.115 56.250 13.435 56.570 ;
      LAYER met4 ;
        RECT 13.115 56.250 13.435 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 60.350 13.030 60.670 ;
      LAYER met4 ;
        RECT 12.710 60.350 13.030 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 59.940 13.030 60.260 ;
      LAYER met4 ;
        RECT 12.710 59.940 13.030 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 59.530 13.030 59.850 ;
      LAYER met4 ;
        RECT 12.710 59.530 13.030 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 59.120 13.030 59.440 ;
      LAYER met4 ;
        RECT 12.710 59.120 13.030 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 58.710 13.030 59.030 ;
      LAYER met4 ;
        RECT 12.710 58.710 13.030 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 58.300 13.030 58.620 ;
      LAYER met4 ;
        RECT 12.710 58.300 13.030 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 57.890 13.030 58.210 ;
      LAYER met4 ;
        RECT 12.710 57.890 13.030 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 57.480 13.030 57.800 ;
      LAYER met4 ;
        RECT 12.710 57.480 13.030 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 57.070 13.030 57.390 ;
      LAYER met4 ;
        RECT 12.710 57.070 13.030 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 56.660 13.030 56.980 ;
      LAYER met4 ;
        RECT 12.710 56.660 13.030 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.710 56.250 13.030 56.570 ;
      LAYER met4 ;
        RECT 12.710 56.250 13.030 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 60.350 12.625 60.670 ;
      LAYER met4 ;
        RECT 12.305 60.350 12.625 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 59.940 12.625 60.260 ;
      LAYER met4 ;
        RECT 12.305 59.940 12.625 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 59.530 12.625 59.850 ;
      LAYER met4 ;
        RECT 12.305 59.530 12.625 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 59.120 12.625 59.440 ;
      LAYER met4 ;
        RECT 12.305 59.120 12.625 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 58.710 12.625 59.030 ;
      LAYER met4 ;
        RECT 12.305 58.710 12.625 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 58.300 12.625 58.620 ;
      LAYER met4 ;
        RECT 12.305 58.300 12.625 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 57.890 12.625 58.210 ;
      LAYER met4 ;
        RECT 12.305 57.890 12.625 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 57.480 12.625 57.800 ;
      LAYER met4 ;
        RECT 12.305 57.480 12.625 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 57.070 12.625 57.390 ;
      LAYER met4 ;
        RECT 12.305 57.070 12.625 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 56.660 12.625 56.980 ;
      LAYER met4 ;
        RECT 12.305 56.660 12.625 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.305 56.250 12.625 56.570 ;
      LAYER met4 ;
        RECT 12.305 56.250 12.625 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 60.350 12.220 60.670 ;
      LAYER met4 ;
        RECT 11.900 60.350 12.220 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 59.940 12.220 60.260 ;
      LAYER met4 ;
        RECT 11.900 59.940 12.220 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 59.530 12.220 59.850 ;
      LAYER met4 ;
        RECT 11.900 59.530 12.220 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 59.120 12.220 59.440 ;
      LAYER met4 ;
        RECT 11.900 59.120 12.220 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 58.710 12.220 59.030 ;
      LAYER met4 ;
        RECT 11.900 58.710 12.220 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 58.300 12.220 58.620 ;
      LAYER met4 ;
        RECT 11.900 58.300 12.220 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 57.890 12.220 58.210 ;
      LAYER met4 ;
        RECT 11.900 57.890 12.220 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 57.480 12.220 57.800 ;
      LAYER met4 ;
        RECT 11.900 57.480 12.220 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 57.070 12.220 57.390 ;
      LAYER met4 ;
        RECT 11.900 57.070 12.220 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 56.660 12.220 56.980 ;
      LAYER met4 ;
        RECT 11.900 56.660 12.220 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.900 56.250 12.220 56.570 ;
      LAYER met4 ;
        RECT 11.900 56.250 12.220 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 60.350 11.815 60.670 ;
      LAYER met4 ;
        RECT 11.495 60.350 11.815 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 59.940 11.815 60.260 ;
      LAYER met4 ;
        RECT 11.495 59.940 11.815 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 59.530 11.815 59.850 ;
      LAYER met4 ;
        RECT 11.495 59.530 11.815 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 59.120 11.815 59.440 ;
      LAYER met4 ;
        RECT 11.495 59.120 11.815 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 58.710 11.815 59.030 ;
      LAYER met4 ;
        RECT 11.495 58.710 11.815 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 58.300 11.815 58.620 ;
      LAYER met4 ;
        RECT 11.495 58.300 11.815 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 57.890 11.815 58.210 ;
      LAYER met4 ;
        RECT 11.495 57.890 11.815 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 57.480 11.815 57.800 ;
      LAYER met4 ;
        RECT 11.495 57.480 11.815 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 57.070 11.815 57.390 ;
      LAYER met4 ;
        RECT 11.495 57.070 11.815 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 56.660 11.815 56.980 ;
      LAYER met4 ;
        RECT 11.495 56.660 11.815 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.495 56.250 11.815 56.570 ;
      LAYER met4 ;
        RECT 11.495 56.250 11.815 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 60.350 11.410 60.670 ;
      LAYER met4 ;
        RECT 11.090 60.350 11.410 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 59.940 11.410 60.260 ;
      LAYER met4 ;
        RECT 11.090 59.940 11.410 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 59.530 11.410 59.850 ;
      LAYER met4 ;
        RECT 11.090 59.530 11.410 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 59.120 11.410 59.440 ;
      LAYER met4 ;
        RECT 11.090 59.120 11.410 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 58.710 11.410 59.030 ;
      LAYER met4 ;
        RECT 11.090 58.710 11.410 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 58.300 11.410 58.620 ;
      LAYER met4 ;
        RECT 11.090 58.300 11.410 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 57.890 11.410 58.210 ;
      LAYER met4 ;
        RECT 11.090 57.890 11.410 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 57.480 11.410 57.800 ;
      LAYER met4 ;
        RECT 11.090 57.480 11.410 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 57.070 11.410 57.390 ;
      LAYER met4 ;
        RECT 11.090 57.070 11.410 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 56.660 11.410 56.980 ;
      LAYER met4 ;
        RECT 11.090 56.660 11.410 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.090 56.250 11.410 56.570 ;
      LAYER met4 ;
        RECT 11.090 56.250 11.410 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 60.350 11.005 60.670 ;
      LAYER met4 ;
        RECT 10.685 60.350 11.005 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 59.940 11.005 60.260 ;
      LAYER met4 ;
        RECT 10.685 59.940 11.005 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 59.530 11.005 59.850 ;
      LAYER met4 ;
        RECT 10.685 59.530 11.005 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 59.120 11.005 59.440 ;
      LAYER met4 ;
        RECT 10.685 59.120 11.005 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 58.710 11.005 59.030 ;
      LAYER met4 ;
        RECT 10.685 58.710 11.005 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 58.300 11.005 58.620 ;
      LAYER met4 ;
        RECT 10.685 58.300 11.005 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 57.890 11.005 58.210 ;
      LAYER met4 ;
        RECT 10.685 57.890 11.005 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 57.480 11.005 57.800 ;
      LAYER met4 ;
        RECT 10.685 57.480 11.005 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 57.070 11.005 57.390 ;
      LAYER met4 ;
        RECT 10.685 57.070 11.005 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 56.660 11.005 56.980 ;
      LAYER met4 ;
        RECT 10.685 56.660 11.005 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.685 56.250 11.005 56.570 ;
      LAYER met4 ;
        RECT 10.685 56.250 11.005 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 60.350 10.600 60.670 ;
      LAYER met4 ;
        RECT 10.280 60.350 10.600 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 59.940 10.600 60.260 ;
      LAYER met4 ;
        RECT 10.280 59.940 10.600 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 59.530 10.600 59.850 ;
      LAYER met4 ;
        RECT 10.280 59.530 10.600 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 59.120 10.600 59.440 ;
      LAYER met4 ;
        RECT 10.280 59.120 10.600 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 58.710 10.600 59.030 ;
      LAYER met4 ;
        RECT 10.280 58.710 10.600 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 58.300 10.600 58.620 ;
      LAYER met4 ;
        RECT 10.280 58.300 10.600 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 57.890 10.600 58.210 ;
      LAYER met4 ;
        RECT 10.280 57.890 10.600 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 57.480 10.600 57.800 ;
      LAYER met4 ;
        RECT 10.280 57.480 10.600 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 57.070 10.600 57.390 ;
      LAYER met4 ;
        RECT 10.280 57.070 10.600 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 56.660 10.600 56.980 ;
      LAYER met4 ;
        RECT 10.280 56.660 10.600 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.280 56.250 10.600 56.570 ;
      LAYER met4 ;
        RECT 10.280 56.250 10.600 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 60.350 10.195 60.670 ;
      LAYER met4 ;
        RECT 9.875 60.350 10.195 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 59.940 10.195 60.260 ;
      LAYER met4 ;
        RECT 9.875 59.940 10.195 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 59.530 10.195 59.850 ;
      LAYER met4 ;
        RECT 9.875 59.530 10.195 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 59.120 10.195 59.440 ;
      LAYER met4 ;
        RECT 9.875 59.120 10.195 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 58.710 10.195 59.030 ;
      LAYER met4 ;
        RECT 9.875 58.710 10.195 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 58.300 10.195 58.620 ;
      LAYER met4 ;
        RECT 9.875 58.300 10.195 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 57.890 10.195 58.210 ;
      LAYER met4 ;
        RECT 9.875 57.890 10.195 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 57.480 10.195 57.800 ;
      LAYER met4 ;
        RECT 9.875 57.480 10.195 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 57.070 10.195 57.390 ;
      LAYER met4 ;
        RECT 9.875 57.070 10.195 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 56.660 10.195 56.980 ;
      LAYER met4 ;
        RECT 9.875 56.660 10.195 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.875 56.250 10.195 56.570 ;
      LAYER met4 ;
        RECT 9.875 56.250 10.195 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 60.350 9.790 60.670 ;
      LAYER met4 ;
        RECT 9.470 60.350 9.790 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 59.940 9.790 60.260 ;
      LAYER met4 ;
        RECT 9.470 59.940 9.790 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 59.530 9.790 59.850 ;
      LAYER met4 ;
        RECT 9.470 59.530 9.790 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 59.120 9.790 59.440 ;
      LAYER met4 ;
        RECT 9.470 59.120 9.790 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 58.710 9.790 59.030 ;
      LAYER met4 ;
        RECT 9.470 58.710 9.790 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 58.300 9.790 58.620 ;
      LAYER met4 ;
        RECT 9.470 58.300 9.790 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 57.890 9.790 58.210 ;
      LAYER met4 ;
        RECT 9.470 57.890 9.790 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 57.480 9.790 57.800 ;
      LAYER met4 ;
        RECT 9.470 57.480 9.790 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 57.070 9.790 57.390 ;
      LAYER met4 ;
        RECT 9.470 57.070 9.790 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 56.660 9.790 56.980 ;
      LAYER met4 ;
        RECT 9.470 56.660 9.790 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.470 56.250 9.790 56.570 ;
      LAYER met4 ;
        RECT 9.470 56.250 9.790 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 60.350 9.385 60.670 ;
      LAYER met4 ;
        RECT 9.065 60.350 9.385 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 59.940 9.385 60.260 ;
      LAYER met4 ;
        RECT 9.065 59.940 9.385 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 59.530 9.385 59.850 ;
      LAYER met4 ;
        RECT 9.065 59.530 9.385 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 59.120 9.385 59.440 ;
      LAYER met4 ;
        RECT 9.065 59.120 9.385 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 58.710 9.385 59.030 ;
      LAYER met4 ;
        RECT 9.065 58.710 9.385 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 58.300 9.385 58.620 ;
      LAYER met4 ;
        RECT 9.065 58.300 9.385 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 57.890 9.385 58.210 ;
      LAYER met4 ;
        RECT 9.065 57.890 9.385 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 57.480 9.385 57.800 ;
      LAYER met4 ;
        RECT 9.065 57.480 9.385 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 57.070 9.385 57.390 ;
      LAYER met4 ;
        RECT 9.065 57.070 9.385 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 56.660 9.385 56.980 ;
      LAYER met4 ;
        RECT 9.065 56.660 9.385 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.065 56.250 9.385 56.570 ;
      LAYER met4 ;
        RECT 9.065 56.250 9.385 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 60.350 8.980 60.670 ;
      LAYER met4 ;
        RECT 8.660 60.350 8.980 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 59.940 8.980 60.260 ;
      LAYER met4 ;
        RECT 8.660 59.940 8.980 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 59.530 8.980 59.850 ;
      LAYER met4 ;
        RECT 8.660 59.530 8.980 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 59.120 8.980 59.440 ;
      LAYER met4 ;
        RECT 8.660 59.120 8.980 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 58.710 8.980 59.030 ;
      LAYER met4 ;
        RECT 8.660 58.710 8.980 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 58.300 8.980 58.620 ;
      LAYER met4 ;
        RECT 8.660 58.300 8.980 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 57.890 8.980 58.210 ;
      LAYER met4 ;
        RECT 8.660 57.890 8.980 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 57.480 8.980 57.800 ;
      LAYER met4 ;
        RECT 8.660 57.480 8.980 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 57.070 8.980 57.390 ;
      LAYER met4 ;
        RECT 8.660 57.070 8.980 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 56.660 8.980 56.980 ;
      LAYER met4 ;
        RECT 8.660 56.660 8.980 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.660 56.250 8.980 56.570 ;
      LAYER met4 ;
        RECT 8.660 56.250 8.980 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 60.350 8.575 60.670 ;
      LAYER met4 ;
        RECT 8.255 60.350 8.575 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 59.940 8.575 60.260 ;
      LAYER met4 ;
        RECT 8.255 59.940 8.575 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 59.530 8.575 59.850 ;
      LAYER met4 ;
        RECT 8.255 59.530 8.575 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 59.120 8.575 59.440 ;
      LAYER met4 ;
        RECT 8.255 59.120 8.575 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 58.710 8.575 59.030 ;
      LAYER met4 ;
        RECT 8.255 58.710 8.575 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 58.300 8.575 58.620 ;
      LAYER met4 ;
        RECT 8.255 58.300 8.575 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 57.890 8.575 58.210 ;
      LAYER met4 ;
        RECT 8.255 57.890 8.575 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 57.480 8.575 57.800 ;
      LAYER met4 ;
        RECT 8.255 57.480 8.575 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 57.070 8.575 57.390 ;
      LAYER met4 ;
        RECT 8.255 57.070 8.575 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 56.660 8.575 56.980 ;
      LAYER met4 ;
        RECT 8.255 56.660 8.575 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.255 56.250 8.575 56.570 ;
      LAYER met4 ;
        RECT 8.255 56.250 8.575 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 60.350 8.170 60.670 ;
      LAYER met4 ;
        RECT 7.850 60.350 8.170 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 59.940 8.170 60.260 ;
      LAYER met4 ;
        RECT 7.850 59.940 8.170 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 59.530 8.170 59.850 ;
      LAYER met4 ;
        RECT 7.850 59.530 8.170 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 59.120 8.170 59.440 ;
      LAYER met4 ;
        RECT 7.850 59.120 8.170 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 58.710 8.170 59.030 ;
      LAYER met4 ;
        RECT 7.850 58.710 8.170 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 58.300 8.170 58.620 ;
      LAYER met4 ;
        RECT 7.850 58.300 8.170 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 57.890 8.170 58.210 ;
      LAYER met4 ;
        RECT 7.850 57.890 8.170 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 57.480 8.170 57.800 ;
      LAYER met4 ;
        RECT 7.850 57.480 8.170 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 57.070 8.170 57.390 ;
      LAYER met4 ;
        RECT 7.850 57.070 8.170 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 56.660 8.170 56.980 ;
      LAYER met4 ;
        RECT 7.850 56.660 8.170 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.850 56.250 8.170 56.570 ;
      LAYER met4 ;
        RECT 7.850 56.250 8.170 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 60.350 7.765 60.670 ;
      LAYER met4 ;
        RECT 7.445 60.350 7.765 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 59.940 7.765 60.260 ;
      LAYER met4 ;
        RECT 7.445 59.940 7.765 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 59.530 7.765 59.850 ;
      LAYER met4 ;
        RECT 7.445 59.530 7.765 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 59.120 7.765 59.440 ;
      LAYER met4 ;
        RECT 7.445 59.120 7.765 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 58.710 7.765 59.030 ;
      LAYER met4 ;
        RECT 7.445 58.710 7.765 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 58.300 7.765 58.620 ;
      LAYER met4 ;
        RECT 7.445 58.300 7.765 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 57.890 7.765 58.210 ;
      LAYER met4 ;
        RECT 7.445 57.890 7.765 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 57.480 7.765 57.800 ;
      LAYER met4 ;
        RECT 7.445 57.480 7.765 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 57.070 7.765 57.390 ;
      LAYER met4 ;
        RECT 7.445 57.070 7.765 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 56.660 7.765 56.980 ;
      LAYER met4 ;
        RECT 7.445 56.660 7.765 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.445 56.250 7.765 56.570 ;
      LAYER met4 ;
        RECT 7.445 56.250 7.765 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 60.350 7.360 60.670 ;
      LAYER met4 ;
        RECT 7.040 60.350 7.360 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 59.940 7.360 60.260 ;
      LAYER met4 ;
        RECT 7.040 59.940 7.360 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 59.530 7.360 59.850 ;
      LAYER met4 ;
        RECT 7.040 59.530 7.360 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 59.120 7.360 59.440 ;
      LAYER met4 ;
        RECT 7.040 59.120 7.360 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 58.710 7.360 59.030 ;
      LAYER met4 ;
        RECT 7.040 58.710 7.360 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 58.300 7.360 58.620 ;
      LAYER met4 ;
        RECT 7.040 58.300 7.360 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 57.890 7.360 58.210 ;
      LAYER met4 ;
        RECT 7.040 57.890 7.360 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 57.480 7.360 57.800 ;
      LAYER met4 ;
        RECT 7.040 57.480 7.360 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 57.070 7.360 57.390 ;
      LAYER met4 ;
        RECT 7.040 57.070 7.360 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 56.660 7.360 56.980 ;
      LAYER met4 ;
        RECT 7.040 56.660 7.360 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.040 56.250 7.360 56.570 ;
      LAYER met4 ;
        RECT 7.040 56.250 7.360 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 60.350 6.955 60.670 ;
      LAYER met4 ;
        RECT 6.635 60.350 6.955 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 59.940 6.955 60.260 ;
      LAYER met4 ;
        RECT 6.635 59.940 6.955 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 59.530 6.955 59.850 ;
      LAYER met4 ;
        RECT 6.635 59.530 6.955 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 59.120 6.955 59.440 ;
      LAYER met4 ;
        RECT 6.635 59.120 6.955 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 58.710 6.955 59.030 ;
      LAYER met4 ;
        RECT 6.635 58.710 6.955 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 58.300 6.955 58.620 ;
      LAYER met4 ;
        RECT 6.635 58.300 6.955 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 57.890 6.955 58.210 ;
      LAYER met4 ;
        RECT 6.635 57.890 6.955 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 57.480 6.955 57.800 ;
      LAYER met4 ;
        RECT 6.635 57.480 6.955 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 57.070 6.955 57.390 ;
      LAYER met4 ;
        RECT 6.635 57.070 6.955 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 56.660 6.955 56.980 ;
      LAYER met4 ;
        RECT 6.635 56.660 6.955 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 56.250 6.955 56.570 ;
      LAYER met4 ;
        RECT 6.635 56.250 6.955 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 60.350 6.550 60.670 ;
      LAYER met4 ;
        RECT 6.230 60.350 6.550 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 59.940 6.550 60.260 ;
      LAYER met4 ;
        RECT 6.230 59.940 6.550 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 59.530 6.550 59.850 ;
      LAYER met4 ;
        RECT 6.230 59.530 6.550 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 59.120 6.550 59.440 ;
      LAYER met4 ;
        RECT 6.230 59.120 6.550 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 58.710 6.550 59.030 ;
      LAYER met4 ;
        RECT 6.230 58.710 6.550 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 58.300 6.550 58.620 ;
      LAYER met4 ;
        RECT 6.230 58.300 6.550 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 57.890 6.550 58.210 ;
      LAYER met4 ;
        RECT 6.230 57.890 6.550 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 57.480 6.550 57.800 ;
      LAYER met4 ;
        RECT 6.230 57.480 6.550 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 57.070 6.550 57.390 ;
      LAYER met4 ;
        RECT 6.230 57.070 6.550 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 56.660 6.550 56.980 ;
      LAYER met4 ;
        RECT 6.230 56.660 6.550 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.230 56.250 6.550 56.570 ;
      LAYER met4 ;
        RECT 6.230 56.250 6.550 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 60.350 6.145 60.670 ;
      LAYER met4 ;
        RECT 5.825 60.350 6.145 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 59.940 6.145 60.260 ;
      LAYER met4 ;
        RECT 5.825 59.940 6.145 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 59.530 6.145 59.850 ;
      LAYER met4 ;
        RECT 5.825 59.530 6.145 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 59.120 6.145 59.440 ;
      LAYER met4 ;
        RECT 5.825 59.120 6.145 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 58.710 6.145 59.030 ;
      LAYER met4 ;
        RECT 5.825 58.710 6.145 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 58.300 6.145 58.620 ;
      LAYER met4 ;
        RECT 5.825 58.300 6.145 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 57.890 6.145 58.210 ;
      LAYER met4 ;
        RECT 5.825 57.890 6.145 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 57.480 6.145 57.800 ;
      LAYER met4 ;
        RECT 5.825 57.480 6.145 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 57.070 6.145 57.390 ;
      LAYER met4 ;
        RECT 5.825 57.070 6.145 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 56.660 6.145 56.980 ;
      LAYER met4 ;
        RECT 5.825 56.660 6.145 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.825 56.250 6.145 56.570 ;
      LAYER met4 ;
        RECT 5.825 56.250 6.145 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 60.350 5.740 60.670 ;
      LAYER met4 ;
        RECT 5.420 60.350 5.740 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 59.940 5.740 60.260 ;
      LAYER met4 ;
        RECT 5.420 59.940 5.740 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 59.530 5.740 59.850 ;
      LAYER met4 ;
        RECT 5.420 59.530 5.740 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 59.120 5.740 59.440 ;
      LAYER met4 ;
        RECT 5.420 59.120 5.740 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 58.710 5.740 59.030 ;
      LAYER met4 ;
        RECT 5.420 58.710 5.740 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 58.300 5.740 58.620 ;
      LAYER met4 ;
        RECT 5.420 58.300 5.740 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 57.890 5.740 58.210 ;
      LAYER met4 ;
        RECT 5.420 57.890 5.740 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 57.480 5.740 57.800 ;
      LAYER met4 ;
        RECT 5.420 57.480 5.740 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 57.070 5.740 57.390 ;
      LAYER met4 ;
        RECT 5.420 57.070 5.740 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 56.660 5.740 56.980 ;
      LAYER met4 ;
        RECT 5.420 56.660 5.740 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.420 56.250 5.740 56.570 ;
      LAYER met4 ;
        RECT 5.420 56.250 5.740 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 60.350 5.335 60.670 ;
      LAYER met4 ;
        RECT 5.015 60.350 5.335 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 59.940 5.335 60.260 ;
      LAYER met4 ;
        RECT 5.015 59.940 5.335 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 59.530 5.335 59.850 ;
      LAYER met4 ;
        RECT 5.015 59.530 5.335 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 59.120 5.335 59.440 ;
      LAYER met4 ;
        RECT 5.015 59.120 5.335 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 58.710 5.335 59.030 ;
      LAYER met4 ;
        RECT 5.015 58.710 5.335 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 58.300 5.335 58.620 ;
      LAYER met4 ;
        RECT 5.015 58.300 5.335 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 57.890 5.335 58.210 ;
      LAYER met4 ;
        RECT 5.015 57.890 5.335 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 57.480 5.335 57.800 ;
      LAYER met4 ;
        RECT 5.015 57.480 5.335 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 57.070 5.335 57.390 ;
      LAYER met4 ;
        RECT 5.015 57.070 5.335 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 56.660 5.335 56.980 ;
      LAYER met4 ;
        RECT 5.015 56.660 5.335 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.015 56.250 5.335 56.570 ;
      LAYER met4 ;
        RECT 5.015 56.250 5.335 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 60.350 4.930 60.670 ;
      LAYER met4 ;
        RECT 4.610 60.350 4.930 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 59.940 4.930 60.260 ;
      LAYER met4 ;
        RECT 4.610 59.940 4.930 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 59.530 4.930 59.850 ;
      LAYER met4 ;
        RECT 4.610 59.530 4.930 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 59.120 4.930 59.440 ;
      LAYER met4 ;
        RECT 4.610 59.120 4.930 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 58.710 4.930 59.030 ;
      LAYER met4 ;
        RECT 4.610 58.710 4.930 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 58.300 4.930 58.620 ;
      LAYER met4 ;
        RECT 4.610 58.300 4.930 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 57.890 4.930 58.210 ;
      LAYER met4 ;
        RECT 4.610 57.890 4.930 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 57.480 4.930 57.800 ;
      LAYER met4 ;
        RECT 4.610 57.480 4.930 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 57.070 4.930 57.390 ;
      LAYER met4 ;
        RECT 4.610 57.070 4.930 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 56.660 4.930 56.980 ;
      LAYER met4 ;
        RECT 4.610 56.660 4.930 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.610 56.250 4.930 56.570 ;
      LAYER met4 ;
        RECT 4.610 56.250 4.930 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 60.350 4.525 60.670 ;
      LAYER met4 ;
        RECT 4.205 60.350 4.525 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 59.940 4.525 60.260 ;
      LAYER met4 ;
        RECT 4.205 59.940 4.525 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 59.530 4.525 59.850 ;
      LAYER met4 ;
        RECT 4.205 59.530 4.525 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 59.120 4.525 59.440 ;
      LAYER met4 ;
        RECT 4.205 59.120 4.525 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 58.710 4.525 59.030 ;
      LAYER met4 ;
        RECT 4.205 58.710 4.525 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 58.300 4.525 58.620 ;
      LAYER met4 ;
        RECT 4.205 58.300 4.525 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 57.890 4.525 58.210 ;
      LAYER met4 ;
        RECT 4.205 57.890 4.525 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 57.480 4.525 57.800 ;
      LAYER met4 ;
        RECT 4.205 57.480 4.525 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 57.070 4.525 57.390 ;
      LAYER met4 ;
        RECT 4.205 57.070 4.525 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 56.660 4.525 56.980 ;
      LAYER met4 ;
        RECT 4.205 56.660 4.525 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.205 56.250 4.525 56.570 ;
      LAYER met4 ;
        RECT 4.205 56.250 4.525 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 60.350 4.120 60.670 ;
      LAYER met4 ;
        RECT 3.800 60.350 4.120 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 59.940 4.120 60.260 ;
      LAYER met4 ;
        RECT 3.800 59.940 4.120 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 59.530 4.120 59.850 ;
      LAYER met4 ;
        RECT 3.800 59.530 4.120 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 59.120 4.120 59.440 ;
      LAYER met4 ;
        RECT 3.800 59.120 4.120 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 58.710 4.120 59.030 ;
      LAYER met4 ;
        RECT 3.800 58.710 4.120 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 58.300 4.120 58.620 ;
      LAYER met4 ;
        RECT 3.800 58.300 4.120 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 57.890 4.120 58.210 ;
      LAYER met4 ;
        RECT 3.800 57.890 4.120 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 57.480 4.120 57.800 ;
      LAYER met4 ;
        RECT 3.800 57.480 4.120 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 57.070 4.120 57.390 ;
      LAYER met4 ;
        RECT 3.800 57.070 4.120 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 56.660 4.120 56.980 ;
      LAYER met4 ;
        RECT 3.800 56.660 4.120 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 56.250 4.120 56.570 ;
      LAYER met4 ;
        RECT 3.800 56.250 4.120 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 60.350 3.715 60.670 ;
      LAYER met4 ;
        RECT 3.395 60.350 3.715 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 59.940 3.715 60.260 ;
      LAYER met4 ;
        RECT 3.395 59.940 3.715 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 59.530 3.715 59.850 ;
      LAYER met4 ;
        RECT 3.395 59.530 3.715 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 59.120 3.715 59.440 ;
      LAYER met4 ;
        RECT 3.395 59.120 3.715 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 58.710 3.715 59.030 ;
      LAYER met4 ;
        RECT 3.395 58.710 3.715 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 58.300 3.715 58.620 ;
      LAYER met4 ;
        RECT 3.395 58.300 3.715 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 57.890 3.715 58.210 ;
      LAYER met4 ;
        RECT 3.395 57.890 3.715 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 57.480 3.715 57.800 ;
      LAYER met4 ;
        RECT 3.395 57.480 3.715 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 57.070 3.715 57.390 ;
      LAYER met4 ;
        RECT 3.395 57.070 3.715 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 56.660 3.715 56.980 ;
      LAYER met4 ;
        RECT 3.395 56.660 3.715 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 56.250 3.715 56.570 ;
      LAYER met4 ;
        RECT 3.395 56.250 3.715 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 60.350 3.310 60.670 ;
      LAYER met4 ;
        RECT 2.990 60.350 3.310 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 59.940 3.310 60.260 ;
      LAYER met4 ;
        RECT 2.990 59.940 3.310 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 59.530 3.310 59.850 ;
      LAYER met4 ;
        RECT 2.990 59.530 3.310 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 59.120 3.310 59.440 ;
      LAYER met4 ;
        RECT 2.990 59.120 3.310 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 58.710 3.310 59.030 ;
      LAYER met4 ;
        RECT 2.990 58.710 3.310 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 58.300 3.310 58.620 ;
      LAYER met4 ;
        RECT 2.990 58.300 3.310 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 57.890 3.310 58.210 ;
      LAYER met4 ;
        RECT 2.990 57.890 3.310 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 57.480 3.310 57.800 ;
      LAYER met4 ;
        RECT 2.990 57.480 3.310 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 57.070 3.310 57.390 ;
      LAYER met4 ;
        RECT 2.990 57.070 3.310 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 56.660 3.310 56.980 ;
      LAYER met4 ;
        RECT 2.990 56.660 3.310 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.990 56.250 3.310 56.570 ;
      LAYER met4 ;
        RECT 2.990 56.250 3.310 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 60.350 2.900 60.670 ;
      LAYER met4 ;
        RECT 2.580 60.350 2.900 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 59.940 2.900 60.260 ;
      LAYER met4 ;
        RECT 2.580 59.940 2.900 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 59.530 2.900 59.850 ;
      LAYER met4 ;
        RECT 2.580 59.530 2.900 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 59.120 2.900 59.440 ;
      LAYER met4 ;
        RECT 2.580 59.120 2.900 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 58.710 2.900 59.030 ;
      LAYER met4 ;
        RECT 2.580 58.710 2.900 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 58.300 2.900 58.620 ;
      LAYER met4 ;
        RECT 2.580 58.300 2.900 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 57.890 2.900 58.210 ;
      LAYER met4 ;
        RECT 2.580 57.890 2.900 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 57.480 2.900 57.800 ;
      LAYER met4 ;
        RECT 2.580 57.480 2.900 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 57.070 2.900 57.390 ;
      LAYER met4 ;
        RECT 2.580 57.070 2.900 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 56.660 2.900 56.980 ;
      LAYER met4 ;
        RECT 2.580 56.660 2.900 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.580 56.250 2.900 56.570 ;
      LAYER met4 ;
        RECT 2.580 56.250 2.900 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 60.350 2.490 60.670 ;
      LAYER met4 ;
        RECT 2.170 60.350 2.490 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 59.940 2.490 60.260 ;
      LAYER met4 ;
        RECT 2.170 59.940 2.490 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 59.530 2.490 59.850 ;
      LAYER met4 ;
        RECT 2.170 59.530 2.490 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 59.120 2.490 59.440 ;
      LAYER met4 ;
        RECT 2.170 59.120 2.490 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 58.710 2.490 59.030 ;
      LAYER met4 ;
        RECT 2.170 58.710 2.490 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 58.300 2.490 58.620 ;
      LAYER met4 ;
        RECT 2.170 58.300 2.490 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 57.890 2.490 58.210 ;
      LAYER met4 ;
        RECT 2.170 57.890 2.490 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 57.480 2.490 57.800 ;
      LAYER met4 ;
        RECT 2.170 57.480 2.490 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 57.070 2.490 57.390 ;
      LAYER met4 ;
        RECT 2.170 57.070 2.490 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 56.660 2.490 56.980 ;
      LAYER met4 ;
        RECT 2.170 56.660 2.490 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.170 56.250 2.490 56.570 ;
      LAYER met4 ;
        RECT 2.170 56.250 2.490 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 60.350 2.080 60.670 ;
      LAYER met4 ;
        RECT 1.760 60.350 2.080 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 59.940 2.080 60.260 ;
      LAYER met4 ;
        RECT 1.760 59.940 2.080 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 59.530 2.080 59.850 ;
      LAYER met4 ;
        RECT 1.760 59.530 2.080 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 59.120 2.080 59.440 ;
      LAYER met4 ;
        RECT 1.760 59.120 2.080 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 58.710 2.080 59.030 ;
      LAYER met4 ;
        RECT 1.760 58.710 2.080 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 58.300 2.080 58.620 ;
      LAYER met4 ;
        RECT 1.760 58.300 2.080 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 57.890 2.080 58.210 ;
      LAYER met4 ;
        RECT 1.760 57.890 2.080 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 57.480 2.080 57.800 ;
      LAYER met4 ;
        RECT 1.760 57.480 2.080 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 57.070 2.080 57.390 ;
      LAYER met4 ;
        RECT 1.760 57.070 2.080 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 56.660 2.080 56.980 ;
      LAYER met4 ;
        RECT 1.760 56.660 2.080 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.760 56.250 2.080 56.570 ;
      LAYER met4 ;
        RECT 1.760 56.250 2.080 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 60.350 1.670 60.670 ;
      LAYER met4 ;
        RECT 1.350 60.350 1.670 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 59.940 1.670 60.260 ;
      LAYER met4 ;
        RECT 1.350 59.940 1.670 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 59.530 1.670 59.850 ;
      LAYER met4 ;
        RECT 1.350 59.530 1.670 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 59.120 1.670 59.440 ;
      LAYER met4 ;
        RECT 1.350 59.120 1.670 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 58.710 1.670 59.030 ;
      LAYER met4 ;
        RECT 1.350 58.710 1.670 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 58.300 1.670 58.620 ;
      LAYER met4 ;
        RECT 1.350 58.300 1.670 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 57.890 1.670 58.210 ;
      LAYER met4 ;
        RECT 1.350 57.890 1.670 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 57.480 1.670 57.800 ;
      LAYER met4 ;
        RECT 1.350 57.480 1.670 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 57.070 1.670 57.390 ;
      LAYER met4 ;
        RECT 1.350 57.070 1.670 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 56.660 1.670 56.980 ;
      LAYER met4 ;
        RECT 1.350 56.660 1.670 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.350 56.250 1.670 56.570 ;
      LAYER met4 ;
        RECT 1.350 56.250 1.670 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 60.350 1.260 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 59.940 1.260 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 59.530 1.260 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 59.120 1.260 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 58.710 1.260 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 58.300 1.260 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 57.890 1.260 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 57.480 1.260 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 57.070 1.260 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 56.660 1.260 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.940 56.250 1.260 56.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 60.350 0.850 60.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 59.940 0.850 60.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 59.530 0.850 59.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 59.120 0.850 59.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 58.710 0.850 59.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 58.300 0.850 58.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 57.890 0.850 58.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 57.480 0.850 57.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 57.070 0.850 57.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 56.660 0.850 56.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.530 56.250 0.850 56.570 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
  END VSWITCH
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
  END VCCHIB
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
  END VDDIO_Q
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  OBS
      LAYER met3 ;
        RECT 0.500 56.240 24.400 198.000 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 94.585 75.000 172.185 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__overlay_vssio_lvc

#--------EOF---------

MACRO sky130_fd_io__top_gpio_ovtv2
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_gpio_ovtv2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730 58.335 140.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 58.235 140.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730 31.985 140.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 31.885 140.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
  END VSWITCH
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730 25.935 140.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730 175.785 140.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.365 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 175.785 140.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 25.835 140.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.365 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
  END VSSIO
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730 41.685 140.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 41.585 140.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
  END VSSD
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 138.730 36.840 140.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730 47.735 140.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 2.040 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 51.645 140.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 140.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 140.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 36.735 140.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 2.040 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
  END VSSA
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730 64.185 140.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 64.085 140.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730 70.035 140.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 138.730 19.885 140.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 19.785 140.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 70.035 140.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
  END VDDIO
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 139.035 15.035 140.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 139.035 14.935 140.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
  END VDDA
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730 2.135 140.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 2.035 140.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
  END VCCHIB
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 138.730 8.985 140.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.730 8.885 140.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
  END VCCD
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 17.930 117.530 86.325 162.905 ;
    END
  END PAD
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.930 53.125 140.000 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 38.675 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.710 48.365 140.000 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 85.865 51.345 ;
    END
  END AMUXBUS_B
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.125 0.000 129.455 20.955 ;
    END
  END DM[0]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.275 0.000 128.605 20.180 ;
    END
  END DM[1]
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.395 0.000 108.725 20.640 ;
    END
  END DM[2]
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.545 0.000 107.875 8.060 ;
    END
  END INP_DIS
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.665 0.000 87.995 20.980 ;
    END
  END VTRIP_SEL
  PIN IB_MODE_SEL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 86.815 0.000 87.145 20.980 ;
    END
  END IB_MODE_SEL[0]
  PIN IB_MODE_SEL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.935 0.000 67.265 20.980 ;
    END
  END IB_MODE_SEL[1]
  PIN SLEW_CTL[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.085 0.000 66.415 20.980 ;
    END
  END SLEW_CTL[0]
  PIN SLEW_CTL[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.205 0.000 46.535 20.980 ;
    END
  END SLEW_CTL[1]
  PIN HYS_TRIM
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.355 0.000 45.685 8.060 ;
    END
  END HYS_TRIM
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.355 0.000 27.685 14.055 ;
    END
  END HLD_OVR
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.135 0.000 22.465 30.150 ;
    END
  END ENABLE_H
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 19.635 0.000 19.965 17.985 ;
    END
  END HLD_H_N
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.770 0.000 9.100 7.915 ;
    END
  END ENABLE_VDDA_H
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.115 0.000 8.445 14.070 ;
    END
  END ANALOG_EN
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.110 0.000 7.440 0.670 ;
    END
  END ENABLE_INP_H
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.380 0.000 20.710 11.310 ;
    END
  END IN
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 24.380 0.000 24.710 0.940 ;
    END
  END IN_H
  PIN VINREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 44.035 0.000 44.365 4.885 ;
    END
  END VINREF
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 74.125 0.000 74.455 14.865 ;
    END
  END OUT
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.235 0.000 65.565 1.165 ;
    END
  END ANALOG_POL
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 51.655 0.000 51.985 8.060 ;
    END
  END ANALOG_SEL
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.140 0.000 125.470 11.965 ;
    END
  END SLOW
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 124.445 0.000 124.775 8.060 ;
    END
  END OE_N
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.975 0.000 130.305 61.655 ;
    END
  END TIE_HI_ESD
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.290 0.000 115.890 39.035 ;
    END
  END TIE_LO_ESD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1.600 0.000 2.200 5.470 ;
    END
  END PAD_A_ESD_0_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.330 0.000 0.930 71.380 ;
    END
  END PAD_A_ESD_1_H
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2.885 0.000 3.485 5.900 ;
    END
  END PAD_A_NOESD_H
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.765 0.000 6.365 12.470 ;
    END
  END ENABLE_VSWITCH_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.845 0.000 96.215 20.755 ;
    END
  END ENABLE_VDDIO
  OBS
      LAYER nwell ;
        RECT 118.950 184.430 140.420 185.605 ;
        RECT 130.895 183.580 140.420 184.430 ;
        RECT 133.940 180.105 140.420 183.580 ;
        RECT 133.900 174.850 140.420 180.105 ;
        RECT 133.175 161.940 140.420 174.850 ;
        RECT 133.740 128.090 140.420 161.940 ;
        RECT 132.500 122.180 140.420 128.090 ;
        RECT 118.950 117.425 140.420 122.180 ;
      LAYER pwell ;
        RECT 114.115 114.365 140.130 116.895 ;
        RECT 131.245 110.270 140.130 114.365 ;
      LAYER nwell ;
        RECT 6.155 107.630 141.055 109.740 ;
        RECT 138.945 67.930 141.055 107.630 ;
        RECT 6.155 66.420 141.055 67.930 ;
        RECT 132.725 63.655 140.680 65.015 ;
        RECT 139.320 54.255 140.680 63.655 ;
        RECT 132.725 52.895 140.680 54.255 ;
      LAYER pwell ;
        RECT 11.470 18.640 140.130 20.430 ;
        RECT 32.115 17.020 140.130 18.640 ;
      LAYER nwell ;
        RECT -0.400 10.495 11.880 11.925 ;
        RECT -0.400 1.430 1.030 10.495 ;
        RECT -0.400 0.000 11.880 1.430 ;
      LAYER li1 ;
        RECT 0.230 184.675 140.000 199.780 ;
        RECT 0.230 117.690 140.085 184.675 ;
        RECT 0.230 116.765 140.000 117.690 ;
        RECT 0.230 110.400 140.145 116.765 ;
        RECT 0.230 109.110 140.000 110.400 ;
        RECT 0.230 67.170 140.475 109.110 ;
        RECT 0.230 66.750 140.425 67.170 ;
        RECT 0.230 64.685 140.000 66.750 ;
        RECT 0.230 53.225 140.350 64.685 ;
        RECT 0.230 0.200 140.000 53.225 ;
      LAYER met1 ;
        RECT 0.080 184.720 140.000 199.810 ;
        RECT 0.080 183.205 140.145 184.720 ;
        RECT 0.080 117.630 140.115 183.205 ;
        POLYGON 140.115 183.205 140.145 183.205 140.115 183.175 ;
        RECT 0.080 108.870 140.000 117.630 ;
        RECT 0.080 67.170 140.475 108.870 ;
        RECT 0.080 64.685 140.000 67.170 ;
        RECT 0.080 53.225 140.350 64.685 ;
        RECT 0.080 0.000 140.000 53.225 ;
      LAYER met2 ;
        RECT 0.080 184.720 140.000 199.955 ;
        RECT 0.080 182.890 140.130 184.720 ;
        RECT 0.080 68.140 140.000 182.890 ;
        RECT 0.080 63.715 140.325 68.140 ;
        RECT 0.080 0.000 140.000 63.715 ;
      LAYER met3 ;
        RECT 0.330 71.780 140.000 199.715 ;
        RECT 1.330 62.055 140.000 71.780 ;
        RECT 1.330 39.435 129.575 62.055 ;
        RECT 1.330 30.550 114.890 39.435 ;
        RECT 1.330 18.385 21.735 30.550 ;
        RECT 1.330 14.470 19.235 18.385 ;
        RECT 1.330 12.870 7.715 14.470 ;
        RECT 1.330 6.300 5.365 12.870 ;
        RECT 1.330 5.870 2.485 6.300 ;
        RECT 3.885 0.000 5.365 6.300 ;
        RECT 6.765 1.070 7.715 12.870 ;
        RECT 8.845 8.315 19.235 14.470 ;
        RECT 20.365 11.710 21.735 18.385 ;
        RECT 9.500 0.000 19.235 8.315 ;
        RECT 21.110 0.000 21.735 11.710 ;
        RECT 22.865 21.380 114.890 30.550 ;
        RECT 22.865 14.455 45.805 21.380 ;
        RECT 22.865 1.340 26.955 14.455 ;
        RECT 22.865 0.000 23.980 1.340 ;
        RECT 25.110 0.000 26.955 1.340 ;
        RECT 28.085 8.460 45.805 14.455 ;
        RECT 46.935 8.460 65.685 21.380 ;
        RECT 28.085 5.285 44.955 8.460 ;
        RECT 28.085 0.000 43.635 5.285 ;
        RECT 44.765 0.000 44.955 5.285 ;
        RECT 46.935 0.000 51.255 8.460 ;
        RECT 52.385 1.565 65.685 8.460 ;
        RECT 67.665 15.265 86.415 21.380 ;
        RECT 52.385 0.000 64.835 1.565 ;
        RECT 67.665 0.000 73.725 15.265 ;
        RECT 74.855 0.000 86.415 15.265 ;
        RECT 88.395 21.155 114.890 21.380 ;
        RECT 88.395 0.000 95.445 21.155 ;
        RECT 96.615 21.040 114.890 21.155 ;
        RECT 96.615 8.460 107.995 21.040 ;
        RECT 96.615 0.000 107.145 8.460 ;
        RECT 109.125 0.000 114.890 21.040 ;
        RECT 116.290 21.355 129.575 39.435 ;
        RECT 116.290 20.580 128.725 21.355 ;
        RECT 116.290 12.365 127.875 20.580 ;
        RECT 116.290 8.460 124.740 12.365 ;
        RECT 116.290 0.000 124.045 8.460 ;
        RECT 125.870 0.000 127.875 12.365 ;
        RECT 130.705 0.000 140.000 62.055 ;
      LAYER met4 ;
        RECT 1.765 175.385 138.330 200.000 ;
        RECT 0.965 95.400 139.035 175.385 ;
        RECT 1.670 69.635 138.330 95.400 ;
        RECT 0.965 68.935 139.035 69.635 ;
        RECT 1.670 63.685 138.330 68.935 ;
        RECT 0.965 63.085 139.035 63.685 ;
        RECT 1.670 57.835 138.330 63.085 ;
        RECT 0.965 57.135 139.035 57.835 ;
        RECT 39.075 52.725 48.530 56.005 ;
        RECT 2.440 51.745 138.330 52.725 ;
        RECT 86.265 48.465 99.310 51.745 ;
        RECT 0.965 46.635 139.035 47.335 ;
        RECT 1.670 41.185 138.330 46.635 ;
        RECT 0.965 40.585 139.035 41.185 ;
        RECT 1.670 36.335 138.330 40.585 ;
        RECT 0.965 35.735 139.035 36.335 ;
        RECT 1.670 31.485 138.330 35.735 ;
        RECT 0.965 30.885 139.035 31.485 ;
        RECT 1.670 25.435 138.330 30.885 ;
        RECT 0.965 24.835 139.035 25.435 ;
        RECT 1.670 19.385 138.330 24.835 ;
        RECT 0.965 18.785 139.035 19.385 ;
        RECT 1.365 14.535 138.635 18.785 ;
        RECT 0.965 13.935 139.035 14.535 ;
        RECT 1.670 8.485 138.330 13.935 ;
        RECT 0.965 7.885 139.035 8.485 ;
        RECT 1.670 1.635 138.330 7.885 ;
        RECT 0.965 1.160 139.035 1.635 ;
      LAYER met5 ;
        RECT 2.965 174.185 137.130 200.000 ;
        RECT 0.000 164.505 140.000 174.185 ;
        RECT 0.000 115.930 16.330 164.505 ;
        RECT 87.925 115.930 140.000 164.505 ;
        RECT 0.000 96.585 140.000 115.930 ;
        RECT 2.870 58.335 137.130 96.585 ;
        RECT 3.640 46.135 137.130 58.335 ;
        RECT 2.870 18.285 137.130 46.135 ;
        RECT 2.565 15.035 137.435 18.285 ;
        RECT 2.870 2.135 137.130 15.035 ;
  END
END sky130_fd_io__top_gpio_ovtv2

#--------EOF---------

MACRO sky130_fd_io__top_gpiov2
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_gpiov2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.200 104.560 73.800 167.010 ;
    END
  END PAD
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 13.910 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.705 41.585 80.000 46.235 ;
    END
  END VSSD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 52.145 51.345 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.465 48.365 80.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 36.440 56.105 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.760 53.125 80.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 6.860 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.945 64.085 80.000 68.535 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.460 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 7.430 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 68.030 70.035 80.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.735 19.785 80.000 24.435 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 22.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.850 31.885 80.000 35.335 ;
    END
  END VSWITCH
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 19.330 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.530 25.835 80.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.230 175.785 80.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 25.550 200.000 ;
    END
  END VSSIO
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 24.590 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.570 14.935 80.000 18.385 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 34.235 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.265 8.885 80.000 13.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 11.150 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.810 2.035 80.000 7.485 ;
    END
  END VCCHIB
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 2.610 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 2.610 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 2.610 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 5.435 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.310 36.735 80.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 56.405 80.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 47.735 80.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.090 51.645 80.000 52.825 ;
    END
  END VSSA
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 69.845 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.575 58.235 80.000 62.685 ;
    END
  END VSSIO_Q
  PIN PAD_A_NOESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 106.585 5.470 118.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.820 0.000 63.890 14.845 ;
    END
    PORT
      LAYER met4 ;
        RECT 9.810 121.205 12.500 121.250 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.830 104.560 9.855 106.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.570 120.010 9.800 121.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 7.515 118.955 8.570 120.010 ;
    END
  END PAD_A_NOESD_H
  PIN ANALOG_POL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.865 0.000 46.195 36.805 ;
    END
  END ANALOG_POL
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.580 0.000 78.910 184.775 ;
    END
  END ENABLE_VDDIO
  PIN IN_H
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.400 0.000 1.020 178.485 ;
    END
  END IN_H
  PIN IN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.240 0.000 79.570 189.560 ;
    END
  END IN
  PIN DM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.855 0.000 50.115 0.545 ;
    END
  END DM[0]
  PIN DM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.835 0.000 67.095 1.195 ;
    END
  END DM[1]
  PIN DM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.490 0.000 28.750 4.070 ;
    END
  END DM[2]
  PIN HLD_H_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.815 0.000 32.075 3.340 ;
    END
  END HLD_H_N
  PIN HLD_OVR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.600 0.000 26.860 2.705 ;
    END
  END HLD_OVR
  PIN INP_DIS
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.245 0.000 45.505 5.090 ;
    END
  END INP_DIS
  PIN ENABLE_VDDA_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.755 0.000 13.015 5.350 ;
    END
  END ENABLE_VDDA_H
  PIN VTRIP_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.130 0.000 6.390 1.550 ;
    END
  END VTRIP_SEL
  PIN OE_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.375 0.000 3.605 4.475 ;
    END
  END OE_N
  PIN OUT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.355 0.000 22.615 6.425 ;
    END
  END OUT
  PIN SLOW
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.610 0.000 77.870 1.185 ;
    END
  END SLOW
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.715 0.000 79.915 177.870 ;
    END
  END TIE_LO_ESD
  PIN PAD_A_ESD_0_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.280 0.000 76.920 2.055 ;
    END
  END PAD_A_ESD_0_H
  PIN ANALOG_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.750 0.000 31.010 2.265 ;
    END
  END ANALOG_SEL
  PIN ENABLE_INP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.390 0.000 38.650 3.090 ;
    END
  END ENABLE_INP_H
  PIN PAD_A_ESD_1_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.275 0.000 68.925 2.270 ;
    END
  END PAD_A_ESD_1_H
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.705 0.000 78.905 1.215 ;
    END
  END TIE_HI_ESD
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.460 0.000 35.720 1.550 ;
    END
  END ENABLE_H
  PIN IB_MODE_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.420 0.000 5.650 4.475 ;
    END
  END IB_MODE_SEL
  PIN ENABLE_VSWITCH_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.310 0.000 16.570 2.320 ;
    END
  END ENABLE_VSWITCH_H
  PIN ANALOG_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 62.430 0.000 62.690 1.305 ;
    END
  END ANALOG_EN
  OBS
      LAYER nwell ;
        RECT -0.415 173.545 80.435 178.975 ;
        RECT -0.415 170.475 7.515 173.545 ;
        RECT 66.970 170.475 80.435 173.545 ;
        RECT -0.415 170.230 80.435 170.475 ;
        RECT -0.415 168.515 80.440 170.230 ;
        RECT -0.415 146.690 6.385 168.515 ;
        RECT 78.630 146.690 80.440 168.515 ;
        RECT -0.415 144.880 80.440 146.690 ;
      LAYER pwell ;
        RECT -0.290 140.685 80.290 144.565 ;
      LAYER nwell ;
        RECT 46.040 140.380 80.440 140.385 ;
        RECT -0.415 130.665 80.440 140.380 ;
      LAYER pwell ;
        RECT -0.215 129.315 40.245 130.355 ;
        RECT 66.910 129.315 80.290 130.355 ;
        RECT -0.215 125.135 80.290 129.315 ;
        RECT -0.215 103.550 5.735 125.135 ;
        RECT 77.865 103.550 80.290 125.135 ;
        RECT -0.215 101.965 80.290 103.550 ;
        RECT -0.215 96.255 5.215 101.965 ;
        RECT 39.385 100.820 80.290 101.965 ;
        RECT 52.880 99.520 80.290 100.820 ;
        RECT 76.770 97.985 80.290 99.520 ;
        RECT 39.385 96.255 80.290 97.985 ;
        RECT -0.215 95.975 80.290 96.255 ;
        RECT -0.215 95.260 45.840 95.975 ;
        RECT -0.215 94.955 46.590 95.260 ;
        RECT -0.215 92.935 9.300 94.955 ;
      LAYER nwell ;
        RECT 46.940 94.245 80.670 95.165 ;
        RECT 62.650 93.735 80.670 94.245 ;
        RECT -0.415 91.820 2.795 92.400 ;
        RECT -0.415 88.485 5.975 91.820 ;
        RECT -0.120 88.280 5.975 88.485 ;
        RECT -0.120 87.740 8.420 88.280 ;
        RECT -0.120 86.660 8.495 87.740 ;
        RECT -0.120 85.580 4.530 86.660 ;
        RECT 79.240 84.345 80.670 93.735 ;
        RECT 46.940 83.165 80.670 84.345 ;
        RECT -0.715 79.805 24.815 81.235 ;
        RECT -0.715 62.340 0.715 79.805 ;
        RECT 79.240 73.775 80.670 83.165 ;
        RECT 62.650 73.265 80.670 73.775 ;
        RECT 46.940 72.595 80.670 73.265 ;
        RECT 79.125 66.045 80.670 72.595 ;
        RECT 70.335 65.195 80.670 66.045 ;
        RECT -0.715 61.020 3.810 62.340 ;
        RECT -0.715 60.770 13.535 61.020 ;
        RECT -0.715 60.180 10.460 60.770 ;
        RECT -0.715 58.020 0.715 60.180 ;
        RECT -0.715 56.590 23.515 58.020 ;
        RECT 79.125 52.050 80.670 65.195 ;
        RECT 70.335 50.620 80.670 52.050 ;
        RECT 48.915 34.265 80.450 36.055 ;
        RECT 58.275 32.410 80.450 34.265 ;
        RECT 64.830 29.785 80.450 32.410 ;
        RECT 64.830 23.080 80.450 25.345 ;
        RECT 4.580 19.155 80.450 23.080 ;
        RECT -0.415 5.665 3.110 9.325 ;
      LAYER li1 ;
        RECT 0.000 178.645 80.000 199.705 ;
        RECT -0.085 170.090 80.105 178.645 ;
        RECT -0.115 145.215 80.105 170.090 ;
        RECT -0.115 145.155 80.000 145.215 ;
        RECT 0.000 144.435 80.000 145.155 ;
        RECT -0.160 140.815 80.160 144.435 ;
        RECT 0.000 140.150 80.000 140.815 ;
        RECT -0.115 140.055 80.000 140.150 ;
        RECT -0.115 131.275 80.085 140.055 ;
        RECT -0.085 130.995 80.085 131.275 ;
        RECT 0.000 130.225 80.000 130.995 ;
        RECT -0.085 130.220 80.160 130.225 ;
        RECT -0.115 96.105 80.160 130.220 ;
        RECT -0.115 95.895 80.000 96.105 ;
        RECT -0.085 94.580 80.000 95.895 ;
        RECT -0.085 93.065 80.085 94.580 ;
        RECT 0.000 92.070 80.085 93.065 ;
        RECT -0.085 88.815 80.085 92.070 ;
        RECT 0.000 80.605 80.085 88.815 ;
        RECT -0.085 57.220 80.085 80.605 ;
        RECT 0.000 51.250 80.085 57.220 ;
        RECT 0.000 35.725 80.000 51.250 ;
        RECT 0.000 30.115 80.120 35.725 ;
        RECT 0.000 25.015 80.000 30.115 ;
        RECT 0.000 19.485 80.120 25.015 ;
        RECT 0.000 8.995 80.000 19.485 ;
        RECT -0.085 5.995 80.000 8.995 ;
        RECT 0.000 0.230 80.000 5.995 ;
      LAYER met1 ;
        RECT 0.000 180.975 80.000 200.000 ;
        RECT 0.000 178.900 80.020 180.975 ;
        RECT 0.000 170.090 80.000 178.900 ;
        RECT -0.115 131.275 80.145 170.090 ;
        RECT 0.000 130.220 80.000 131.275 ;
        RECT -0.115 95.895 80.145 130.220 ;
        RECT 0.000 94.580 80.000 95.895 ;
        RECT 0.000 91.480 80.060 94.580 ;
        RECT -0.145 89.750 80.060 91.480 ;
        RECT 0.000 80.635 80.060 89.750 ;
        RECT -0.115 72.930 80.060 80.635 ;
        POLYGON 80.060 72.985 80.115 72.930 80.060 72.930 ;
        RECT -0.115 57.190 80.115 72.930 ;
        RECT 0.000 51.220 80.115 57.190 ;
        RECT 0.000 35.725 80.000 51.220 ;
        RECT 0.000 30.120 80.115 35.725 ;
        RECT 0.000 25.015 80.000 30.120 ;
        RECT 0.000 19.485 80.115 25.015 ;
        RECT 0.000 1.585 80.000 19.485 ;
        RECT 0.000 0.260 62.150 1.585 ;
        RECT 62.970 0.260 80.000 1.585 ;
      LAYER met2 ;
        RECT 0.210 178.150 79.915 200.000 ;
        RECT 0.210 6.705 79.435 178.150 ;
        RECT 0.210 5.630 22.075 6.705 ;
        RECT 0.210 4.755 12.475 5.630 ;
        RECT 0.210 0.250 3.095 4.755 ;
        RECT 3.885 0.250 5.140 4.755 ;
        RECT 5.930 1.830 12.475 4.755 ;
        RECT 6.670 0.250 12.475 1.830 ;
        RECT 13.295 2.600 22.075 5.630 ;
        RECT 13.295 0.250 16.030 2.600 ;
        RECT 16.850 0.250 22.075 2.600 ;
        RECT 22.895 5.370 79.435 6.705 ;
        RECT 22.895 4.350 44.965 5.370 ;
        RECT 22.895 2.985 28.210 4.350 ;
        RECT 22.895 0.250 26.320 2.985 ;
        RECT 27.140 0.250 28.210 2.985 ;
        RECT 29.030 3.620 44.965 4.350 ;
        RECT 29.030 2.545 31.535 3.620 ;
        RECT 29.030 0.250 30.470 2.545 ;
        RECT 31.290 0.250 31.535 2.545 ;
        RECT 32.355 3.370 44.965 3.620 ;
        RECT 32.355 1.830 38.110 3.370 ;
        RECT 32.355 0.250 35.180 1.830 ;
        RECT 36.000 0.250 38.110 1.830 ;
        RECT 38.930 0.250 44.965 3.370 ;
        RECT 45.785 2.550 79.435 5.370 ;
        RECT 45.785 1.475 67.995 2.550 ;
        RECT 45.785 0.825 66.555 1.475 ;
        RECT 45.785 0.250 49.575 0.825 ;
        RECT 50.395 0.250 66.555 0.825 ;
        RECT 67.375 0.250 67.995 1.475 ;
        RECT 69.205 2.335 79.435 2.550 ;
        RECT 69.205 0.250 76.000 2.335 ;
        RECT 77.200 1.495 79.435 2.335 ;
        RECT 77.200 1.465 78.425 1.495 ;
        RECT 77.200 0.250 77.330 1.465 ;
        RECT 78.150 0.250 78.425 1.465 ;
        RECT 79.185 0.250 79.435 1.495 ;
      LAYER met3 ;
        RECT 0.400 189.960 79.570 200.000 ;
        RECT 0.400 185.175 78.840 189.960 ;
        RECT 0.400 178.885 78.180 185.175 ;
        RECT 1.420 37.205 78.180 178.885 ;
        RECT 1.420 0.245 45.465 37.205 ;
        RECT 46.595 15.245 78.180 37.205 ;
        RECT 46.595 0.245 62.420 15.245 ;
        RECT 64.290 0.245 78.180 15.245 ;
      LAYER met4 ;
        RECT 25.950 175.385 65.830 200.000 ;
        RECT 1.345 121.650 78.165 175.385 ;
        RECT 1.345 121.640 9.410 121.650 ;
        RECT 1.345 120.410 8.170 121.640 ;
        RECT 12.900 120.805 78.165 121.650 ;
        RECT 1.345 119.355 7.115 120.410 ;
        RECT 10.200 119.610 78.165 120.805 ;
        RECT 1.345 106.185 1.600 119.355 ;
        RECT 5.870 118.555 7.115 119.355 ;
        RECT 8.970 118.555 78.165 119.610 ;
        RECT 5.870 106.985 78.165 118.555 ;
        RECT 5.870 106.185 7.430 106.985 ;
        RECT 1.345 104.160 7.430 106.185 ;
        RECT 10.255 104.160 78.165 106.985 ;
        RECT 1.345 95.400 78.165 104.160 ;
        RECT 1.860 69.635 67.630 95.400 ;
        RECT 1.345 68.935 78.165 69.635 ;
        RECT 7.260 63.685 60.545 68.935 ;
        RECT 1.345 63.085 78.165 63.685 ;
        RECT 70.245 57.835 71.175 63.085 ;
        RECT 1.345 57.135 78.165 57.835 ;
        RECT 3.010 56.505 46.690 57.135 ;
        RECT 36.840 52.725 38.360 56.505 ;
        RECT 3.010 51.745 46.690 52.725 ;
        RECT 52.545 48.465 54.065 51.245 ;
        RECT 3.010 47.335 46.690 47.965 ;
        RECT 1.345 46.635 78.165 47.335 ;
        RECT 14.310 41.185 55.305 46.635 ;
        RECT 1.345 40.585 78.165 41.185 ;
        RECT 5.835 36.335 66.910 40.585 ;
        RECT 1.345 35.735 78.165 36.335 ;
        RECT 22.670 31.485 23.450 35.735 ;
        RECT 1.345 30.885 78.165 31.485 ;
        RECT 19.730 25.435 21.130 30.885 ;
        RECT 1.345 24.835 78.165 25.435 ;
        RECT 7.830 19.385 71.335 24.835 ;
        RECT 1.345 18.785 78.165 19.385 ;
        RECT 24.990 14.535 51.170 18.785 ;
        RECT 1.345 13.935 78.165 14.535 ;
        RECT 34.635 8.485 69.865 13.935 ;
        RECT 1.345 7.885 78.165 8.485 ;
        RECT 11.550 1.635 76.410 7.885 ;
        RECT 1.345 0.535 78.165 1.635 ;
      LAYER met5 ;
        RECT 9.800 168.610 75.200 173.485 ;
        RECT 9.800 98.085 75.200 102.960 ;
  END
END sky130_fd_io__top_gpiov2

#--------EOF---------

MACRO sky130_fd_io__top_ground_hvc_wpad
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_ground_hvc_wpad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
  END VSSA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
  END VDDIO
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
  END VDDA
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
  END VDDIO_Q
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
  END VSSIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
  END VSWITCH
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
  END VSSIO_Q
  PIN G_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 6.200 104.175 68.800 166.625 ;
    END
  END G_PAD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 50.390 0.000 74.290 25.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 0.000 48.890 12.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 169.135 59.285 169.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 110.440 59.285 169.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 107.960 59.285 110.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 169.135 53.285 172.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.855 106.010 50.995 108.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 174.680 60.945 190.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.285 173.020 60.945 174.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 172.645 59.285 174.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.400 104.555 48.855 106.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 102.415 47.400 104.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.040 99.715 59.285 107.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.550 99.505 45.260 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 170.460 48.855 170.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 110.620 48.855 170.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 108.150 48.855 110.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.965 170.460 42.855 175.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 105.655 42.855 110.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.965 175.350 48.855 190.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 104.555 46.715 106.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.840 102.135 45.260 104.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.135 42.840 102.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 100.215 42.840 102.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 100.105 42.840 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.840 99.505 43.550 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 98.300 51.040 99.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.890 96.150 51.040 98.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 96.150 48.890 96.300 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.495 0.000 24.395 2.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.895 0.000 36.895 12.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.945 89.470 36.895 99.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.070 98.795 29.525 100.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 100.250 28.070 102.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 175.350 36.820 195.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.230 174.760 36.820 175.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.540 174.070 36.230 174.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.875 173.405 35.540 174.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.225 172.755 34.875 173.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.930 170.460 34.225 172.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 158.470 31.930 172.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 104.790 31.930 104.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.930 99.895 36.895 104.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 91.890 24.395 92.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 92.540 29.525 96.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.110 96.200 21.500 98.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.305 98.590 19.110 101.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 101.395 16.305 102.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.500 169.130 25.010 172.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 158.470 21.500 172.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 104.600 21.500 104.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.500 100.250 25.930 104.680 ;
    END
  END SRC_BDY_HVC
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895 0.000 27.895 0.535 ;
    END
  END OGC_HVC
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.495 0.000 24.395 32.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 0.000 74.290 90.185 ;
    END
  END G_CORE
  OBS
      LAYER li1 ;
        RECT 1.070 1.000 72.775 199.695 ;
      LAYER met1 ;
        RECT 0.185 0.970 73.620 199.725 ;
      LAYER met2 ;
        RECT 0.265 25.940 74.290 195.075 ;
        RECT 0.265 2.335 50.110 25.940 ;
        RECT 24.675 0.980 50.110 2.335 ;
      LAYER met3 ;
        RECT 0.240 174.950 25.530 195.100 ;
        RECT 37.220 190.440 74.290 195.100 ;
        RECT 37.220 190.420 49.375 190.440 ;
        RECT 0.240 174.470 35.140 174.950 ;
        RECT 0.240 173.805 34.475 174.470 ;
        RECT 37.220 174.360 37.565 190.420 ;
        RECT 49.255 174.950 49.375 190.420 ;
        RECT 0.240 173.190 33.825 173.805 ;
        RECT 36.630 173.670 37.565 174.360 ;
        RECT 0.240 158.070 15.100 173.190 ;
        RECT 21.900 173.040 25.530 173.190 ;
        RECT 32.330 173.155 33.825 173.190 ;
        RECT 25.410 168.730 25.530 173.040 ;
        RECT 35.940 173.005 37.565 173.670 ;
        RECT 35.275 172.355 37.565 173.005 ;
        RECT 34.625 170.060 37.565 172.355 ;
        RECT 43.255 171.010 49.375 174.950 ;
        RECT 61.345 172.620 74.290 190.440 ;
        RECT 59.685 172.245 74.290 172.620 ;
        RECT 21.900 158.070 25.530 168.730 ;
        RECT 32.330 158.070 42.455 170.060 ;
        RECT 0.240 111.020 42.455 158.070 ;
        RECT 49.255 168.735 49.375 171.010 ;
        RECT 53.685 169.685 74.290 172.245 ;
        RECT 0.240 105.260 37.490 111.020 ;
        RECT 49.255 108.550 52.885 168.735 ;
        RECT 51.395 108.360 52.885 108.550 ;
        RECT 0.240 105.080 25.530 105.260 ;
        RECT 37.295 105.255 37.490 105.260 ;
        RECT 43.255 106.410 48.455 107.750 ;
        RECT 43.255 105.255 44.860 106.410 ;
        RECT 0.240 104.200 15.100 105.080 ;
        RECT 37.295 104.955 44.860 105.255 ;
        RECT 0.240 102.600 21.100 104.200 ;
        RECT 26.330 102.790 31.530 104.390 ;
        RECT 0.240 100.995 15.100 102.600 ;
        RECT 16.705 101.795 21.100 102.600 ;
        RECT 0.240 98.190 15.905 100.995 ;
        RECT 19.510 99.850 21.100 101.795 ;
        RECT 28.470 100.650 31.530 102.790 ;
        RECT 19.510 98.990 27.670 99.850 ;
        RECT 21.900 98.395 27.670 98.990 ;
        RECT 29.925 99.495 31.530 100.650 ;
        RECT 37.295 102.685 42.440 104.955 ;
        RECT 49.255 104.155 50.640 105.610 ;
        RECT 29.925 98.395 31.545 99.495 ;
        RECT 0.240 95.800 18.710 98.190 ;
        RECT 21.900 97.055 31.545 98.395 ;
        RECT 21.900 95.800 23.345 97.055 ;
        RECT 0.240 91.490 23.345 95.800 ;
        RECT 29.925 92.140 31.545 97.055 ;
        RECT 24.795 91.490 31.545 92.140 ;
        RECT 0.240 89.070 31.545 91.490 ;
        RECT 37.295 97.900 37.490 102.685 ;
        RECT 47.800 102.015 50.640 104.155 ;
        RECT 45.660 101.735 50.640 102.015 ;
        RECT 43.240 100.615 50.640 101.735 ;
        RECT 43.950 99.905 44.150 100.615 ;
        RECT 45.660 99.905 50.640 100.615 ;
        RECT 59.685 99.315 74.290 169.685 ;
        RECT 37.295 96.700 48.490 97.900 ;
        RECT 37.295 95.750 37.490 96.700 ;
        RECT 51.440 95.750 74.290 99.315 ;
        RECT 37.295 90.585 74.290 95.750 ;
        RECT 37.295 89.070 49.990 90.585 ;
        RECT 0.240 32.915 49.990 89.070 ;
        RECT 24.795 12.825 49.990 32.915 ;
        RECT 24.795 12.380 25.495 12.825 ;
        RECT 37.295 12.780 49.990 12.825 ;
        RECT 37.295 12.380 37.490 12.780 ;
        RECT 49.290 12.380 49.990 12.780 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 168.225 75.000 174.185 ;
        RECT 0.000 102.575 4.600 168.225 ;
        RECT 70.400 102.575 75.000 168.225 ;
        RECT 0.000 96.585 75.000 102.575 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__top_ground_hvc_wpad

#--------EOF---------

MACRO sky130_fd_io__top_ground_lvc_wpad
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_ground_lvc_wpad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
  END VSSIO
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
  END VSSA
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
  END VSSIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
  END VCCHIB
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
  END VCCD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
  END VDDIO_Q
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
  END VSSD
  PIN G_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 9.315 100.140 65.955 167.570 ;
    END
  END G_PAD
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 0.000 20.495 1.485 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 0.000 74.700 3.660 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 0.000 44.440 0.325 ;
    END
  END BDY2_B2B
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 0.000 49.255 22.900 ;
    END
  END DRN_LVC2
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 0.000 36.880 20.220 ;
    END
  END DRN_LVC1
  PIN G_CORE
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 50.755 0.000 74.700 84.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 0.000 24.500 70.755 ;
    END
  END G_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210 0.000 27.700 0.170 ;
    END
  END OGC_LVC
  OBS
      LAYER li1 ;
        RECT 0.240 1.020 74.755 197.780 ;
      LAYER met1 ;
        RECT 0.120 0.450 74.785 197.840 ;
        RECT 0.120 0.000 25.930 0.450 ;
        RECT 27.980 0.000 74.785 0.450 ;
      LAYER met2 ;
        RECT 0.500 3.940 74.700 194.430 ;
        RECT 0.500 1.765 54.435 3.940 ;
        RECT 20.775 0.605 54.435 1.765 ;
        RECT 20.775 0.000 34.160 0.605 ;
        RECT 44.720 0.000 54.435 0.605 ;
      LAYER met3 ;
        RECT 0.500 84.865 74.700 189.515 ;
        RECT 0.500 71.155 50.355 84.865 ;
        RECT 24.900 23.300 50.355 71.155 ;
        RECT 24.900 20.620 37.980 23.300 ;
        RECT 24.900 17.790 25.600 20.620 ;
        RECT 37.280 17.790 37.980 20.620 ;
        RECT 49.655 17.790 50.355 23.300 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 169.170 75.000 172.185 ;
        RECT 0.000 98.540 7.715 169.170 ;
        RECT 67.555 98.540 75.000 169.170 ;
        RECT 0.000 94.585 75.000 98.540 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__top_ground_lvc_wpad

#--------EOF---------

MACRO sky130_fd_io__top_power_hvc_wpad
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_power_hvc_wpad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN P_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 11.330 97.700 63.670 173.100 ;
    END
  END P_PAD
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 61.110 0.000 74.290 190.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 107.960 59.285 190.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.805 107.815 59.140 107.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.660 107.665 58.990 107.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.510 107.515 58.840 107.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.360 107.365 58.690 107.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.210 107.215 58.540 107.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.060 107.065 58.390 107.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.910 106.915 58.240 107.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.760 106.765 58.090 106.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.610 106.615 57.940 106.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.460 106.465 57.790 106.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.310 106.315 57.640 106.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.160 106.165 57.490 106.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.010 106.015 57.340 106.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.860 105.865 57.190 106.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.710 105.715 57.040 105.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.560 105.565 56.890 105.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.410 105.415 56.740 105.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.260 105.265 56.590 105.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.110 105.115 56.440 105.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.960 104.965 56.290 105.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.810 104.815 56.140 104.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.660 104.665 55.990 104.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.510 104.515 55.840 104.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.360 104.365 55.690 104.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.210 104.215 55.540 104.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.060 104.065 55.390 104.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.910 103.915 55.240 104.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.760 103.765 55.090 103.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.610 103.615 54.940 103.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.460 103.465 54.790 103.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.310 103.315 54.640 103.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.160 103.165 54.490 103.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.010 103.015 54.340 103.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.860 102.865 54.190 103.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.710 102.715 54.040 102.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.560 102.565 53.890 102.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.410 102.415 53.740 102.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 102.315 53.640 102.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 102.165 53.490 102.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 102.015 53.340 102.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 101.865 53.190 102.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 101.715 53.040 101.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 101.565 52.890 101.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 101.415 52.740 101.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 101.265 52.590 101.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 101.115 52.440 101.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.965 52.290 101.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.815 52.140 100.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.665 51.990 100.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.515 51.840 100.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.365 51.690 100.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.215 51.540 100.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 100.165 51.490 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.210 100.015 51.340 100.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.060 99.865 51.190 100.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.910 98.300 51.040 99.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 108.150 48.855 190.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.385 108.055 48.760 108.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.290 107.905 48.610 108.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.140 107.755 48.460 107.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.990 107.605 48.310 107.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.840 107.455 48.160 107.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.690 107.305 48.010 107.455 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.540 107.155 47.860 107.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.390 107.005 47.710 107.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.240 106.855 47.560 107.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.090 106.705 47.410 106.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.940 106.555 47.260 106.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.790 106.405 47.110 106.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.640 106.255 46.960 106.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.490 106.105 46.810 106.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.340 105.955 46.660 106.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.190 105.805 46.510 105.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.040 105.655 46.360 105.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 105.585 46.290 105.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 105.435 46.140 105.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 105.285 45.990 105.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 105.135 45.840 105.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.985 45.690 105.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.835 45.540 104.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.685 45.390 104.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.535 45.240 104.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.385 45.090 104.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.235 44.940 104.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 104.085 44.790 104.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.935 44.640 104.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.785 44.490 103.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.635 44.340 103.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.485 44.190 103.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.335 44.040 103.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.185 43.890 103.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 103.035 43.740 103.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.885 43.590 103.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.735 43.440 102.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.585 43.290 102.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.435 43.140 102.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.285 42.990 102.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 0.000 42.840 102.285 ;
    END
  END DRN_HVC
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895 0.000 27.895 0.535 ;
    END
  END OGC_HVC
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495 0.000 24.395 36.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 0.000 74.290 50.000 ;
    END
  END P_CORE
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.670 36.115 56.915 39.665 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.260 39.665 56.845 39.735 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.190 39.735 56.775 39.805 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.120 39.805 56.705 39.875 ;
    END
    PORT
      LAYER met2 ;
        RECT 53.050 39.875 56.635 39.945 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.980 39.945 56.565 40.015 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.910 40.015 56.495 40.085 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.840 40.085 56.425 40.155 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.770 40.155 56.355 40.225 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.700 40.225 56.285 40.295 ;
    END
    PORT
      LAYER met2 ;
        RECT 52.630 40.295 56.230 40.350 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.090 0.000 14.120 195.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.945 0.000 36.895 99.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.425 99.895 36.745 100.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.275 100.045 36.595 100.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.125 100.195 36.445 100.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.975 100.345 36.295 100.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.825 100.495 36.145 100.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.675 100.645 35.995 100.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.525 100.795 35.845 100.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.375 100.945 35.695 101.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.225 101.095 35.545 101.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.075 101.245 35.395 101.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.925 101.395 35.245 101.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.775 101.545 35.095 101.695 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.625 101.695 34.945 101.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.475 101.845 34.795 101.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.325 101.995 34.645 102.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.175 102.145 34.495 102.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.025 102.295 34.400 102.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 175.350 36.820 200.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 175.260 36.730 175.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 175.110 36.580 175.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.960 36.430 175.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.810 36.280 174.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.660 36.130 174.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.510 35.980 174.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.360 35.830 174.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.210 35.680 174.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.060 35.530 174.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.910 35.380 174.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.760 35.230 173.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.610 35.080 173.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.460 34.930 173.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.310 34.780 173.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.160 34.630 173.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.010 34.480 173.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.860 34.330 173.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.710 34.180 172.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.560 34.030 172.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.410 33.880 172.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.260 33.730 172.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.110 33.580 172.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.960 33.430 172.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.810 33.280 171.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.660 33.130 171.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.510 32.980 171.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.360 32.830 171.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.210 32.680 171.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 171.060 32.530 171.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 170.910 32.380 171.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 170.760 32.230 170.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 170.610 32.080 170.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 102.390 31.930 170.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.895 92.390 30.160 92.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.820 92.465 30.085 92.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 92.540 29.525 96.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.045 96.655 29.375 96.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.895 96.805 29.225 96.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.745 96.955 29.075 97.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.595 97.105 28.925 97.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.445 97.255 28.775 97.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.295 97.405 28.625 97.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.145 97.555 28.475 97.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.995 97.705 28.325 97.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.845 97.855 28.175 98.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.695 98.005 28.025 98.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.545 98.155 27.875 98.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.395 98.305 27.725 98.455 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.245 98.455 27.575 98.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.095 98.605 27.425 98.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.945 98.755 27.275 98.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.795 98.905 27.125 99.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.645 99.055 26.975 99.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.495 99.205 26.825 99.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.345 99.355 26.675 99.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 99.505 26.525 99.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.045 99.655 26.375 99.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.895 99.805 26.225 99.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.745 99.955 26.075 100.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.595 100.105 25.925 100.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.445 100.255 25.775 100.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.295 100.405 25.625 100.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.145 100.555 25.475 100.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.995 100.705 25.325 100.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.845 100.855 25.175 101.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.695 101.005 25.025 101.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.545 101.155 24.875 101.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.395 101.305 24.725 101.455 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.245 101.455 24.575 101.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.095 101.605 24.425 101.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.945 101.755 24.275 101.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.795 101.905 24.125 102.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.645 102.055 23.980 102.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 172.640 25.010 200.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 172.580 24.950 172.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 172.430 24.800 172.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 172.280 24.650 172.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 172.130 24.500 172.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.980 24.350 172.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.830 24.200 171.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.680 24.050 171.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.530 23.900 171.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.380 23.750 171.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.230 23.600 171.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 171.080 23.450 171.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.930 23.300 171.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.780 23.150 170.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.630 23.000 170.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.480 22.850 170.630 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.330 22.700 170.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.180 22.550 170.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 170.030 22.400 170.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 169.880 22.250 170.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 169.730 22.100 169.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 169.580 21.950 169.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 169.430 21.800 169.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 169.280 21.650 169.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 102.200 21.500 169.280 ;
    END
  END SRC_BDY_HVC
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 75.000 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 75.000 7.385 ;
    END
  END VCCHIB
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 75.000 18.285 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 75.000 94.985 ;
    END
  END VDDIO
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 75.000 68.435 ;
    END
  END VDDIO_Q
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.835 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 75.000 56.735 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 75.000 46.135 ;
    END
  END VSSD
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 75.000 30.385 ;
    END
  END VSSIO
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 75.000 62.585 ;
    END
  END VSSIO_Q
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 75.000 35.235 ;
    END
  END VSWITCH
  OBS
      LAYER li1 ;
        RECT 1.070 1.000 72.775 199.695 ;
      LAYER met1 ;
        RECT 0.000 0.000 75.000 200.000 ;
      LAYER met2 ;
        RECT 0.000 195.355 75.000 200.000 ;
        RECT 0.000 46.980 0.725 195.355 ;
      LAYER met2 ;
        RECT 0.725 46.980 0.810 195.355 ;
      LAYER met2 ;
        RECT 0.000 46.940 0.730 46.980 ;
      LAYER met2 ;
        RECT 0.730 46.940 0.810 46.980 ;
      LAYER met2 ;
        RECT 0.000 46.900 0.770 46.940 ;
      LAYER met2 ;
        RECT 0.770 46.900 0.810 46.940 ;
      LAYER met2 ;
        RECT 0.000 36.970 0.810 46.900 ;
        RECT 0.000 2.170 0.725 36.970 ;
      LAYER met2 ;
        RECT 0.725 2.170 0.810 36.970 ;
      LAYER met2 ;
        RECT 0.000 0.000 0.215 2.170 ;
      LAYER met2 ;
        RECT 0.215 0.000 0.810 2.170 ;
        RECT 14.400 190.295 75.000 195.355 ;
        RECT 14.400 40.630 60.830 190.295 ;
        RECT 14.400 40.015 52.350 40.630 ;
        RECT 56.510 40.575 60.830 40.630 ;
        RECT 56.565 40.505 60.830 40.575 ;
        RECT 56.635 40.435 60.830 40.505 ;
        RECT 56.705 40.365 60.830 40.435 ;
        RECT 56.775 40.295 60.830 40.365 ;
        RECT 56.845 40.225 60.830 40.295 ;
        RECT 56.915 40.155 60.830 40.225 ;
        RECT 56.985 40.085 60.830 40.155 ;
        RECT 57.055 40.015 60.830 40.085 ;
        RECT 14.400 39.945 52.420 40.015 ;
        RECT 57.125 39.945 60.830 40.015 ;
        RECT 14.400 39.875 52.490 39.945 ;
        RECT 14.400 39.805 52.560 39.875 ;
        RECT 14.400 39.735 52.630 39.805 ;
        RECT 14.400 39.665 52.700 39.735 ;
        RECT 14.400 39.595 52.770 39.665 ;
        RECT 14.400 39.525 52.840 39.595 ;
        RECT 14.400 39.455 52.910 39.525 ;
        RECT 14.400 39.385 52.980 39.455 ;
        RECT 14.400 35.835 54.390 39.385 ;
        RECT 57.195 35.835 60.830 39.945 ;
        RECT 14.400 0.815 60.830 35.835 ;
        RECT 14.400 0.000 25.615 0.815 ;
        RECT 28.175 0.000 60.830 0.815 ;
        RECT 74.570 0.000 75.000 190.295 ;
      LAYER met3 ;
        RECT 0.000 185.105 2.760 200.000 ;
      LAYER met3 ;
        RECT 2.760 185.105 15.100 200.000 ;
      LAYER met3 ;
        RECT 0.000 184.955 2.850 185.105 ;
      LAYER met3 ;
        RECT 2.850 184.955 15.100 185.105 ;
      LAYER met3 ;
        RECT 0.000 184.805 3.000 184.955 ;
      LAYER met3 ;
        RECT 3.000 184.805 15.100 184.955 ;
      LAYER met3 ;
        RECT 0.000 184.655 3.150 184.805 ;
      LAYER met3 ;
        RECT 3.150 184.655 15.100 184.805 ;
      LAYER met3 ;
        RECT 0.000 184.505 3.300 184.655 ;
      LAYER met3 ;
        RECT 3.300 184.505 15.100 184.655 ;
      LAYER met3 ;
        RECT 0.000 184.355 3.450 184.505 ;
      LAYER met3 ;
        RECT 3.450 184.355 15.100 184.505 ;
      LAYER met3 ;
        RECT 0.000 184.205 3.600 184.355 ;
      LAYER met3 ;
        RECT 3.600 184.205 15.100 184.355 ;
      LAYER met3 ;
        RECT 0.000 184.055 3.750 184.205 ;
      LAYER met3 ;
        RECT 3.750 184.055 15.100 184.205 ;
      LAYER met3 ;
        RECT 0.000 183.905 3.900 184.055 ;
      LAYER met3 ;
        RECT 3.900 183.905 15.100 184.055 ;
      LAYER met3 ;
        RECT 0.000 183.755 4.050 183.905 ;
      LAYER met3 ;
        RECT 4.050 183.755 15.100 183.905 ;
      LAYER met3 ;
        RECT 0.000 183.605 4.200 183.755 ;
      LAYER met3 ;
        RECT 4.200 183.605 15.100 183.755 ;
      LAYER met3 ;
        RECT 0.000 183.455 4.350 183.605 ;
      LAYER met3 ;
        RECT 4.350 183.455 15.100 183.605 ;
      LAYER met3 ;
        RECT 0.000 183.305 4.500 183.455 ;
      LAYER met3 ;
        RECT 4.500 183.305 15.100 183.455 ;
      LAYER met3 ;
        RECT 0.000 183.155 4.650 183.305 ;
      LAYER met3 ;
        RECT 4.650 183.155 15.100 183.305 ;
      LAYER met3 ;
        RECT 0.000 183.005 4.800 183.155 ;
      LAYER met3 ;
        RECT 4.800 183.005 15.100 183.155 ;
      LAYER met3 ;
        RECT 0.000 182.855 4.950 183.005 ;
      LAYER met3 ;
        RECT 4.950 182.855 15.100 183.005 ;
      LAYER met3 ;
        RECT 0.000 182.705 5.100 182.855 ;
      LAYER met3 ;
        RECT 5.100 182.705 15.100 182.855 ;
      LAYER met3 ;
        RECT 0.000 182.555 5.250 182.705 ;
      LAYER met3 ;
        RECT 5.250 182.555 15.100 182.705 ;
      LAYER met3 ;
        RECT 0.000 182.405 5.400 182.555 ;
      LAYER met3 ;
        RECT 5.400 182.405 15.100 182.555 ;
      LAYER met3 ;
        RECT 0.000 182.255 5.550 182.405 ;
      LAYER met3 ;
        RECT 5.550 182.255 15.100 182.405 ;
      LAYER met3 ;
        RECT 0.000 182.105 5.700 182.255 ;
      LAYER met3 ;
        RECT 5.700 182.105 15.100 182.255 ;
      LAYER met3 ;
        RECT 0.000 181.955 5.850 182.105 ;
      LAYER met3 ;
        RECT 5.850 181.955 15.100 182.105 ;
      LAYER met3 ;
        RECT 0.000 181.805 6.000 181.955 ;
      LAYER met3 ;
        RECT 6.000 181.805 15.100 181.955 ;
      LAYER met3 ;
        RECT 0.000 181.655 6.150 181.805 ;
      LAYER met3 ;
        RECT 6.150 181.655 15.100 181.805 ;
      LAYER met3 ;
        RECT 0.000 181.505 6.300 181.655 ;
      LAYER met3 ;
        RECT 6.300 181.505 15.100 181.655 ;
      LAYER met3 ;
        RECT 0.000 181.355 6.450 181.505 ;
      LAYER met3 ;
        RECT 6.450 181.355 15.100 181.505 ;
      LAYER met3 ;
        RECT 0.000 181.205 6.600 181.355 ;
      LAYER met3 ;
        RECT 6.600 181.205 15.100 181.355 ;
      LAYER met3 ;
        RECT 0.000 181.055 6.750 181.205 ;
      LAYER met3 ;
        RECT 6.750 181.055 15.100 181.205 ;
      LAYER met3 ;
        RECT 0.000 180.905 6.900 181.055 ;
      LAYER met3 ;
        RECT 6.900 180.905 15.100 181.055 ;
      LAYER met3 ;
        RECT 0.000 180.755 7.050 180.905 ;
      LAYER met3 ;
        RECT 7.050 180.755 15.100 180.905 ;
      LAYER met3 ;
        RECT 0.000 180.605 7.200 180.755 ;
      LAYER met3 ;
        RECT 7.200 180.605 15.100 180.755 ;
      LAYER met3 ;
        RECT 0.000 180.455 7.350 180.605 ;
      LAYER met3 ;
        RECT 7.350 180.455 15.100 180.605 ;
      LAYER met3 ;
        RECT 0.000 180.305 7.500 180.455 ;
      LAYER met3 ;
        RECT 7.500 180.305 15.100 180.455 ;
      LAYER met3 ;
        RECT 0.000 180.155 7.650 180.305 ;
      LAYER met3 ;
        RECT 7.650 180.155 15.100 180.305 ;
      LAYER met3 ;
        RECT 0.000 180.005 7.800 180.155 ;
      LAYER met3 ;
        RECT 7.800 180.005 15.100 180.155 ;
      LAYER met3 ;
        RECT 0.000 179.855 7.950 180.005 ;
      LAYER met3 ;
        RECT 7.950 179.855 15.100 180.005 ;
      LAYER met3 ;
        RECT 0.000 179.705 8.100 179.855 ;
      LAYER met3 ;
        RECT 8.100 179.705 15.100 179.855 ;
      LAYER met3 ;
        RECT 0.000 179.555 8.250 179.705 ;
      LAYER met3 ;
        RECT 8.250 179.555 15.100 179.705 ;
      LAYER met3 ;
        RECT 0.000 179.405 8.400 179.555 ;
      LAYER met3 ;
        RECT 8.400 179.405 15.100 179.555 ;
      LAYER met3 ;
        RECT 0.000 179.255 8.550 179.405 ;
      LAYER met3 ;
        RECT 8.550 179.255 15.100 179.405 ;
      LAYER met3 ;
        RECT 0.000 179.105 8.700 179.255 ;
      LAYER met3 ;
        RECT 8.700 179.105 15.100 179.255 ;
      LAYER met3 ;
        RECT 0.000 178.955 8.850 179.105 ;
      LAYER met3 ;
        RECT 8.850 178.955 15.100 179.105 ;
      LAYER met3 ;
        RECT 0.000 178.805 9.000 178.955 ;
      LAYER met3 ;
        RECT 9.000 178.805 15.100 178.955 ;
      LAYER met3 ;
        RECT 0.000 178.655 9.150 178.805 ;
      LAYER met3 ;
        RECT 9.150 178.655 15.100 178.805 ;
      LAYER met3 ;
        RECT 0.000 178.505 9.300 178.655 ;
      LAYER met3 ;
        RECT 9.300 178.505 15.100 178.655 ;
      LAYER met3 ;
        RECT 0.000 178.355 9.450 178.505 ;
      LAYER met3 ;
        RECT 9.450 178.355 15.100 178.505 ;
      LAYER met3 ;
        RECT 0.000 178.205 9.600 178.355 ;
      LAYER met3 ;
        RECT 9.600 178.205 15.100 178.355 ;
      LAYER met3 ;
        RECT 0.000 178.055 9.750 178.205 ;
      LAYER met3 ;
        RECT 9.750 178.055 15.100 178.205 ;
      LAYER met3 ;
        RECT 0.000 177.905 9.900 178.055 ;
      LAYER met3 ;
        RECT 9.900 177.905 15.100 178.055 ;
      LAYER met3 ;
        RECT 0.000 177.755 10.050 177.905 ;
      LAYER met3 ;
        RECT 10.050 177.755 15.100 177.905 ;
      LAYER met3 ;
        RECT 0.000 177.605 10.200 177.755 ;
      LAYER met3 ;
        RECT 10.200 177.605 15.100 177.755 ;
      LAYER met3 ;
        RECT 0.000 177.455 10.350 177.605 ;
      LAYER met3 ;
        RECT 10.350 177.455 15.100 177.605 ;
      LAYER met3 ;
        RECT 0.000 177.305 10.500 177.455 ;
      LAYER met3 ;
        RECT 10.500 177.305 15.100 177.455 ;
      LAYER met3 ;
        RECT 0.000 177.155 10.650 177.305 ;
      LAYER met3 ;
        RECT 10.650 177.155 15.100 177.305 ;
      LAYER met3 ;
        RECT 0.000 177.005 10.800 177.155 ;
      LAYER met3 ;
        RECT 10.800 177.005 15.100 177.155 ;
      LAYER met3 ;
        RECT 0.000 176.855 10.950 177.005 ;
      LAYER met3 ;
        RECT 10.950 176.855 15.100 177.005 ;
      LAYER met3 ;
        RECT 0.000 176.705 11.100 176.855 ;
      LAYER met3 ;
        RECT 11.100 176.705 15.100 176.855 ;
      LAYER met3 ;
        RECT 0.000 176.555 11.250 176.705 ;
      LAYER met3 ;
        RECT 11.250 176.555 15.100 176.705 ;
      LAYER met3 ;
        RECT 0.000 176.405 11.400 176.555 ;
      LAYER met3 ;
        RECT 11.400 176.405 15.100 176.555 ;
      LAYER met3 ;
        RECT 0.000 176.255 11.550 176.405 ;
      LAYER met3 ;
        RECT 11.550 176.255 15.100 176.405 ;
      LAYER met3 ;
        RECT 0.000 176.105 11.700 176.255 ;
      LAYER met3 ;
        RECT 11.700 176.105 15.100 176.255 ;
      LAYER met3 ;
        RECT 0.000 175.955 11.850 176.105 ;
      LAYER met3 ;
        RECT 11.850 175.955 15.100 176.105 ;
      LAYER met3 ;
        RECT 0.000 175.805 12.000 175.955 ;
      LAYER met3 ;
        RECT 12.000 175.805 15.100 175.955 ;
      LAYER met3 ;
        RECT 0.000 175.655 12.150 175.805 ;
      LAYER met3 ;
        RECT 12.150 175.655 15.100 175.805 ;
      LAYER met3 ;
        RECT 0.000 175.505 12.300 175.655 ;
      LAYER met3 ;
        RECT 12.300 175.505 15.100 175.655 ;
      LAYER met3 ;
        RECT 0.000 175.355 12.450 175.505 ;
      LAYER met3 ;
        RECT 12.450 175.355 15.100 175.505 ;
      LAYER met3 ;
        RECT 0.000 175.205 12.600 175.355 ;
      LAYER met3 ;
        RECT 12.600 175.205 15.100 175.355 ;
      LAYER met3 ;
        RECT 0.000 175.055 12.750 175.205 ;
      LAYER met3 ;
        RECT 12.750 175.055 15.100 175.205 ;
      LAYER met3 ;
        RECT 0.000 174.905 12.900 175.055 ;
      LAYER met3 ;
        RECT 12.900 174.905 15.100 175.055 ;
      LAYER met3 ;
        RECT 0.000 174.755 13.050 174.905 ;
      LAYER met3 ;
        RECT 13.050 174.755 15.100 174.905 ;
      LAYER met3 ;
        RECT 0.000 174.605 13.200 174.755 ;
      LAYER met3 ;
        RECT 13.200 174.605 15.100 174.755 ;
      LAYER met3 ;
        RECT 0.000 174.455 13.350 174.605 ;
      LAYER met3 ;
        RECT 13.350 174.455 15.100 174.605 ;
      LAYER met3 ;
        RECT 0.000 174.305 13.500 174.455 ;
      LAYER met3 ;
        RECT 13.500 174.305 15.100 174.455 ;
      LAYER met3 ;
        RECT 0.000 174.155 13.650 174.305 ;
      LAYER met3 ;
        RECT 13.650 174.155 15.100 174.305 ;
      LAYER met3 ;
        RECT 0.000 174.005 13.800 174.155 ;
      LAYER met3 ;
        RECT 13.800 174.005 15.100 174.155 ;
      LAYER met3 ;
        RECT 0.000 173.855 13.950 174.005 ;
      LAYER met3 ;
        RECT 13.950 173.855 15.100 174.005 ;
      LAYER met3 ;
        RECT 0.000 173.705 14.100 173.855 ;
      LAYER met3 ;
        RECT 14.100 173.705 15.100 173.855 ;
      LAYER met3 ;
        RECT 0.000 173.555 14.250 173.705 ;
      LAYER met3 ;
        RECT 14.250 173.555 15.100 173.705 ;
      LAYER met3 ;
        RECT 0.000 173.455 2.760 173.555 ;
      LAYER met3 ;
        RECT 2.760 173.455 15.100 173.555 ;
      LAYER met3 ;
        RECT 0.000 46.630 0.195 173.455 ;
      LAYER met3 ;
        RECT 0.195 101.800 15.100 173.455 ;
        RECT 25.410 172.240 25.530 200.000 ;
        RECT 37.220 190.440 75.000 200.000 ;
        RECT 37.220 190.420 52.885 190.440 ;
        RECT 37.220 174.950 42.455 190.420 ;
        RECT 37.130 174.860 42.455 174.950 ;
        RECT 36.980 174.710 42.455 174.860 ;
        RECT 36.830 174.560 42.455 174.710 ;
        RECT 36.680 174.410 42.455 174.560 ;
        RECT 36.530 174.260 42.455 174.410 ;
        RECT 36.380 174.110 42.455 174.260 ;
        RECT 36.230 173.960 42.455 174.110 ;
        RECT 36.080 173.810 42.455 173.960 ;
        RECT 35.930 173.660 42.455 173.810 ;
        RECT 35.780 173.510 42.455 173.660 ;
        RECT 35.630 173.360 42.455 173.510 ;
        RECT 35.480 173.210 42.455 173.360 ;
        RECT 35.330 173.060 42.455 173.210 ;
        RECT 35.180 172.910 42.455 173.060 ;
        RECT 35.030 172.760 42.455 172.910 ;
        RECT 34.880 172.610 42.455 172.760 ;
        RECT 34.730 172.460 42.455 172.610 ;
        RECT 34.580 172.310 42.455 172.460 ;
        RECT 25.350 172.180 25.530 172.240 ;
        RECT 25.200 172.030 25.530 172.180 ;
        RECT 34.430 172.160 42.455 172.310 ;
        RECT 25.050 171.880 25.530 172.030 ;
        RECT 34.280 172.010 42.455 172.160 ;
        RECT 24.900 171.730 25.530 171.880 ;
        RECT 34.130 171.860 42.455 172.010 ;
        RECT 24.750 171.580 25.530 171.730 ;
        RECT 33.980 171.710 42.455 171.860 ;
        RECT 24.600 171.430 25.530 171.580 ;
        RECT 33.830 171.560 42.455 171.710 ;
        RECT 24.450 171.280 25.530 171.430 ;
        RECT 33.680 171.410 42.455 171.560 ;
        RECT 24.300 171.130 25.530 171.280 ;
        RECT 33.530 171.260 42.455 171.410 ;
        RECT 24.150 170.980 25.530 171.130 ;
        RECT 33.380 171.110 42.455 171.260 ;
        RECT 24.000 170.830 25.530 170.980 ;
        RECT 33.230 170.960 42.455 171.110 ;
        RECT 23.850 170.680 25.530 170.830 ;
        RECT 33.080 170.810 42.455 170.960 ;
        RECT 23.700 170.530 25.530 170.680 ;
        RECT 32.930 170.660 42.455 170.810 ;
        RECT 23.550 170.380 25.530 170.530 ;
        RECT 32.780 170.510 42.455 170.660 ;
        RECT 23.400 170.230 25.530 170.380 ;
        RECT 32.630 170.360 42.455 170.510 ;
        RECT 23.250 170.080 25.530 170.230 ;
        RECT 32.480 170.210 42.455 170.360 ;
        RECT 23.100 169.930 25.530 170.080 ;
        RECT 22.950 169.780 25.530 169.930 ;
        RECT 22.800 169.630 25.530 169.780 ;
        RECT 22.650 169.480 25.530 169.630 ;
        RECT 22.500 169.330 25.530 169.480 ;
        RECT 22.350 169.180 25.530 169.330 ;
        RECT 22.200 169.030 25.530 169.180 ;
        RECT 22.050 168.880 25.530 169.030 ;
        RECT 21.900 102.600 25.530 168.880 ;
        RECT 32.330 108.550 42.455 170.210 ;
        RECT 32.330 108.455 39.985 108.550 ;
        RECT 32.330 108.305 39.890 108.455 ;
        RECT 49.255 108.360 52.885 190.420 ;
        RECT 32.330 108.155 39.740 108.305 ;
        RECT 49.255 108.215 50.405 108.360 ;
        RECT 32.330 108.005 39.590 108.155 ;
        RECT 49.255 108.065 50.260 108.215 ;
        RECT 32.330 107.855 39.440 108.005 ;
        RECT 49.255 107.915 50.110 108.065 ;
        RECT 32.330 107.705 39.290 107.855 ;
        RECT 49.255 107.765 49.960 107.915 ;
        RECT 49.255 107.750 49.810 107.765 ;
        RECT 32.330 107.555 39.140 107.705 ;
        RECT 49.160 107.655 49.810 107.750 ;
        RECT 49.010 107.615 49.810 107.655 ;
        RECT 32.330 107.405 38.990 107.555 ;
        RECT 49.010 107.505 49.660 107.615 ;
        RECT 59.685 107.560 75.000 190.440 ;
        RECT 48.860 107.465 49.660 107.505 ;
        RECT 32.330 107.255 38.840 107.405 ;
        RECT 48.860 107.355 49.510 107.465 ;
        RECT 59.540 107.415 75.000 107.560 ;
        RECT 48.710 107.315 49.510 107.355 ;
        RECT 32.330 107.105 38.690 107.255 ;
        RECT 48.710 107.205 49.360 107.315 ;
        RECT 59.390 107.265 75.000 107.415 ;
        RECT 48.560 107.165 49.360 107.205 ;
        RECT 32.330 106.955 38.540 107.105 ;
        RECT 48.560 107.055 49.210 107.165 ;
        RECT 59.240 107.115 75.000 107.265 ;
        RECT 48.410 107.015 49.210 107.055 ;
        RECT 32.330 106.805 38.390 106.955 ;
        RECT 48.410 106.905 49.060 107.015 ;
        RECT 59.090 106.965 75.000 107.115 ;
        RECT 48.260 106.865 49.060 106.905 ;
        RECT 32.330 106.655 38.240 106.805 ;
        RECT 48.260 106.755 48.910 106.865 ;
        RECT 58.940 106.815 75.000 106.965 ;
        RECT 48.110 106.715 48.910 106.755 ;
        RECT 32.330 106.505 38.090 106.655 ;
        RECT 48.110 106.605 48.760 106.715 ;
        RECT 58.790 106.665 75.000 106.815 ;
        RECT 47.960 106.565 48.760 106.605 ;
        RECT 32.330 106.355 37.940 106.505 ;
        RECT 47.960 106.455 48.610 106.565 ;
        RECT 58.640 106.515 75.000 106.665 ;
        RECT 47.810 106.415 48.610 106.455 ;
        RECT 32.330 106.205 37.790 106.355 ;
        RECT 47.810 106.305 48.460 106.415 ;
        RECT 58.490 106.365 75.000 106.515 ;
        RECT 47.660 106.265 48.460 106.305 ;
        RECT 32.330 106.055 37.640 106.205 ;
        RECT 47.660 106.155 48.310 106.265 ;
        RECT 58.340 106.215 75.000 106.365 ;
        RECT 47.510 106.115 48.310 106.155 ;
        RECT 32.330 102.790 37.490 106.055 ;
        RECT 47.510 106.005 48.160 106.115 ;
        RECT 58.190 106.065 75.000 106.215 ;
        RECT 47.360 105.965 48.160 106.005 ;
        RECT 47.360 105.855 48.010 105.965 ;
        RECT 58.040 105.915 75.000 106.065 ;
        RECT 47.210 105.815 48.010 105.855 ;
        RECT 47.210 105.705 47.860 105.815 ;
        RECT 57.890 105.765 75.000 105.915 ;
        RECT 47.060 105.665 47.860 105.705 ;
        RECT 47.060 105.555 47.710 105.665 ;
        RECT 57.740 105.615 75.000 105.765 ;
        RECT 46.910 105.515 47.710 105.555 ;
        RECT 46.910 105.405 47.560 105.515 ;
        RECT 57.590 105.465 75.000 105.615 ;
        RECT 46.760 105.365 47.560 105.405 ;
        RECT 46.760 105.255 47.410 105.365 ;
        RECT 57.440 105.315 75.000 105.465 ;
        RECT 46.690 105.215 47.410 105.255 ;
        RECT 46.690 105.185 47.260 105.215 ;
        RECT 46.540 105.065 47.260 105.185 ;
        RECT 57.290 105.165 75.000 105.315 ;
        RECT 46.540 105.035 47.110 105.065 ;
        RECT 46.390 104.915 47.110 105.035 ;
        RECT 57.140 105.015 75.000 105.165 ;
        RECT 46.390 104.885 46.960 104.915 ;
        RECT 46.240 104.765 46.960 104.885 ;
        RECT 56.990 104.865 75.000 105.015 ;
        RECT 46.240 104.735 46.810 104.765 ;
        RECT 46.090 104.615 46.810 104.735 ;
        RECT 56.840 104.715 75.000 104.865 ;
        RECT 46.090 104.585 46.660 104.615 ;
        RECT 45.940 104.465 46.660 104.585 ;
        RECT 56.690 104.565 75.000 104.715 ;
        RECT 45.940 104.435 46.510 104.465 ;
        RECT 45.790 104.315 46.510 104.435 ;
        RECT 56.540 104.415 75.000 104.565 ;
        RECT 45.790 104.285 46.360 104.315 ;
        RECT 45.640 104.165 46.360 104.285 ;
        RECT 56.390 104.265 75.000 104.415 ;
        RECT 45.640 104.135 46.210 104.165 ;
        RECT 45.490 104.015 46.210 104.135 ;
        RECT 56.240 104.115 75.000 104.265 ;
        RECT 45.490 103.985 46.060 104.015 ;
        RECT 45.340 103.865 46.060 103.985 ;
        RECT 56.090 103.965 75.000 104.115 ;
        RECT 45.340 103.835 45.910 103.865 ;
        RECT 45.190 103.715 45.910 103.835 ;
        RECT 55.940 103.815 75.000 103.965 ;
        RECT 45.190 103.685 45.760 103.715 ;
        RECT 45.040 103.565 45.760 103.685 ;
        RECT 55.790 103.665 75.000 103.815 ;
        RECT 45.040 103.535 45.610 103.565 ;
        RECT 44.890 103.415 45.610 103.535 ;
        RECT 55.640 103.515 75.000 103.665 ;
        RECT 44.890 103.385 45.460 103.415 ;
        RECT 44.740 103.265 45.460 103.385 ;
        RECT 55.490 103.365 75.000 103.515 ;
        RECT 44.740 103.235 45.310 103.265 ;
        RECT 44.590 103.115 45.310 103.235 ;
        RECT 55.340 103.215 75.000 103.365 ;
        RECT 44.590 103.085 45.160 103.115 ;
        RECT 44.440 102.965 45.160 103.085 ;
        RECT 55.190 103.065 75.000 103.215 ;
        RECT 44.440 102.935 45.010 102.965 ;
        RECT 34.800 102.695 37.490 102.790 ;
        RECT 44.290 102.815 45.010 102.935 ;
        RECT 55.040 102.915 75.000 103.065 ;
        RECT 44.290 102.785 44.860 102.815 ;
        RECT 24.380 102.455 25.530 102.600 ;
        RECT 34.895 102.545 37.490 102.695 ;
        RECT 44.140 102.635 44.860 102.785 ;
        RECT 54.890 102.765 75.000 102.915 ;
        RECT 24.525 102.305 25.530 102.455 ;
        RECT 35.045 102.395 37.490 102.545 ;
        RECT 43.990 102.485 44.860 102.635 ;
        RECT 54.740 102.615 75.000 102.765 ;
        RECT 24.675 102.155 25.530 102.305 ;
        RECT 35.195 102.245 37.490 102.395 ;
        RECT 43.840 102.335 44.860 102.485 ;
        RECT 54.590 102.465 75.000 102.615 ;
        RECT 24.825 102.005 25.530 102.155 ;
        RECT 35.345 102.095 37.490 102.245 ;
        RECT 43.690 102.185 44.860 102.335 ;
        RECT 54.440 102.315 75.000 102.465 ;
        RECT 24.975 101.990 25.530 102.005 ;
        RECT 24.975 101.895 25.625 101.990 ;
        RECT 35.495 101.945 37.490 102.095 ;
        RECT 43.540 102.035 44.860 102.185 ;
        RECT 54.290 102.165 75.000 102.315 ;
        RECT 24.975 101.855 25.775 101.895 ;
        RECT 0.195 101.655 15.245 101.800 ;
        RECT 25.125 101.745 25.775 101.855 ;
        RECT 35.645 101.795 37.490 101.945 ;
        RECT 43.390 101.885 44.860 102.035 ;
        RECT 54.140 102.015 75.000 102.165 ;
        RECT 54.040 101.915 75.000 102.015 ;
        RECT 25.125 101.705 25.925 101.745 ;
        RECT 0.195 101.505 15.395 101.655 ;
        RECT 25.275 101.595 25.925 101.705 ;
        RECT 35.795 101.645 37.490 101.795 ;
        RECT 25.275 101.555 26.075 101.595 ;
        RECT 0.195 101.355 15.545 101.505 ;
        RECT 25.425 101.445 26.075 101.555 ;
        RECT 35.945 101.495 37.490 101.645 ;
        RECT 25.425 101.405 26.225 101.445 ;
        RECT 0.195 101.205 15.695 101.355 ;
        RECT 25.575 101.295 26.225 101.405 ;
        RECT 36.095 101.345 37.490 101.495 ;
        RECT 25.575 101.255 26.375 101.295 ;
        RECT 0.195 101.055 15.845 101.205 ;
        RECT 25.725 101.145 26.375 101.255 ;
        RECT 36.245 101.195 37.490 101.345 ;
        RECT 25.725 101.105 26.525 101.145 ;
        RECT 0.195 100.905 15.995 101.055 ;
        RECT 25.875 100.995 26.525 101.105 ;
        RECT 36.395 101.045 37.490 101.195 ;
        RECT 25.875 100.955 26.675 100.995 ;
        RECT 0.195 100.755 16.145 100.905 ;
        RECT 26.025 100.845 26.675 100.955 ;
        RECT 36.545 100.895 37.490 101.045 ;
        RECT 26.025 100.805 26.825 100.845 ;
        RECT 0.195 100.605 16.295 100.755 ;
        RECT 26.175 100.695 26.825 100.805 ;
        RECT 36.695 100.745 37.490 100.895 ;
        RECT 26.175 100.655 26.975 100.695 ;
        RECT 0.195 100.455 16.445 100.605 ;
        RECT 26.325 100.545 26.975 100.655 ;
        RECT 36.845 100.595 37.490 100.745 ;
        RECT 26.325 100.505 27.125 100.545 ;
        RECT 0.195 100.305 16.595 100.455 ;
        RECT 26.475 100.395 27.125 100.505 ;
        RECT 36.995 100.445 37.490 100.595 ;
        RECT 26.475 100.355 27.275 100.395 ;
        RECT 0.195 100.155 16.745 100.305 ;
        RECT 26.625 100.245 27.275 100.355 ;
        RECT 37.145 100.265 37.490 100.445 ;
        RECT 26.625 100.205 27.425 100.245 ;
        RECT 0.195 100.005 16.895 100.155 ;
        RECT 26.775 100.095 27.425 100.205 ;
        RECT 26.775 100.055 27.575 100.095 ;
        RECT 0.195 99.855 17.045 100.005 ;
        RECT 26.925 99.945 27.575 100.055 ;
        RECT 26.925 99.905 27.725 99.945 ;
        RECT 0.195 99.705 17.195 99.855 ;
        RECT 27.075 99.795 27.725 99.905 ;
        RECT 27.075 99.755 27.875 99.795 ;
        RECT 0.195 99.555 17.345 99.705 ;
        RECT 27.225 99.645 27.875 99.755 ;
        RECT 27.225 99.605 28.025 99.645 ;
        RECT 0.195 99.405 17.495 99.555 ;
        RECT 27.375 99.495 28.025 99.605 ;
        RECT 27.375 99.455 31.545 99.495 ;
        RECT 0.195 99.255 17.645 99.405 ;
        RECT 27.525 99.305 31.545 99.455 ;
        RECT 0.195 99.105 17.795 99.255 ;
        RECT 27.675 99.155 31.545 99.305 ;
        RECT 0.195 98.955 17.945 99.105 ;
        RECT 27.825 99.005 31.545 99.155 ;
        RECT 0.195 98.805 18.095 98.955 ;
        RECT 27.975 98.855 31.545 99.005 ;
        RECT 0.195 98.655 18.245 98.805 ;
        RECT 28.125 98.705 31.545 98.855 ;
        RECT 0.195 98.505 18.395 98.655 ;
        RECT 28.275 98.555 31.545 98.705 ;
        RECT 0.195 98.355 18.545 98.505 ;
        RECT 28.425 98.405 31.545 98.555 ;
        RECT 0.195 98.205 18.695 98.355 ;
        RECT 28.575 98.255 31.545 98.405 ;
        RECT 0.195 98.055 18.845 98.205 ;
        RECT 28.725 98.105 31.545 98.255 ;
        RECT 0.195 97.905 18.995 98.055 ;
        RECT 28.875 97.955 31.545 98.105 ;
        RECT 0.195 97.755 19.145 97.905 ;
        RECT 29.025 97.805 31.545 97.955 ;
        RECT 0.195 97.605 19.295 97.755 ;
        RECT 29.175 97.655 31.545 97.805 ;
        RECT 0.195 97.455 19.445 97.605 ;
        RECT 29.325 97.505 31.545 97.655 ;
        RECT 0.195 97.305 19.595 97.455 ;
        RECT 29.475 97.355 31.545 97.505 ;
        RECT 0.195 97.155 19.745 97.305 ;
        RECT 29.625 97.205 31.545 97.355 ;
        RECT 0.195 97.005 19.895 97.155 ;
        RECT 29.775 97.055 31.545 97.205 ;
        RECT 0.195 96.855 20.045 97.005 ;
        RECT 0.195 96.705 20.195 96.855 ;
        RECT 0.195 96.555 20.345 96.705 ;
        RECT 0.195 96.405 20.495 96.555 ;
        RECT 0.195 96.255 20.645 96.405 ;
        RECT 0.195 92.140 23.345 96.255 ;
        RECT 29.925 92.940 31.545 97.055 ;
        RECT 30.485 92.865 31.545 92.940 ;
        RECT 0.195 92.065 23.420 92.140 ;
        RECT 0.195 91.990 23.495 92.065 ;
        RECT 30.560 91.990 31.545 92.865 ;
        RECT 0.195 46.630 31.545 91.990 ;
      LAYER met3 ;
        RECT 0.000 46.480 0.260 46.630 ;
      LAYER met3 ;
        RECT 0.260 46.480 31.545 46.630 ;
      LAYER met3 ;
        RECT 0.000 46.330 0.410 46.480 ;
      LAYER met3 ;
        RECT 0.410 46.330 31.545 46.480 ;
      LAYER met3 ;
        RECT 0.000 46.220 0.560 46.330 ;
      LAYER met3 ;
        RECT 0.560 46.220 31.545 46.330 ;
      LAYER met3 ;
        RECT 0.000 36.635 0.810 46.220 ;
      LAYER met3 ;
        RECT 0.810 36.910 31.545 46.220 ;
      LAYER met3 ;
        RECT 0.000 0.000 0.195 36.635 ;
      LAYER met3 ;
        RECT 24.795 0.000 31.545 36.910 ;
        RECT 37.295 0.000 37.490 100.265 ;
        RECT 43.240 100.565 44.860 101.885 ;
        RECT 53.890 101.765 75.000 101.915 ;
        RECT 53.740 101.615 75.000 101.765 ;
        RECT 53.590 101.465 75.000 101.615 ;
        RECT 53.440 101.315 75.000 101.465 ;
        RECT 53.290 101.165 75.000 101.315 ;
        RECT 53.140 101.015 75.000 101.165 ;
        RECT 52.990 100.865 75.000 101.015 ;
        RECT 52.840 100.715 75.000 100.865 ;
        RECT 52.690 100.565 75.000 100.715 ;
        RECT 43.240 100.415 44.810 100.565 ;
        RECT 52.540 100.415 75.000 100.565 ;
        RECT 43.240 100.265 44.660 100.415 ;
        RECT 52.390 100.265 75.000 100.415 ;
        RECT 43.240 97.900 44.510 100.265 ;
        RECT 52.240 100.115 75.000 100.265 ;
        RECT 52.090 99.965 75.000 100.115 ;
        RECT 51.940 99.815 75.000 99.965 ;
        RECT 51.890 99.765 75.000 99.815 ;
        RECT 51.740 99.615 75.000 99.765 ;
        RECT 51.590 99.465 75.000 99.615 ;
        RECT 51.440 97.900 75.000 99.465 ;
        RECT 43.240 50.400 75.000 97.900 ;
        RECT 43.240 0.000 49.990 50.400 ;
        RECT 74.690 0.000 75.000 50.400 ;
      LAYER met4 ;
        RECT 4.800 97.700 70.200 173.100 ;
      LAYER met5 ;
        RECT 4.800 98.100 9.730 172.970 ;
        RECT 65.270 98.100 70.200 172.970 ;
  END
END sky130_fd_io__top_power_hvc_wpad

#--------EOF---------

MACRO sky130_fd_io__top_power_hvc_wpadv2
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_power_hvc_wpadv2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY X Y R90 ;
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.495 0.000 24.395 32.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 0.000 74.290 90.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.500 101.295 74.290 173.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.500 101.285 74.290 101.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.550 100.345 61.500 101.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.975 99.770 60.550 100.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.425 99.220 59.975 99.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.765 98.560 59.425 99.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.635 93.430 58.765 98.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.390 90.185 53.635 93.430 ;
    END
  END P_CORE
  PIN DRN_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 37.890 0.000 48.890 11.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 50.390 0.000 74.290 25.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 169.135 59.285 169.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 110.440 59.285 169.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.285 107.960 59.285 110.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.685 169.135 53.285 169.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.685 169.735 59.285 169.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 169.735 52.685 172.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.855 106.010 53.285 110.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 185.360 71.625 190.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.530 185.265 71.625 185.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.900 184.635 71.530 185.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.085 183.820 70.900 184.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 183.820 70.085 183.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.635 183.370 70.085 183.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 183.370 69.635 183.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.035 182.770 69.635 183.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 182.770 69.035 182.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.425 182.160 69.035 182.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.810 181.545 68.425 182.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.180 180.915 67.810 181.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.635 180.370 67.180 180.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 180.370 66.635 180.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.585 179.320 66.635 180.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 179.320 65.585 179.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.235 177.970 65.585 179.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 177.970 64.235 178.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.485 177.220 64.235 177.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 177.220 63.485 177.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.700 176.435 63.485 177.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.985 175.720 62.700 176.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 175.720 61.985 175.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.585 173.320 61.985 175.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 173.320 59.585 175.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.285 173.020 59.585 173.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.775 172.645 59.285 173.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.400 104.555 48.855 106.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 102.415 47.400 104.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.340 102.015 59.285 107.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 102.015 53.340 102.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.160 100.835 53.340 102.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.040 99.715 52.160 100.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.550 99.505 45.260 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 170.460 48.855 170.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 110.620 48.855 170.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.855 108.150 48.855 110.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.965 170.460 42.855 175.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 105.655 42.855 110.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.965 175.350 48.855 190.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.260 104.555 46.570 105.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.840 102.135 45.260 104.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 102.135 42.840 102.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 100.215 42.840 102.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 100.105 42.840 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.840 99.505 43.550 100.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 98.300 51.040 99.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.790 97.050 51.040 98.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 97.050 49.790 97.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.890 96.150 49.790 97.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.890 96.150 48.890 96.300 ;
    END
  END DRN_HVC
  PIN SRC_BDY_HVC
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 25.895 0.000 36.895 2.725 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.495 0.000 24.395 2.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.945 89.470 36.895 99.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.070 98.155 30.165 100.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 100.250 28.070 102.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 175.350 36.820 200.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.130 174.660 36.820 175.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.660 36.130 174.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.530 174.060 36.130 174.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 174.060 35.530 174.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.780 173.310 35.530 174.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 173.310 34.780 173.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.180 172.710 34.780 173.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 172.710 34.180 172.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.930 170.460 34.180 172.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 158.470 31.930 172.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 104.790 31.930 104.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.930 99.895 36.895 104.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 91.440 24.845 92.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.745 92.540 29.525 96.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.895 94.105 23.595 96.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.025 96.655 29.525 98.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 96.805 20.895 99.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.930 98.155 28.025 100.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 99.505 18.195 102.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 173.020 25.010 173.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 172.640 25.010 173.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.500 169.130 25.010 172.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 159.510 21.500 171.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.500 104.600 21.500 104.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.500 100.250 25.930 104.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.300 173.020 15.500 174.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.300 174.220 25.010 174.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.250 174.220 14.300 175.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.250 175.270 25.010 175.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.370 175.270 13.250 176.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.710 176.150 12.370 176.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 176.810 11.710 177.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.550 177.970 25.010 178.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.510 177.970 10.550 179.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.680 179.010 9.510 179.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 179.840 8.680 180.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.150 180.370 25.010 180.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 180.370 8.150 181.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.100 181.420 25.010 181.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.050 181.420 7.100 182.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.050 182.470 25.010 182.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.155 182.470 6.050 183.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 183.365 5.155 183.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.550 183.970 25.010 184.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 183.970 4.550 184.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.800 184.720 25.010 184.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.160 184.720 3.800 185.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.160 185.360 25.010 200.000 ;
    END
  END SRC_BDY_HVC
  PIN OGC_HVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 25.895 0.000 27.895 0.535 ;
    END
  END OGC_HVC
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN P_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 6.200 104.175 68.800 166.625 ;
    END
  END P_PAD
  OBS
      LAYER li1 ;
        RECT 0.610 0.970 72.855 199.695 ;
      LAYER met1 ;
        RECT 0.185 0.970 72.915 199.725 ;
      LAYER met2 ;
        RECT 0.265 25.940 74.290 195.075 ;
        RECT 0.265 2.335 50.110 25.940 ;
        RECT 24.675 0.980 50.110 2.335 ;
      LAYER met3 ;
        RECT 0.240 184.320 2.760 185.360 ;
        RECT 0.240 183.570 3.400 184.320 ;
        RECT 25.410 183.570 25.530 185.360 ;
        RECT 0.240 182.965 4.150 183.570 ;
        RECT 6.450 183.020 25.530 183.570 ;
        RECT 0.240 182.070 4.755 182.965 ;
        RECT 25.410 182.070 25.530 183.020 ;
        RECT 0.240 181.020 5.650 182.070 ;
        RECT 7.500 181.970 25.530 182.070 ;
        RECT 25.410 181.020 25.530 181.970 ;
        RECT 0.240 179.970 6.700 181.020 ;
        RECT 8.550 180.920 25.530 181.020 ;
        RECT 25.410 179.970 25.530 180.920 ;
        RECT 0.240 179.440 7.750 179.970 ;
        RECT 0.240 178.610 8.280 179.440 ;
        RECT 9.910 179.410 25.530 179.970 ;
        RECT 0.240 177.570 9.110 178.610 ;
        RECT 10.950 178.520 25.530 179.410 ;
        RECT 25.410 177.570 25.530 178.520 ;
        RECT 0.240 176.410 10.150 177.570 ;
        RECT 12.110 177.210 25.530 177.570 ;
        RECT 12.770 176.550 25.530 177.210 ;
        RECT 0.240 175.750 11.310 176.410 ;
        RECT 13.650 175.820 25.530 176.550 ;
        RECT 0.240 174.870 11.970 175.750 ;
        RECT 25.410 174.870 25.530 175.820 ;
        RECT 0.240 173.820 12.850 174.870 ;
        RECT 14.700 174.770 25.530 174.870 ;
        RECT 25.410 173.820 25.530 174.770 ;
        RECT 37.220 174.260 37.565 185.360 ;
        RECT 49.255 184.960 49.375 185.360 ;
        RECT 49.255 184.370 69.685 184.960 ;
        RECT 72.025 184.865 74.290 185.360 ;
        RECT 49.255 182.370 49.375 184.370 ;
        RECT 71.930 184.235 74.290 184.865 ;
        RECT 71.300 183.420 74.290 184.235 ;
        RECT 70.485 182.970 74.290 183.420 ;
        RECT 70.035 182.370 74.290 182.970 ;
        RECT 49.255 181.945 67.410 182.370 ;
        RECT 49.255 181.315 66.780 181.945 ;
        RECT 69.435 181.760 74.290 182.370 ;
        RECT 49.255 180.995 66.235 181.315 ;
        RECT 68.825 181.145 74.290 181.760 ;
        RECT 49.255 179.970 49.375 180.995 ;
        RECT 68.210 180.515 74.290 181.145 ;
        RECT 67.580 179.970 74.290 180.515 ;
        RECT 49.255 179.870 65.185 179.970 ;
        RECT 49.255 178.920 49.375 179.870 ;
        RECT 67.035 178.920 74.290 179.970 ;
        RECT 49.255 178.520 63.835 178.920 ;
        RECT 49.255 176.820 49.375 178.520 ;
        RECT 65.985 177.570 74.290 178.920 ;
        RECT 64.635 176.820 74.290 177.570 ;
        RECT 49.255 176.325 61.585 176.820 ;
        RECT 49.255 174.950 49.375 176.325 ;
        RECT 63.885 176.035 74.290 176.820 ;
        RECT 63.100 175.320 74.290 176.035 ;
        RECT 0.240 172.620 13.900 173.820 ;
        RECT 15.900 173.570 25.530 173.820 ;
        RECT 36.530 173.660 37.565 174.260 ;
        RECT 0.240 172.240 15.100 172.620 ;
        RECT 0.240 172.070 21.100 172.240 ;
        RECT 0.240 159.110 15.100 172.070 ;
        RECT 25.410 168.730 25.530 173.570 ;
        RECT 35.930 172.910 37.565 173.660 ;
        RECT 35.180 172.310 37.565 172.910 ;
        RECT 34.580 170.060 37.565 172.310 ;
        RECT 43.255 171.010 49.375 174.950 ;
        RECT 62.385 173.720 74.290 175.320 ;
        RECT 59.985 172.620 61.100 172.920 ;
        RECT 59.685 172.245 61.100 172.620 ;
        RECT 21.900 159.110 25.530 168.730 ;
        RECT 0.240 158.070 25.530 159.110 ;
        RECT 32.330 158.070 42.455 170.060 ;
        RECT 0.240 111.020 42.455 158.070 ;
        RECT 49.255 169.335 49.375 171.010 ;
        RECT 53.085 170.285 61.100 172.245 ;
        RECT 49.255 168.735 52.285 169.335 ;
        RECT 0.240 105.260 37.490 111.020 ;
        RECT 49.255 110.840 52.885 168.735 ;
        RECT 0.240 105.080 25.530 105.260 ;
        RECT 37.295 105.255 37.490 105.260 ;
        RECT 43.255 106.410 48.455 107.750 ;
        RECT 43.255 106.265 47.000 106.410 ;
        RECT 43.255 105.255 44.860 106.265 ;
        RECT 0.240 104.200 15.100 105.080 ;
        RECT 37.295 104.955 44.860 105.255 ;
        RECT 46.970 104.955 47.000 106.265 ;
        RECT 0.240 102.600 21.100 104.200 ;
        RECT 26.330 102.790 31.530 104.390 ;
        RECT 0.240 99.105 15.100 102.600 ;
        RECT 18.595 99.905 21.100 102.600 ;
        RECT 28.470 100.650 31.530 102.790 ;
        RECT 0.240 96.405 17.795 99.105 ;
        RECT 21.295 97.755 25.530 99.850 ;
        RECT 30.565 99.495 31.530 100.650 ;
        RECT 37.295 102.685 42.440 104.955 ;
        RECT 49.255 104.155 52.940 105.610 ;
        RECT 30.565 97.755 31.545 99.495 ;
        RECT 21.295 97.205 27.625 97.755 ;
        RECT 23.995 97.055 27.625 97.205 ;
        RECT 0.240 93.705 20.495 96.405 ;
        RECT 0.240 91.040 23.345 93.705 ;
        RECT 29.925 92.140 31.545 97.755 ;
        RECT 25.245 91.040 31.545 92.140 ;
        RECT 0.240 89.070 31.545 91.040 ;
        RECT 37.295 97.900 37.490 102.685 ;
        RECT 47.800 102.565 52.940 104.155 ;
        RECT 43.240 101.615 44.860 101.735 ;
        RECT 59.685 101.695 61.100 170.285 ;
        RECT 59.685 101.615 60.150 101.695 ;
        RECT 43.240 101.235 51.760 101.615 ;
        RECT 43.240 100.615 50.640 101.235 ;
        RECT 43.950 99.905 44.150 100.615 ;
        RECT 45.660 99.905 50.640 100.615 ;
        RECT 53.740 100.745 60.150 101.615 ;
        RECT 53.740 100.435 59.575 100.745 ;
        RECT 52.560 100.170 59.575 100.435 ;
        RECT 52.560 99.620 59.025 100.170 ;
        RECT 61.900 99.945 74.290 100.885 ;
        RECT 52.560 99.315 58.365 99.620 ;
        RECT 60.950 99.370 74.290 99.945 ;
        RECT 51.440 98.960 58.365 99.315 ;
        RECT 37.295 97.600 49.390 97.900 ;
        RECT 37.295 95.750 37.490 97.600 ;
        RECT 51.440 96.650 53.235 98.960 ;
        RECT 60.375 98.820 74.290 99.370 ;
        RECT 59.825 98.160 74.290 98.820 ;
        RECT 50.190 95.750 53.235 96.650 ;
        RECT 37.295 93.830 53.235 95.750 ;
        RECT 37.295 89.070 49.990 93.830 ;
        RECT 59.165 93.030 74.290 98.160 ;
        RECT 54.035 90.585 74.290 93.030 ;
        RECT 0.240 32.915 49.990 89.070 ;
        RECT 24.795 11.730 49.990 32.915 ;
        RECT 24.795 3.125 37.490 11.730 ;
        RECT 24.795 2.725 25.495 3.125 ;
        RECT 37.295 2.725 37.490 3.125 ;
        RECT 49.290 2.725 49.990 11.730 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 168.225 75.000 174.185 ;
        RECT 0.000 102.575 4.600 168.225 ;
        RECT 70.400 102.575 75.000 168.225 ;
        RECT 0.000 96.585 75.000 102.575 ;
        RECT 2.870 36.840 72.130 96.585 ;
        RECT 0.000 36.835 75.000 36.840 ;
        RECT 2.870 18.285 72.130 36.835 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__top_power_hvc_wpadv2

#--------EOF---------

MACRO sky130_fd_io__top_power_lvc_wpad
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_power_lvc_wpad ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 198.000 ;
  SYMMETRY X Y R90 ;
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 23.835 1.270 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 23.835 75.000 28.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 173.785 75.000 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 173.785 1.270 198.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 23.935 75.000 28.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 23.935 1.270 28.385 ;
    END
  END VSSIO
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 49.645 75.000 50.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 45.735 75.000 46.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 54.405 75.000 54.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 34.735 1.270 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 34.735 75.000 38.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 49.645 1.270 50.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 34.840 75.000 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 45.735 75.000 54.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 34.840 1.270 38.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 45.735 1.270 54.735 ;
    END
  END VSSA
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 56.235 1.270 60.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 56.235 75.000 60.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 56.335 1.270 60.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 56.335 75.000 60.585 ;
    END
  END VSSIO_Q
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 0.035 1.270 5.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 0.035 75.000 5.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 0.135 75.000 5.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 0.135 1.270 5.385 ;
    END
  END VCCHIB
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 6.885 1.270 11.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 6.885 75.000 11.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 6.985 75.000 11.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 6.985 1.270 11.435 ;
    END
  END VCCD
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 12.935 0.965 16.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.035 12.935 75.000 16.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 13.035 75.000 16.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 13.035 0.965 16.285 ;
    END
  END VDDA
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 17.785 1.270 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 17.785 75.000 22.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 68.035 1.270 93.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 68.035 75.000 93.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 68.035 75.000 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 17.885 75.000 22.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 68.035 1.270 92.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 17.885 1.270 22.335 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 29.885 1.270 33.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 29.885 75.000 33.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 29.985 75.000 33.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 29.985 1.270 33.235 ;
    END
  END VSWITCH
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 0.000 62.085 1.270 66.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 62.085 75.000 66.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 62.185 75.000 66.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 62.185 1.270 66.435 ;
    END
  END VDDIO_Q
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 51.125 75.000 54.105 ;
    END
  END AMUXBUS_A
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 46.365 75.000 49.345 ;
    END
  END AMUXBUS_B
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 39.585 1.270 44.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 39.585 75.000 44.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 39.685 75.000 44.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 39.685 1.270 44.135 ;
    END
  END VSSD
  PIN P_PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 9.315 100.140 65.955 167.570 ;
    END
  END P_PAD
  PIN SRC_BDY_LVC1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 0.500 0.000 20.495 1.485 ;
    END
  END SRC_BDY_LVC1
  PIN SRC_BDY_LVC2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.715 0.000 74.700 3.660 ;
    END
  END SRC_BDY_LVC2
  PIN BDY2_B2B
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 34.440 0.000 44.440 0.325 ;
    END
  END BDY2_B2B
  PIN DRN_LVC2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 38.380 0.000 49.255 22.900 ;
    END
  END DRN_LVC2
  PIN DRN_LVC1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 26.000 0.000 36.880 20.220 ;
    END
  END DRN_LVC1
  PIN P_CORE
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 50.755 0.000 74.700 84.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.500 0.000 24.500 70.755 ;
    END
  END P_CORE
  PIN OGC_LVC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 26.210 0.000 27.700 0.170 ;
    END
  END OGC_LVC
  OBS
      LAYER li1 ;
        RECT 0.240 1.020 74.755 197.780 ;
      LAYER met1 ;
        RECT 0.120 0.450 74.785 197.840 ;
        RECT 0.120 0.000 25.930 0.450 ;
        RECT 27.980 0.000 74.785 0.450 ;
      LAYER met2 ;
        RECT 0.500 3.940 74.700 194.430 ;
        RECT 0.500 1.765 54.435 3.940 ;
        RECT 20.775 0.605 54.435 1.765 ;
        RECT 20.775 0.000 34.160 0.605 ;
        RECT 44.720 0.000 54.435 0.605 ;
      LAYER met3 ;
        RECT 0.500 84.865 74.700 189.515 ;
        RECT 0.500 71.155 50.355 84.865 ;
        RECT 24.900 23.300 50.355 71.155 ;
        RECT 24.900 20.620 37.980 23.300 ;
        RECT 24.900 17.790 25.600 20.620 ;
        RECT 37.280 17.790 37.980 20.620 ;
        RECT 49.655 17.790 50.355 23.300 ;
      LAYER met4 ;
        RECT 1.670 173.385 73.330 198.000 ;
        RECT 0.965 93.400 74.035 173.385 ;
        RECT 1.670 67.635 73.330 93.400 ;
        RECT 0.965 66.935 74.035 67.635 ;
        RECT 1.670 61.685 73.330 66.935 ;
        RECT 0.965 61.085 74.035 61.685 ;
        RECT 1.670 55.835 73.330 61.085 ;
        RECT 0.965 55.135 74.035 55.835 ;
        RECT 1.670 49.745 73.330 50.725 ;
        RECT 0.965 44.635 74.035 45.335 ;
        RECT 1.670 39.185 73.330 44.635 ;
        RECT 0.965 38.585 74.035 39.185 ;
        RECT 1.670 34.335 73.330 38.585 ;
        RECT 0.965 33.735 74.035 34.335 ;
        RECT 1.670 29.485 73.330 33.735 ;
        RECT 0.965 28.885 74.035 29.485 ;
        RECT 1.670 23.435 73.330 28.885 ;
        RECT 0.965 22.835 74.035 23.435 ;
        RECT 1.670 17.385 73.330 22.835 ;
        RECT 0.965 16.785 74.035 17.385 ;
        RECT 1.365 12.535 73.635 16.785 ;
        RECT 0.965 11.935 74.035 12.535 ;
        RECT 1.670 6.485 73.330 11.935 ;
        RECT 0.965 5.885 74.035 6.485 ;
        RECT 1.670 0.035 73.330 5.885 ;
      LAYER met5 ;
        RECT 2.870 172.185 72.130 198.000 ;
        RECT 0.000 169.170 75.000 172.185 ;
        RECT 0.000 98.540 7.715 169.170 ;
        RECT 67.555 98.540 75.000 169.170 ;
        RECT 0.000 94.585 75.000 98.540 ;
        RECT 2.870 34.840 72.130 94.585 ;
        RECT 0.000 34.835 75.000 34.840 ;
        RECT 2.870 16.285 72.130 34.835 ;
        RECT 2.565 13.035 72.435 16.285 ;
        RECT 2.870 0.135 72.130 13.035 ;
  END
END sky130_fd_io__top_power_lvc_wpad

#--------EOF---------

MACRO sky130_fd_io__top_xres4v2
  CLASS PAD ;
  FOREIGN sky130_fd_io__top_xres4v2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 200.000 ;
  SYMMETRY R90 ;
  PIN PAD_A_ESD_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.245 0.000 18.910 0.565 ;
    END
    PORT
      LAYER met2 ;
        RECT 17.245 0.000 18.910 0.565 ;
    END
  END PAD_A_ESD_H
  PIN XRES_H_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.935 0.000 29.665 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 28.935 0.000 29.665 0.330 ;
    END
  END XRES_H_N
  PIN FILT_IN_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.075 0.000 21.225 1.410 ;
    END
    PORT
      LAYER met2 ;
        RECT 20.075 0.000 21.225 1.410 ;
    END
  END FILT_IN_H
  PIN ENABLE_VDDIO
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.400 0.000 8.920 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 8.425 0.000 8.895 0.330 ;
    END
  END ENABLE_VDDIO
  PIN TIE_WEAK_HI_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.190 0.000 73.260 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 72.215 0.000 73.235 0.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.190 49.985 73.925 64.465 ;
    END
  END TIE_WEAK_HI_H
  PIN ENABLE_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.285 0.000 12.545 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 12.285 0.000 12.545 0.330 ;
    END
  END ENABLE_H
  PIN PULLUP_H
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.555 0.000 15.135 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 14.555 0.000 15.135 0.330 ;
    END
  END PULLUP_H
  PIN EN_VDDIO_SIG_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.360 0.000 22.660 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 22.360 0.000 22.660 0.330 ;
    END
    PORT
      LAYER met2 ;
        RECT 29.320 5.360 29.580 11.085 ;
    END
  END EN_VDDIO_SIG_H
  PIN TIE_LO_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.580 0.000 28.230 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 27.580 0.000 28.230 0.330 ;
    END
  END TIE_LO_ESD
  PIN TIE_HI_ESD
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.505 0.000 31.155 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 30.505 0.000 31.155 0.330 ;
    END
  END TIE_HI_ESD
  PIN DISABLE_PULLUP_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.760 0.000 33.020 0.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 32.760 0.000 33.020 0.330 ;
    END
  END DISABLE_PULLUP_H
  PIN INP_SEL_H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 24.905 0.000 25.135 9.975 ;
    END
  END INP_SEL_H
  PIN VSSIO
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 25.835 75.000 30.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 25.835 1.270 30.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 175.785 1.270 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 25.935 75.000 30.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 175.785 75.000 200.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 25.935 1.270 30.385 ;
    END
  END VSSIO
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 36.735 75.000 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 56.405 75.000 56.735 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 47.735 75.000 48.065 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 51.645 75.000 52.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 36.735 1.270 40.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 51.645 1.270 52.825 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 47.735 75.000 56.735 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 36.840 75.000 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 36.840 1.270 40.085 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 47.735 1.270 56.735 ;
    END
  END VSSA
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 41.585 75.000 46.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 41.585 1.270 46.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 41.685 75.000 46.135 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 41.685 1.270 46.135 ;
    END
  END VSSD
  PIN AMUXBUS_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 48.365 75.000 51.345 ;
    END
  END AMUXBUS_B
  PIN AMUXBUS_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.000 53.125 75.000 56.105 ;
    END
  END AMUXBUS_A
  PIN VDDIO_Q
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 64.085 75.000 68.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 64.085 1.270 68.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 64.185 75.000 68.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 64.185 1.270 68.435 ;
    END
  END VDDIO_Q
  PIN VDDIO
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 70.035 75.000 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.730 19.785 75.000 24.435 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 70.035 1.270 95.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 19.785 1.270 24.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 19.885 75.000 24.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 70.035 75.000 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 70.035 1.270 94.985 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 19.885 1.270 24.335 ;
    END
  END VDDIO
  PIN VSWITCH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 31.885 75.000 35.335 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 31.885 1.270 35.335 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 31.985 75.000 35.235 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 31.985 1.270 35.235 ;
    END
  END VSWITCH
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 74.035 14.935 75.000 18.385 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 14.935 0.965 18.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 74.035 15.035 75.000 18.285 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 15.035 0.965 18.285 ;
    END
  END VDDA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 8.885 75.000 13.535 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 8.885 1.270 13.535 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 8.985 75.000 13.435 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 8.985 1.270 13.435 ;
    END
  END VCCD
  PIN VCCHIB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 73.730 2.035 75.000 7.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 2.035 1.270 7.485 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 2.135 75.000 7.385 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 2.135 1.270 7.385 ;
    END
  END VCCHIB
  PIN VSSIO_Q
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 73.730 58.235 75.000 62.685 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.000 58.235 1.270 62.685 ;
    END
    PORT
      LAYER met5 ;
        RECT 73.730 58.335 75.000 62.585 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.000 58.335 1.270 62.585 ;
    END
  END VSSIO_Q
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 17.250 108.455 54.435 164.285 ;
    END
  END PAD
  OBS
      LAYER nwell ;
        RECT -0.515 168.515 75.620 170.210 ;
        RECT -0.515 146.690 1.675 168.515 ;
        RECT 73.095 146.690 75.620 168.515 ;
        RECT -0.515 144.880 75.620 146.690 ;
      LAYER pwell ;
        RECT -0.290 140.685 75.290 144.565 ;
      LAYER nwell ;
        RECT -0.330 130.665 75.330 140.380 ;
      LAYER pwell ;
        RECT -0.130 129.315 41.750 130.355 ;
        RECT 61.910 129.315 75.130 130.355 ;
        RECT -0.130 124.135 75.130 129.315 ;
        RECT -0.130 102.525 1.435 124.135 ;
        RECT 73.560 102.525 75.130 124.135 ;
        RECT -0.130 99.230 75.130 102.525 ;
        RECT -0.130 97.995 58.470 99.230 ;
        RECT 71.930 97.995 75.130 99.230 ;
        RECT -0.130 96.735 75.130 97.995 ;
        RECT -0.130 96.730 58.470 96.735 ;
      LAYER li1 ;
        RECT 0.000 144.435 75.000 199.220 ;
        RECT -0.160 140.815 75.160 144.435 ;
        RECT 0.000 130.225 75.000 140.815 ;
        RECT -0.265 101.395 75.000 130.225 ;
        RECT 0.000 0.185 75.000 101.395 ;
      LAYER met1 ;
        RECT 0.000 170.090 75.000 199.210 ;
        RECT -0.145 131.275 75.145 170.090 ;
        RECT 0.000 130.220 75.000 131.275 ;
        RECT -0.145 95.895 75.145 130.220 ;
        RECT 0.000 10.255 75.000 95.895 ;
        RECT 0.000 0.610 24.625 10.255 ;
        RECT 0.000 0.185 12.005 0.610 ;
        RECT 12.825 0.185 14.275 0.610 ;
        RECT 15.415 0.185 22.080 0.610 ;
        RECT 22.940 0.185 24.625 0.610 ;
        RECT 25.415 0.610 75.000 10.255 ;
        RECT 25.415 0.185 27.300 0.610 ;
        RECT 28.510 0.185 30.225 0.610 ;
        RECT 31.435 0.185 32.480 0.610 ;
        RECT 33.300 0.185 75.000 0.610 ;
      LAYER met2 ;
        RECT 0.340 11.365 74.915 199.210 ;
        RECT 0.340 5.080 29.040 11.365 ;
        RECT 29.860 5.080 74.915 11.365 ;
        RECT 0.340 1.690 74.915 5.080 ;
        RECT 0.340 0.845 19.795 1.690 ;
        RECT 0.340 0.610 16.965 0.845 ;
        RECT 0.340 0.000 8.145 0.610 ;
        RECT 9.175 0.000 12.005 0.610 ;
        RECT 12.825 0.000 14.275 0.610 ;
        RECT 15.415 0.000 16.965 0.610 ;
        RECT 19.190 0.000 19.795 0.845 ;
        RECT 21.505 0.610 74.915 1.690 ;
        RECT 21.505 0.000 22.080 0.610 ;
        RECT 22.940 0.000 27.300 0.610 ;
        RECT 28.510 0.000 28.655 0.610 ;
        RECT 29.945 0.000 30.225 0.610 ;
        RECT 31.435 0.000 32.480 0.610 ;
        RECT 33.300 0.000 71.935 0.610 ;
        RECT 73.515 0.000 74.915 0.610 ;
      LAYER met3 ;
        RECT 0.965 64.865 74.700 200.000 ;
        RECT 0.965 49.585 71.790 64.865 ;
        RECT 74.325 49.585 74.700 64.865 ;
        RECT 0.965 1.810 74.700 49.585 ;
        RECT 0.965 0.965 19.675 1.810 ;
        RECT 0.965 0.730 16.845 0.965 ;
        RECT 0.965 0.330 8.000 0.730 ;
        RECT 9.320 0.330 16.845 0.730 ;
        RECT 19.310 0.330 19.675 0.965 ;
        RECT 21.625 0.730 74.700 1.810 ;
        RECT 21.625 0.330 28.535 0.730 ;
        RECT 30.065 0.330 71.790 0.730 ;
        RECT 73.660 0.330 74.700 0.730 ;
      LAYER met4 ;
        RECT 1.670 175.385 73.330 200.000 ;
        RECT 0.965 95.400 74.035 175.385 ;
        RECT 1.670 69.635 73.330 95.400 ;
        RECT 0.965 68.935 74.035 69.635 ;
        RECT 1.670 63.685 73.330 68.935 ;
        RECT 0.965 63.085 74.035 63.685 ;
        RECT 1.670 57.835 73.330 63.085 ;
        RECT 0.965 57.135 74.035 57.835 ;
        RECT 1.670 51.745 73.330 52.725 ;
        RECT 0.965 46.635 74.035 47.335 ;
        RECT 1.670 41.185 73.330 46.635 ;
        RECT 0.965 40.585 74.035 41.185 ;
        RECT 1.670 36.335 73.330 40.585 ;
        RECT 0.965 35.735 74.035 36.335 ;
        RECT 1.670 31.485 73.330 35.735 ;
        RECT 0.965 30.885 74.035 31.485 ;
        RECT 1.670 25.435 73.330 30.885 ;
        RECT 0.965 24.835 74.035 25.435 ;
        RECT 1.670 19.385 73.330 24.835 ;
        RECT 0.965 18.785 74.035 19.385 ;
        RECT 1.365 14.535 73.635 18.785 ;
        RECT 0.965 13.935 74.035 14.535 ;
        RECT 1.670 8.485 73.330 13.935 ;
        RECT 0.965 7.885 74.035 8.485 ;
        RECT 1.670 2.035 73.330 7.885 ;
      LAYER met5 ;
        RECT 2.870 174.185 72.130 200.000 ;
        RECT 0.000 165.885 75.000 174.185 ;
        RECT 0.000 106.855 15.650 165.885 ;
        RECT 56.035 106.855 75.000 165.885 ;
        RECT 0.000 96.585 75.000 106.855 ;
        RECT 2.870 18.285 72.130 96.585 ;
        RECT 2.565 15.035 72.435 18.285 ;
        RECT 2.870 2.135 72.130 15.035 ;
  END
END sky130_fd_io__top_xres4v2

#--------EOF---------


END LIBRARY
