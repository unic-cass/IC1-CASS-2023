magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 130 827
rect 384 261 596 827
rect 850 261 1326 827
<< pwell >>
rect 511 1050 1111 1067
rect 3 893 89 1050
rect 511 893 1285 1050
rect 511 885 1111 893
rect 3 38 89 195
rect 601 192 1253 203
rect 398 56 1253 192
rect 601 21 1253 56
<< scnmos >>
rect 590 911 620 1041
rect 676 911 706 1041
rect 762 911 792 1041
rect 848 911 878 1041
rect 1002 911 1032 1041
rect 477 82 507 166
rect 684 47 714 177
rect 770 47 800 177
rect 856 47 886 177
rect 942 47 972 177
rect 1036 47 1066 177
rect 1140 47 1170 177
<< scpmoshvt >>
rect 941 618 971 776
rect 1032 618 1062 776
rect 475 297 505 497
rect 941 312 971 470
rect 1036 297 1066 497
rect 1140 297 1170 497
<< ndiff >>
rect 537 1025 590 1041
rect 537 991 545 1025
rect 579 991 590 1025
rect 537 957 590 991
rect 537 923 545 957
rect 579 923 590 957
rect 537 911 590 923
rect 620 1032 676 1041
rect 620 998 631 1032
rect 665 998 676 1032
rect 620 964 676 998
rect 620 930 631 964
rect 665 930 676 964
rect 620 911 676 930
rect 706 1032 762 1041
rect 706 998 717 1032
rect 751 998 762 1032
rect 706 964 762 998
rect 706 930 717 964
rect 751 930 762 964
rect 706 911 762 930
rect 792 1032 848 1041
rect 792 998 803 1032
rect 837 998 848 1032
rect 792 964 848 998
rect 792 930 803 964
rect 837 930 848 964
rect 792 911 848 930
rect 878 1032 1002 1041
rect 878 930 889 1032
rect 991 930 1002 1032
rect 878 911 1002 930
rect 1032 1025 1085 1041
rect 1032 991 1043 1025
rect 1077 991 1085 1025
rect 1032 957 1085 991
rect 1032 923 1043 957
rect 1077 923 1085 957
rect 1032 911 1085 923
rect 627 169 684 177
rect 424 141 477 166
rect 424 107 432 141
rect 466 107 477 141
rect 424 82 477 107
rect 507 141 560 166
rect 507 107 518 141
rect 552 107 560 141
rect 507 82 560 107
rect 627 135 639 169
rect 673 135 684 169
rect 627 101 684 135
rect 627 67 639 101
rect 673 67 684 101
rect 627 47 684 67
rect 714 169 770 177
rect 714 135 725 169
rect 759 135 770 169
rect 714 101 770 135
rect 714 67 725 101
rect 759 67 770 101
rect 714 47 770 67
rect 800 101 856 177
rect 800 67 811 101
rect 845 67 856 101
rect 800 47 856 67
rect 886 169 942 177
rect 886 135 897 169
rect 931 135 942 169
rect 886 101 942 135
rect 886 67 897 101
rect 931 67 942 101
rect 886 47 942 67
rect 972 169 1036 177
rect 972 135 983 169
rect 1017 135 1036 169
rect 972 101 1036 135
rect 972 67 983 101
rect 1017 67 1036 101
rect 972 47 1036 67
rect 1066 169 1140 177
rect 1066 135 1077 169
rect 1111 135 1140 169
rect 1066 101 1140 135
rect 1066 67 1077 101
rect 1111 67 1140 101
rect 1066 47 1140 67
rect 1170 169 1227 177
rect 1170 135 1181 169
rect 1215 135 1227 169
rect 1170 101 1227 135
rect 1170 67 1181 101
rect 1215 67 1227 101
rect 1170 47 1227 67
<< pdiff >>
rect 886 732 941 776
rect 886 698 896 732
rect 930 698 941 732
rect 886 664 941 698
rect 886 630 894 664
rect 928 630 941 664
rect 886 618 941 630
rect 971 732 1032 776
rect 971 698 984 732
rect 1018 698 1032 732
rect 971 664 1032 698
rect 971 630 984 664
rect 1018 630 1032 664
rect 971 618 1032 630
rect 1062 732 1116 776
rect 1062 698 1074 732
rect 1108 698 1116 732
rect 1062 664 1116 698
rect 1062 630 1074 664
rect 1108 630 1116 664
rect 1062 618 1116 630
rect 420 458 475 497
rect 420 424 428 458
rect 462 424 475 458
rect 420 375 475 424
rect 420 341 428 375
rect 462 341 475 375
rect 420 297 475 341
rect 505 458 560 497
rect 505 424 518 458
rect 552 424 560 458
rect 505 375 560 424
rect 986 470 1036 497
rect 886 458 941 470
rect 886 424 894 458
rect 928 424 941 458
rect 505 341 518 375
rect 552 341 560 375
rect 505 297 560 341
rect 886 375 941 424
rect 886 341 894 375
rect 928 341 941 375
rect 886 312 941 341
rect 971 458 1036 470
rect 971 424 984 458
rect 1018 424 1036 458
rect 971 375 1036 424
rect 971 341 984 375
rect 1018 341 1036 375
rect 971 312 1036 341
rect 986 297 1036 312
rect 1066 458 1140 497
rect 1066 424 1077 458
rect 1111 424 1140 458
rect 1066 375 1140 424
rect 1066 341 1077 375
rect 1111 341 1140 375
rect 1066 297 1140 341
rect 1170 458 1227 497
rect 1170 424 1181 458
rect 1215 424 1227 458
rect 1170 375 1227 424
rect 1170 341 1181 375
rect 1215 341 1227 375
rect 1170 297 1227 341
<< ndiffc >>
rect 545 991 579 1025
rect 545 923 579 957
rect 631 998 665 1032
rect 631 930 665 964
rect 717 998 751 1032
rect 717 930 751 964
rect 803 998 837 1032
rect 803 930 837 964
rect 889 930 991 1032
rect 1043 991 1077 1025
rect 1043 923 1077 957
rect 432 107 466 141
rect 518 107 552 141
rect 639 135 673 169
rect 639 67 673 101
rect 725 135 759 169
rect 725 67 759 101
rect 811 67 845 101
rect 897 135 931 169
rect 897 67 931 101
rect 983 135 1017 169
rect 983 67 1017 101
rect 1077 135 1111 169
rect 1077 67 1111 101
rect 1181 135 1215 169
rect 1181 67 1215 101
<< pdiffc >>
rect 896 698 930 732
rect 894 630 928 664
rect 984 698 1018 732
rect 984 630 1018 664
rect 1074 698 1108 732
rect 1074 630 1108 664
rect 428 424 462 458
rect 428 341 462 375
rect 518 424 552 458
rect 894 424 928 458
rect 518 341 552 375
rect 894 341 928 375
rect 984 424 1018 458
rect 984 341 1018 375
rect 1077 424 1111 458
rect 1077 341 1111 375
rect 1181 424 1215 458
rect 1181 341 1215 375
<< psubdiff >>
rect 29 977 63 1024
rect 29 919 63 943
rect 1225 977 1259 1024
rect 1225 919 1259 943
rect 29 145 63 169
rect 29 64 63 111
<< nsubdiff >>
rect 29 759 63 783
rect 29 675 63 725
rect 420 715 560 743
rect 420 681 434 715
rect 468 681 512 715
rect 546 681 560 715
rect 420 654 560 681
rect 29 608 63 641
rect 1225 759 1259 783
rect 1225 675 1259 725
rect 1225 608 1259 641
<< psubdiffcont >>
rect 29 943 63 977
rect 1225 943 1259 977
rect 29 111 63 145
<< nsubdiffcont >>
rect 29 725 63 759
rect 29 641 63 675
rect 434 681 468 715
rect 512 681 546 715
rect 1225 725 1259 759
rect 1225 641 1259 675
<< poly >>
rect 590 1041 620 1067
rect 676 1041 706 1067
rect 762 1041 792 1067
rect 848 1041 878 1067
rect 1002 1041 1032 1067
rect 590 896 620 911
rect 676 896 706 911
rect 762 896 792 911
rect 848 896 878 911
rect 590 866 878 896
rect 612 785 682 866
rect 1002 824 1032 911
rect 1142 871 1211 875
rect 1140 859 1211 871
rect 1140 825 1167 859
rect 1201 825 1211 859
rect 612 751 628 785
rect 662 751 682 785
rect 612 735 682 751
rect 788 812 1062 824
rect 788 778 804 812
rect 838 794 1062 812
rect 838 778 854 794
rect 788 644 854 778
rect 941 776 971 794
rect 1032 776 1062 794
rect 1140 803 1211 825
rect 788 610 804 644
rect 838 610 854 644
rect 788 603 854 610
rect 941 603 971 618
rect 1032 603 1062 618
rect 788 573 1062 603
rect 475 497 505 523
rect 788 501 971 531
rect 788 499 854 501
rect 788 465 804 499
rect 838 465 854 499
rect 941 470 971 501
rect 1036 497 1066 531
rect 1140 497 1170 803
rect 788 431 854 465
rect 788 397 804 431
rect 838 397 854 431
rect 788 381 854 397
rect 475 245 505 297
rect 941 286 971 312
rect 1036 282 1066 297
rect 1140 282 1170 297
rect 592 267 658 280
rect 592 245 608 267
rect 475 233 608 245
rect 642 245 658 267
rect 642 244 726 245
rect 642 233 972 244
rect 475 214 972 233
rect 475 202 507 214
rect 477 166 507 202
rect 684 177 714 214
rect 770 177 800 214
rect 856 177 886 214
rect 942 177 972 214
rect 1036 217 1170 282
rect 1036 177 1066 217
rect 1140 177 1170 217
rect 477 21 507 82
rect 684 21 714 47
rect 770 21 800 47
rect 856 21 886 47
rect 942 21 972 47
rect 1036 21 1066 47
rect 1140 21 1170 47
<< polycont >>
rect 1167 825 1201 859
rect 628 751 662 785
rect 804 778 838 812
rect 804 610 838 644
rect 804 465 838 499
rect 804 397 838 431
rect 608 233 642 267
<< locali >>
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1288 1105
rect 17 977 75 1071
rect 17 943 29 977
rect 63 943 75 977
rect 17 926 75 943
rect 529 1025 581 1071
rect 529 991 545 1025
rect 579 991 581 1025
rect 529 957 581 991
rect 529 923 545 957
rect 579 923 581 957
rect 529 903 581 923
rect 615 1032 681 1037
rect 615 998 631 1032
rect 665 998 681 1032
rect 615 964 681 998
rect 615 930 631 964
rect 665 930 681 964
rect 615 865 681 930
rect 715 1032 753 1071
rect 715 998 717 1032
rect 751 998 753 1032
rect 715 964 753 998
rect 715 930 717 964
rect 751 930 753 964
rect 715 903 753 930
rect 787 1032 853 1037
rect 787 998 803 1032
rect 837 998 853 1032
rect 787 964 853 998
rect 787 930 803 964
rect 837 930 853 964
rect 787 865 853 930
rect 889 1032 991 1071
rect 889 903 991 930
rect 1027 1025 1097 1032
rect 1027 991 1043 1025
rect 1077 991 1097 1025
rect 1027 964 1097 991
rect 1213 977 1271 1071
rect 1027 957 1139 964
rect 1027 923 1043 957
rect 1077 923 1139 957
rect 1213 943 1225 977
rect 1259 943 1271 977
rect 1213 926 1271 943
rect 1027 892 1139 923
rect 1027 881 1153 892
rect 615 853 853 865
rect 1072 871 1153 881
rect 1072 859 1217 871
rect 629 831 839 853
rect 804 812 838 831
rect 17 759 75 794
rect 17 731 29 759
rect 17 697 28 731
rect 63 725 75 759
rect 612 785 678 793
rect 612 751 628 785
rect 662 751 678 785
rect 804 762 838 778
rect 1072 825 1167 859
rect 1201 825 1217 859
rect 62 697 75 725
rect 17 675 75 697
rect 17 641 29 675
rect 63 641 75 675
rect 17 597 75 641
rect 412 715 562 750
rect 412 681 434 715
rect 468 681 512 715
rect 546 681 562 715
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 378 561
rect 412 532 562 681
rect 412 467 478 532
rect 612 474 678 751
rect 882 732 944 748
rect 882 728 896 732
rect 736 698 896 728
rect 930 698 944 732
rect 736 694 944 698
rect 736 515 770 694
rect 878 664 944 694
rect 804 644 838 660
rect 878 630 894 664
rect 928 630 944 664
rect 878 617 944 630
rect 978 732 1024 748
rect 978 698 984 732
rect 1018 698 1024 732
rect 978 664 1024 698
rect 978 630 984 664
rect 1018 630 1024 664
rect 804 583 838 610
rect 804 549 928 583
rect 736 499 838 515
rect 736 481 804 499
rect 276 458 478 467
rect 276 457 428 458
rect 276 423 284 457
rect 318 423 356 457
rect 390 423 428 457
rect 462 423 478 458
rect 276 413 478 423
rect 412 375 478 413
rect 412 341 428 375
rect 462 341 478 375
rect 412 327 478 341
rect 512 458 678 474
rect 512 424 518 458
rect 552 426 678 458
rect 804 431 838 465
rect 552 424 560 426
rect 512 375 560 424
rect 512 341 518 375
rect 552 341 560 375
rect 17 145 75 162
rect 17 111 29 145
rect 63 111 75 145
rect 17 17 75 111
rect 404 141 470 179
rect 404 107 432 141
rect 466 107 470 141
rect 404 17 470 107
rect 512 141 560 341
rect 594 267 658 308
rect 594 233 608 267
rect 642 233 658 267
rect 594 214 658 233
rect 804 196 838 397
rect 894 458 928 549
rect 894 375 928 424
rect 894 325 928 341
rect 978 561 1024 630
rect 1072 732 1110 825
rect 1072 698 1074 732
rect 1108 698 1110 732
rect 1072 664 1110 698
rect 1072 630 1074 664
rect 1108 630 1110 664
rect 1072 614 1110 630
rect 1213 759 1271 791
rect 1213 731 1225 759
rect 1213 697 1214 731
rect 1259 725 1271 759
rect 1248 697 1271 725
rect 1213 675 1271 697
rect 1213 641 1225 675
rect 1259 641 1271 675
rect 1213 597 1271 641
rect 978 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 978 458 1024 527
rect 978 424 984 458
rect 1018 424 1024 458
rect 978 375 1024 424
rect 978 341 984 375
rect 1018 341 1024 375
rect 978 325 1024 341
rect 1072 458 1127 474
rect 1072 424 1077 458
rect 1111 424 1127 458
rect 1072 375 1127 424
rect 1072 341 1077 375
rect 1111 341 1127 375
rect 1072 196 1127 341
rect 1181 458 1215 527
rect 1181 375 1215 424
rect 1181 322 1215 341
rect 512 107 518 141
rect 552 107 560 141
rect 512 75 560 107
rect 623 169 689 180
rect 623 135 639 169
rect 673 135 689 169
rect 623 101 689 135
rect 623 67 639 101
rect 673 67 689 101
rect 623 17 689 67
rect 723 169 933 196
rect 723 135 725 169
rect 759 146 897 169
rect 759 135 761 146
rect 723 101 761 135
rect 895 135 897 146
rect 931 135 933 169
rect 723 67 725 101
rect 759 67 761 101
rect 723 51 761 67
rect 795 101 861 112
rect 795 67 811 101
rect 845 67 861 101
rect 795 17 861 67
rect 895 101 933 135
rect 895 67 897 101
rect 931 67 933 101
rect 895 51 933 67
rect 967 169 1033 180
rect 967 135 983 169
rect 1017 135 1033 169
rect 967 101 1033 135
rect 967 67 983 101
rect 1017 67 1033 101
rect 967 17 1033 67
rect 1067 169 1127 196
rect 1067 135 1077 169
rect 1111 135 1127 169
rect 1067 101 1127 135
rect 1067 67 1077 101
rect 1111 67 1127 101
rect 1067 51 1127 67
rect 1165 169 1231 180
rect 1165 135 1181 169
rect 1215 135 1231 169
rect 1165 101 1231 135
rect 1165 67 1181 101
rect 1215 67 1231 101
rect 1165 17 1231 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 1071 63 1105
rect 121 1071 155 1105
rect 213 1071 247 1105
rect 305 1071 339 1105
rect 397 1071 431 1105
rect 489 1071 523 1105
rect 581 1071 615 1105
rect 673 1071 707 1105
rect 765 1071 799 1105
rect 857 1071 891 1105
rect 949 1071 983 1105
rect 1041 1071 1075 1105
rect 1133 1071 1167 1105
rect 1225 1071 1259 1105
rect 28 725 29 731
rect 29 725 62 731
rect 28 697 62 725
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 284 423 318 457
rect 356 423 390 457
rect 428 424 462 457
rect 428 423 462 424
rect 1214 725 1225 731
rect 1225 725 1248 731
rect 1214 697 1248 725
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 1105 1288 1136
rect 0 1071 29 1105
rect 63 1071 121 1105
rect 155 1071 213 1105
rect 247 1071 305 1105
rect 339 1071 397 1105
rect 431 1071 489 1105
rect 523 1071 581 1105
rect 615 1071 673 1105
rect 707 1071 765 1105
rect 799 1071 857 1105
rect 891 1071 949 1105
rect 983 1071 1041 1105
rect 1075 1071 1133 1105
rect 1167 1071 1225 1105
rect 1259 1071 1288 1105
rect 0 1040 1288 1071
rect 16 731 74 737
rect 16 728 28 731
rect 14 700 28 728
rect 16 697 28 700
rect 62 728 74 731
rect 1202 731 1260 737
rect 1202 728 1214 731
rect 62 700 1214 728
rect 62 697 74 700
rect 16 691 74 697
rect 1202 697 1214 700
rect 1248 697 1260 731
rect 1202 691 1260 697
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 272 457 474 463
rect 272 456 284 457
rect 14 428 284 456
rect 272 423 284 428
rect 318 423 356 457
rect 390 423 428 457
rect 462 456 474 457
rect 462 428 1274 456
rect 462 423 474 428
rect 272 417 474 423
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
rlabel comment s 0 0 0 0 4 lpflow_lsbuf_lh_hl_isowell_tap_2
flabel comment s 821 764 821 764 0 FreeSans 200 90 0 0 no_jumper_check
flabel metal1 s 66 1071 94 1105 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 98 700 125 728 0 FreeSans 200 0 0 0 VPB
port 3 nsew power bidirectional
flabel metal1 s 82 -11 116 23 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 87 428 99 456 0 FreeSans 200 0 0 0 VPWRIN
port 4 nsew power bidirectional abutment
flabel metal1 s 0 496 1248 544 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 607 268 641 302 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 1087 268 1121 302 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 1087 194 1121 228 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
rlabel locali s 1213 926 1271 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 889 903 991 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 715 903 753 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 529 903 581 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 17 926 75 1071 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 0 1071 1288 1105 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1288 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 1040 1288 1136 1 VGND
port 2 nsew ground bidirectional abutment
rlabel locali s 1181 322 1215 527 1 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 561 1024 748 1 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 527 1288 561 1 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 978 325 1024 527 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 272 456 474 463 1 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 272 417 474 428 1 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 14 428 1274 456 1 VPWRIN
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 1088
string GDS_END 1557648
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1544374
string LEFclass CORE WELLTAP
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
