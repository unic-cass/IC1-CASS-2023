* NGSPICE file created from wb_buttons_leds.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt wb_buttons_leds buttons clk i_wb_addr[0] i_wb_addr[10] i_wb_addr[11] i_wb_addr[12]
+ i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16] i_wb_addr[17] i_wb_addr[18]
+ i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21] i_wb_addr[22] i_wb_addr[23]
+ i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27] i_wb_addr[28] i_wb_addr[29]
+ i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3] i_wb_addr[4] i_wb_addr[5]
+ i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc i_wb_data[0] i_wb_data[10]
+ i_wb_data[11] i_wb_data[12] i_wb_data[13] i_wb_data[14] i_wb_data[15] i_wb_data[16]
+ i_wb_data[17] i_wb_data[18] i_wb_data[19] i_wb_data[1] i_wb_data[20] i_wb_data[21]
+ i_wb_data[22] i_wb_data[23] i_wb_data[24] i_wb_data[25] i_wb_data[26] i_wb_data[27]
+ i_wb_data[28] i_wb_data[29] i_wb_data[2] i_wb_data[30] i_wb_data[31] i_wb_data[3]
+ i_wb_data[4] i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8] i_wb_data[9] i_wb_stb
+ i_wb_we led_enb[0] led_enb[10] led_enb[11] led_enb[1] led_enb[2] led_enb[3] led_enb[4]
+ led_enb[5] led_enb[6] led_enb[7] led_enb[8] led_enb[9] leds[0] leds[10] leds[11]
+ leds[1] leds[2] leds[3] leds[4] leds[5] leds[6] leds[7] leds[8] leds[9] o_wb_ack
+ o_wb_data[0] o_wb_data[10] o_wb_data[11] o_wb_data[12] o_wb_data[13] o_wb_data[14]
+ o_wb_data[15] o_wb_data[16] o_wb_data[17] o_wb_data[18] o_wb_data[19] o_wb_data[1]
+ o_wb_data[20] o_wb_data[21] o_wb_data[22] o_wb_data[23] o_wb_data[24] o_wb_data[25]
+ o_wb_data[26] o_wb_data[27] o_wb_data[28] o_wb_data[29] o_wb_data[2] o_wb_data[30]
+ o_wb_data[31] o_wb_data[3] o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7] o_wb_data[8]
+ o_wb_data[9] o_wb_stall reset vccd1 vssd1
X_09671_ _09631_/Y _09666_/B _09674_/B _09670_/X vssd1 vssd1 vccd1 vccd1 _09819_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_94_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09105_ _12770_/A _11920_/B _09172_/B _17466_/D vssd1 vssd1 vccd1 vccd1 _09106_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_175_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09036_ _17081_/A _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__o21ba_4
XFILLER_191_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout820 _12465_/B vssd1 vssd1 vccd1 vccd1 _12770_/D sky130_fd_sc_hd__buf_12
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout831 _10962_/B vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__buf_12
X_09938_ _10067_/A _09803_/B _09803_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__a21oi_1
Xfanout842 _14906_/A vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__buf_6
Xfanout853 _10963_/D vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__buf_2
Xfanout864 _11377_/C vssd1 vssd1 vccd1 vccd1 _11563_/D sky130_fd_sc_hd__buf_6
Xfanout875 _11377_/D vssd1 vssd1 vccd1 vccd1 _11629_/C sky130_fd_sc_hd__buf_4
Xfanout886 _17480_/Q vssd1 vssd1 vccd1 vccd1 _15402_/A sky130_fd_sc_hd__clkbuf_16
X_09869_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09869_/X sky130_fd_sc_hd__a21o_2
Xfanout897 _10560_/D vssd1 vssd1 vccd1 vccd1 _10062_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11900_ _12107_/A _11900_/B _12258_/B _12090_/B vssd1 vssd1 vccd1 vccd1 _11901_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12880_ _12881_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _13040_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _12031_/A _11831_/B vssd1 vssd1 vccd1 vccd1 _11831_/Y sky130_fd_sc_hd__nand2_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14599_/B _14708_/D vssd1 vssd1 vccd1 vccd1 _14679_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11762_ _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__and2_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13501_ _13501_/A _13501_/B vssd1 vssd1 vccd1 vccd1 _13503_/A sky130_fd_sc_hd__nor2_1
X_10713_ _10713_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10715_/C sky130_fd_sc_hd__xnor2_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _15457_/C _12864_/A _14840_/A vssd1 vssd1 vccd1 vccd1 _14481_/X sky130_fd_sc_hd__mux2_4
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _11693_/A vssd1 vssd1 vccd1 vccd1 _11693_/Y sky130_fd_sc_hd__inv_2
X_16220_ _08776_/C _17075_/A2 _16218_/X _16219_/Y vssd1 vssd1 vccd1 vccd1 _16221_/A
+ sky130_fd_sc_hd__a211o_1
X_13432_ _13431_/A _13431_/B _13431_/C vssd1 vssd1 vccd1 vccd1 _13443_/B sky130_fd_sc_hd__o21ai_4
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _10644_/A _10649_/A _10644_/C vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__or3_4
XFILLER_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _16040_/B _16245_/A _16149_/X vssd1 vssd1 vccd1 vccd1 _16153_/A sky130_fd_sc_hd__a21oi_4
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13363_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _13364_/B sky130_fd_sc_hd__and2_1
X_10575_ _10567_/A _10572_/A _10573_/X _10574_/Y vssd1 vssd1 vccd1 vccd1 _10575_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_166_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ _15131_/A _15102_/B vssd1 vssd1 vccd1 vccd1 _15102_/Y sky130_fd_sc_hd__nand2_1
X_12314_ _12314_/A _12314_/B vssd1 vssd1 vccd1 vccd1 _12316_/C sky130_fd_sc_hd__nand2_2
X_16082_ _15577_/Y _16361_/A _15954_/A vssd1 vssd1 vccd1 vccd1 _16082_/X sky130_fd_sc_hd__o21a_1
X_13294_ _13295_/A _13295_/B _13295_/C vssd1 vssd1 vccd1 vccd1 _13308_/A sky130_fd_sc_hd__a21o_4
XFILLER_177_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15033_ _12025_/B _11813_/B _09350_/B _12597_/B _12060_/S _15095_/B vssd1 vssd1 vccd1
+ vccd1 _15034_/B sky130_fd_sc_hd__mux4_1
XFILLER_170_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12245_ _12245_/A _12245_/B vssd1 vssd1 vccd1 vccd1 _12247_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12176_ _12176_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__nand2_2
XFILLER_122_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11127_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11130_/C sky130_fd_sc_hd__nand2_2
XFILLER_150_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16984_ _16991_/A _17040_/A _16984_/C vssd1 vssd1 vccd1 vccd1 _16986_/B sky130_fd_sc_hd__and3_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15935_ _15935_/A _15935_/B vssd1 vssd1 vccd1 vccd1 _15937_/B sky130_fd_sc_hd__xnor2_1
X_11058_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11059_/C sky130_fd_sc_hd__xnor2_4
XFILLER_7_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10009_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__nand3_1
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15866_ _15866_/A _15866_/B _15866_/C vssd1 vssd1 vccd1 vccd1 _15867_/B sky130_fd_sc_hd__or3_1
XFILLER_92_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17605_ fanout940/X _17605_/D vssd1 vssd1 vccd1 vccd1 _17605_/Q sky130_fd_sc_hd__dfxtp_1
X_14817_ _14775_/X _14816_/X _12560_/A vssd1 vssd1 vccd1 vccd1 _16577_/A sky130_fd_sc_hd__a21bo_1
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15797_ _15797_/A _15797_/B vssd1 vssd1 vccd1 vccd1 _15797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17536_ fanout933/X _17536_/D vssd1 vssd1 vccd1 vccd1 _17536_/Q sky130_fd_sc_hd__dfxtp_1
X_14748_ _14748_/A _14748_/B vssd1 vssd1 vccd1 vccd1 _14750_/B sky130_fd_sc_hd__or2_1
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17467_ fanout928/X _17467_/D vssd1 vssd1 vccd1 vccd1 _17467_/Q sky130_fd_sc_hd__dfxtp_1
X_14679_ _14649_/A _14679_/B vssd1 vssd1 vccd1 vccd1 _14680_/C sky130_fd_sc_hd__nand2b_2
XFILLER_32_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16418_ _16419_/A _16419_/B vssd1 vssd1 vccd1 vccd1 _16519_/B sky130_fd_sc_hd__or2_2
X_17398_ input44/X _17422_/A2 _17397_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17527_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16349_ _16266_/A _16266_/B _16267_/Y vssd1 vssd1 vccd1 vccd1 _16363_/B sky130_fd_sc_hd__a21bo_1
XFILLER_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout127 _17270_/A2 vssd1 vssd1 vccd1 vccd1 _17231_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout149 _14912_/Y vssd1 vssd1 vccd1 vccd1 _15097_/A sky130_fd_sc_hd__buf_4
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _09723_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09725_/C sky130_fd_sc_hd__or2_4
XFILLER_80_1062 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09654_ _09655_/A _09653_/Y _09928_/C _09654_/D vssd1 vssd1 vccd1 vccd1 _09784_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _11900_/B _09892_/D _10036_/D _09584_/A vssd1 vssd1 vccd1 vccd1 _09585_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _10694_/A _10694_/B _10479_/B _10360_/D vssd1 vssd1 vccd1 vccd1 _10374_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09019_ _08905_/A _08905_/C _08905_/B vssd1 vssd1 vccd1 vccd1 _09051_/B sky130_fd_sc_hd__a21o_2
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10291_ _10971_/A _10745_/D _10743_/C _10525_/A vssd1 vssd1 vccd1 vccd1 _10291_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_117_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12030_ _17363_/A _09350_/B _14948_/B vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__a21o_1
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout650 _12025_/B vssd1 vssd1 vccd1 vccd1 _12734_/C sky130_fd_sc_hd__buf_6
Xfanout661 _09654_/D vssd1 vssd1 vccd1 vccd1 _11808_/B sky130_fd_sc_hd__buf_4
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout672 fanout676/X vssd1 vssd1 vccd1 vccd1 _14153_/C sky130_fd_sc_hd__buf_8
X_13981_ _13982_/A _13982_/B vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__and2b_1
Xfanout683 fanout686/X vssd1 vssd1 vccd1 vccd1 _14063_/C sky130_fd_sc_hd__buf_6
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout694 _17500_/Q vssd1 vssd1 vccd1 vccd1 _16722_/A sky130_fd_sc_hd__buf_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15720_ _11700_/Y _16389_/A _15701_/X _15719_/X vssd1 vssd1 vccd1 vccd1 _15720_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12932_ _13117_/B _12932_/B vssd1 vssd1 vccd1 vccd1 _12933_/C sky130_fd_sc_hd__nand2_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15651_ _15651_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15742_/B sky130_fd_sc_hd__xnor2_4
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12863_ _12861_/X _12862_/X _17369_/A vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__mux2_2
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14601_/A _14601_/B _14601_/C vssd1 vssd1 vccd1 vccd1 _14646_/A sky130_fd_sc_hd__o21ai_2
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11814_ _14982_/B _14981_/B _14912_/B vssd1 vssd1 vccd1 vccd1 _11814_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15582_/A _15582_/B vssd1 vssd1 vccd1 vccd1 _15584_/B sky130_fd_sc_hd__xnor2_4
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12794_/A _12794_/B vssd1 vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__nor2_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ input39/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__or3_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14533_/A _14533_/B _14533_/C vssd1 vssd1 vccd1 vccd1 _14534_/B sky130_fd_sc_hd__and3_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11747_/B sky130_fd_sc_hd__xnor2_1
XFILLER_159_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17252_ _17593_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17252_/X sky130_fd_sc_hd__a21o_1
X_14464_ _14463_/B _14463_/C _14463_/A vssd1 vssd1 vccd1 vccd1 _14465_/B sky130_fd_sc_hd__a21o_1
X_11676_ _11676_/A _15011_/A vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__nor2_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16203_ _16203_/A _16203_/B _16099_/X vssd1 vssd1 vccd1 vccd1 _16203_/X sky130_fd_sc_hd__or3b_4
X_13415_ _13415_/A _13415_/B vssd1 vssd1 vccd1 vccd1 _13417_/C sky130_fd_sc_hd__nor2_2
XFILLER_179_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _10713_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__and2_2
X_17183_ input14/X input3/X vssd1 vssd1 vccd1 vccd1 _17428_/C sky130_fd_sc_hd__nor2_8
X_14395_ _14396_/A _14396_/B vssd1 vssd1 vccd1 vccd1 _14395_/Y sky130_fd_sc_hd__nor2_4
XFILLER_183_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16134_ _16136_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _16234_/C sky130_fd_sc_hd__nand2_1
XFILLER_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13346_ _13346_/A _13346_/B _13346_/C vssd1 vssd1 vccd1 vccd1 _13347_/B sky130_fd_sc_hd__and3_1
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10558_ _10559_/A _11370_/C _10559_/B _10560_/A vssd1 vssd1 vccd1 vccd1 _10561_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_182_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16065_ _16171_/A _16814_/B vssd1 vssd1 vccd1 vccd1 _16066_/B sky130_fd_sc_hd__nand2_2
XFILLER_142_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13277_ _17371_/A _13516_/S _12218_/A _13276_/Y _08718_/A vssd1 vssd1 vccd1 vccd1
+ _13277_/X sky130_fd_sc_hd__a311o_1
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10489_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__xnor2_2
X_15016_ _17164_/C _15001_/X _15015_/X vssd1 vssd1 vccd1 vccd1 _15016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12228_ _11824_/Y _11852_/B _15095_/B vssd1 vssd1 vccd1 vccd1 _12229_/C sky130_fd_sc_hd__mux2_2
XFILLER_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12159_ _12488_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _12161_/C sky130_fd_sc_hd__nand2_1
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16967_ _16858_/Y _16914_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16967_/X sky130_fd_sc_hd__o21ba_1
XFILLER_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15918_ _15918_/A _16226_/B _16743_/C _17043_/B vssd1 vssd1 vccd1 vccd1 _15918_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16898_ _16897_/A _16897_/B _16897_/C vssd1 vssd1 vccd1 vccd1 _16900_/B sky130_fd_sc_hd__o21ai_2
XFILLER_92_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15849_ _16165_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _15850_/B sky130_fd_sc_hd__nand2_2
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09370_ _09370_/A _09370_/B _09370_/C vssd1 vssd1 vccd1 vccd1 _09387_/B sky130_fd_sc_hd__nand3_2
XFILLER_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17519_ fanout931/X _17519_/D vssd1 vssd1 vccd1 vccd1 _17519_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09706_ _09706_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09709_/A sky130_fd_sc_hd__nor2_4
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwb_buttons_leds_957 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_957/HI led_enb[10] sky130_fd_sc_hd__conb_1
X_09637_ _09942_/A _09637_/B _11920_/D _09944_/D vssd1 vssd1 vccd1 vccd1 _09640_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _10255_/A _10791_/C vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__nand2_8
XFILLER_167_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _09620_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__nand2_4
X_11530_ _11534_/B _11530_/B _11530_/C vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__and3_2
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11461_ _11460_/B _11461_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__and2b_2
XFILLER_183_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13200_ _13369_/A _13200_/B vssd1 vssd1 vccd1 vccd1 _13202_/C sky130_fd_sc_hd__nor2_2
X_10412_ _10525_/A _10971_/A _10412_/C _10640_/D vssd1 vssd1 vccd1 vccd1 _10415_/A
+ sky130_fd_sc_hd__and4_2
X_14180_ _14180_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14181_/C sky130_fd_sc_hd__xnor2_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11392_ _11393_/B _11393_/C _11393_/A vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__o21ai_2
XFILLER_178_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13131_ _12956_/A _12960_/A _13264_/A _13130_/Y vssd1 vssd1 vccd1 vccd1 _13264_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10343_ _10342_/A _10342_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10343_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10274_ _14785_/A _10013_/B _10272_/X _10269_/X _10145_/B vssd1 vssd1 vccd1 vccd1
+ _10276_/B sky130_fd_sc_hd__a32o_2
X_13062_ _13061_/A _13061_/B _13061_/C vssd1 vssd1 vccd1 vccd1 _13063_/B sky130_fd_sc_hd__a21o_1
XFILLER_140_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12013_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12014_/B sky130_fd_sc_hd__and2_1
XFILLER_132_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16821_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16897_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout480 _15262_/A vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__buf_6
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout491 _12907_/A vssd1 vssd1 vccd1 vccd1 _11902_/A sky130_fd_sc_hd__buf_6
XFILLER_111_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16752_ _16751_/A _16751_/B _16751_/C vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__a21oi_2
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13964_ _13964_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__xnor2_2
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15703_ _15703_/A _15796_/B _15262_/A vssd1 vssd1 vccd1 vccd1 _15705_/B sky130_fd_sc_hd__or3b_4
X_12915_ _12915_/A _12915_/B _12915_/C vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__and3_1
X_16683_ _16683_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16684_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13895_ _13895_/A _13895_/B _13895_/C _14063_/C vssd1 vssd1 vccd1 vccd1 _13896_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15634_ _16917_/A _15621_/Y _15633_/Y _15613_/Y vssd1 vssd1 vccd1 vccd1 _15634_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ _12844_/X _12845_/X _13838_/S vssd1 vssd1 vccd1 vccd1 _12847_/B sky130_fd_sc_hd__mux2_1
XFILLER_181_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _16136_/B _16533_/A _16695_/A _15647_/A vssd1 vssd1 vccd1 vccd1 _15568_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12777_ _12778_/A _12778_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12779_/A sky130_fd_sc_hd__a21oi_1
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17304_/A1 _17328_/A2 _17303_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17481_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14516_ _14518_/A _14518_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14519_/B sky130_fd_sc_hd__a21o_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11728_ _11725_/A _11725_/B _11725_/C vssd1 vssd1 vccd1 vccd1 _11729_/C sky130_fd_sc_hd__a21oi_4
XFILLER_147_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ _15496_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__nor2_4
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17235_ _17555_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__and2_1
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14447_ _14508_/A _14446_/C _14446_/A vssd1 vssd1 vccd1 vccd1 _14459_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11659_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__xnor2_2
XFILLER_128_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ _17166_/A _17166_/B _17166_/C vssd1 vssd1 vccd1 vccd1 _17166_/X sky130_fd_sc_hd__and3_1
X_14378_ _14378_/A _14378_/B _14378_/C vssd1 vssd1 vccd1 vccd1 _14379_/B sky130_fd_sc_hd__and3_1
XFILLER_155_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16117_ _16011_/A _14922_/S _17164_/D _16012_/S vssd1 vssd1 vccd1 vccd1 _16117_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_171_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13329_ _13329_/A _13329_/B _13329_/C vssd1 vssd1 vccd1 vccd1 _13330_/B sky130_fd_sc_hd__nand3_4
XFILLER_192_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17097_ _17096_/A _17096_/B _17096_/C vssd1 vssd1 vccd1 vccd1 _17097_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _16048_/A _16048_/B vssd1 vssd1 vccd1 vccd1 _16051_/A sky130_fd_sc_hd__xnor2_2
XFILLER_89_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _08844_/X _08908_/A _08868_/X _08869_/Y vssd1 vssd1 vccd1 vccd1 _08873_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09422_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__nand2b_2
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09353_ _09353_/A _09491_/A vssd1 vssd1 vccd1 vccd1 _09355_/B sky130_fd_sc_hd__nor2_4
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _12258_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__and2_2
XFILLER_193_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08999_ _08999_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__nor2_4
XFILLER_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _11010_/B _10961_/B _11043_/B vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__or3_4
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12700_ _16011_/B _15095_/B _12700_/C _12700_/D vssd1 vssd1 vccd1 vccd1 _13628_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_141_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13680_ _13680_/A _13680_/B _13680_/C vssd1 vssd1 vccd1 vccd1 _13681_/B sky130_fd_sc_hd__nor3_1
XFILLER_71_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10892_ _11148_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10893_/C sky130_fd_sc_hd__and2_2
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12631_ _12631_/A _12631_/B _12631_/C vssd1 vssd1 vccd1 vccd1 _12631_/Y sky130_fd_sc_hd__nor3_4
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15350_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15352_/B sky130_fd_sc_hd__xnor2_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _12561_/A _12561_/B _12561_/C vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__o21ai_2
X_14301_ _14680_/A _14599_/B _14545_/D _14485_/D vssd1 vssd1 vccd1 vccd1 _14302_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11513_ _11475_/A _11475_/C _11475_/B vssd1 vssd1 vccd1 vccd1 _11514_/C sky130_fd_sc_hd__a21oi_4
X_15281_ _15281_/A _15281_/B vssd1 vssd1 vccd1 vccd1 _15283_/B sky130_fd_sc_hd__xnor2_4
XFILLER_184_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12493_ _12492_/A _12492_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12494_/B sky130_fd_sc_hd__o21a_1
XFILLER_156_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17020_ _16966_/B _16969_/B _16966_/A vssd1 vssd1 vccd1 vccd1 _17066_/B sky130_fd_sc_hd__o21bai_2
X_14232_ _14232_/A _14232_/B vssd1 vssd1 vccd1 vccd1 _14235_/A sky130_fd_sc_hd__xor2_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11444_ _11444_/A _11444_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11444_/Y sky130_fd_sc_hd__nand3_4
XFILLER_184_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14163_ _14237_/A _14237_/B vssd1 vssd1 vccd1 vccd1 _14165_/B sky130_fd_sc_hd__xor2_2
XFILLER_171_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11375_ _11553_/B _11518_/C _11325_/A _11324_/D vssd1 vssd1 vccd1 vccd1 _11376_/C
+ sky130_fd_sc_hd__a22o_2
XFILLER_153_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ _13114_/A _13114_/B vssd1 vssd1 vccd1 vccd1 _13115_/B sky130_fd_sc_hd__nor2_1
XFILLER_180_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _10559_/A _10360_/D _10326_/C vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__nand3_4
XFILLER_124_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14094_ _14254_/A _14175_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14200_/B sky130_fd_sc_hd__and3_1
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13046_/A _13046_/B _13046_/C vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__a21o_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10372_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10188_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10188_/Y sky130_fd_sc_hd__nand3_4
XFILLER_78_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16804_ _15794_/A _16795_/Y _16797_/X _17169_/A1 _16803_/X vssd1 vssd1 vccd1 vccd1
+ _16804_/X sky130_fd_sc_hd__o221a_2
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14996_ _09509_/B _10736_/C _10738_/D _10013_/B _10430_/A _14982_/A vssd1 vssd1 vccd1
+ vccd1 _14998_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13947_ _13948_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _13947_/Y sky130_fd_sc_hd__nand2_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16735_ _16735_/A _16735_/B vssd1 vssd1 vccd1 vccd1 _16735_/Y sky130_fd_sc_hd__nor2_1
XFILLER_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16666_ _16667_/A _16938_/D vssd1 vssd1 vccd1 vccd1 _16670_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _13878_/A _13878_/B vssd1 vssd1 vccd1 vccd1 _13880_/A sky130_fd_sc_hd__nor2_2
X_15617_ _15617_/A _15891_/B _15262_/B vssd1 vssd1 vccd1 vccd1 _15618_/B sky130_fd_sc_hd__or3b_1
X_12829_ _12826_/A _12827_/Y _12676_/A _12677_/Y vssd1 vssd1 vccd1 vccd1 _12829_/Y
+ sky130_fd_sc_hd__a211oi_4
X_16597_ _16597_/A _16597_/B vssd1 vssd1 vccd1 vccd1 _16600_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ _15548_/A vssd1 vssd1 vccd1 vccd1 _17552_/D sky130_fd_sc_hd__clkinv_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15479_ _15564_/A _15479_/B vssd1 vssd1 vccd1 vccd1 _15481_/B sky130_fd_sc_hd__nand2_4
XFILLER_147_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _17440_/Q _17233_/A2 _17216_/X _17217_/X _17372_/C1 vssd1 vssd1 vccd1 vccd1
+ _17440_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17149_ _17119_/B _17086_/A _17038_/C _16315_/A vssd1 vssd1 vccd1 vccd1 _17149_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _09964_/A _09962_/X _09923_/A _09957_/A vssd1 vssd1 vccd1 vccd1 _10091_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_157_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08922_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08853_ _11895_/A _12270_/B _12734_/C _12734_/D vssd1 vssd1 vccd1 vccd1 _08854_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _12088_/A _12088_/B _11870_/B _11867_/C vssd1 vssd1 vccd1 vccd1 _08798_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_85_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09405_ _09409_/C _09647_/B _09268_/A _09266_/Y vssd1 vssd1 vccd1 vccd1 _09411_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_38_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _09344_/A _09316_/X _09334_/A _09335_/Y vssd1 vssd1 vccd1 vccd1 _09339_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ _09268_/A _09266_/Y _09409_/C _09647_/B vssd1 vssd1 vccd1 vccd1 _09411_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09198_ _12166_/A _12340_/B _09198_/C vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__nand3_2
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11162_/C sky130_fd_sc_hd__xnor2_2
XFILLER_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10111_ _10112_/A _10110_/Y _10366_/A _17468_/D vssd1 vssd1 vccd1 vccd1 _10234_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11091_ _11080_/A _11080_/C _11080_/D _11080_/B vssd1 vssd1 vccd1 vccd1 _11145_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_96_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10042_ _10042_/A _10046_/A _10042_/C vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__or3_2
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14850_ _15381_/A _14906_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__and3_1
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _13801_/A _13801_/B vssd1 vssd1 vccd1 vccd1 _13803_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14781_ _16809_/A _15898_/A vssd1 vssd1 vccd1 vccd1 _15895_/B sky130_fd_sc_hd__or2_2
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11993_ _11993_/A _12155_/B _11993_/C vssd1 vssd1 vccd1 vccd1 _12197_/A sky130_fd_sc_hd__nor3_4
XFILLER_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16520_ _16625_/A _16520_/B vssd1 vssd1 vccd1 vccd1 _16522_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13732_ _13936_/A _13732_/B vssd1 vssd1 vccd1 vccd1 _13828_/B sky130_fd_sc_hd__or2_1
XFILLER_28_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ _10995_/B _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10945_/B sky130_fd_sc_hd__o21ai_1
XFILLER_72_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _16354_/B _16356_/B _16354_/A vssd1 vssd1 vccd1 vccd1 _16453_/B sky130_fd_sc_hd__o21ba_2
XFILLER_56_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13663_ _14050_/B _13764_/D _13664_/D _14050_/A vssd1 vssd1 vccd1 vccd1 _13665_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ _11266_/A _11122_/B _11391_/B _11480_/C vssd1 vssd1 vccd1 vccd1 _10878_/A
+ sky130_fd_sc_hd__and4_1
X_15402_ _15402_/A _15402_/B _16695_/A vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__and3_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12611_/X _12612_/Y _12458_/A _12458_/Y vssd1 vssd1 vccd1 vccd1 _12631_/B
+ sky130_fd_sc_hd__o211a_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _16382_/A _16382_/B vssd1 vssd1 vccd1 vccd1 _16562_/B sky130_fd_sc_hd__or2_1
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13594_ _13595_/A _13595_/B vssd1 vssd1 vccd1 vccd1 _13594_/X sky130_fd_sc_hd__and2b_2
XFILLER_185_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _15821_/A _16536_/A _15334_/A vssd1 vssd1 vccd1 vccd1 _15408_/B sky130_fd_sc_hd__and3_1
XFILLER_61_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12545_ _12543_/X _12544_/X _13838_/S vssd1 vssd1 vccd1 vccd1 _12545_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15264_ _15143_/X _15262_/X _15305_/C vssd1 vssd1 vccd1 vccd1 _16446_/A sky130_fd_sc_hd__a21bo_4
XFILLER_177_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12476_ _12476_/A _12476_/B _12476_/C vssd1 vssd1 vccd1 vccd1 _12477_/B sky130_fd_sc_hd__and3_1
X_17003_ _17003_/A _17003_/B _17003_/C vssd1 vssd1 vccd1 vccd1 _17004_/B sky130_fd_sc_hd__nand3_2
X_14215_ _14215_/A _14215_/B vssd1 vssd1 vccd1 vccd1 _14216_/B sky130_fd_sc_hd__nand2_2
XFILLER_8_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11427_ _11506_/A _11553_/A _11561_/D _15402_/A vssd1 vssd1 vccd1 vccd1 _11430_/A
+ sky130_fd_sc_hd__and4_2
XANTENNA_5 _17555_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _17063_/A _15171_/Y _15173_/Y _15194_/X vssd1 vssd1 vccd1 vccd1 _15195_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14146_ _14229_/B _14146_/B vssd1 vssd1 vccd1 vccd1 _14148_/B sky130_fd_sc_hd__nor2_2
XFILLER_153_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11358_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__nor2_2
XFILLER_180_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ _10431_/A _10309_/B _10309_/C vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__and3_2
XFILLER_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14077_ _14077_/A _14077_/B vssd1 vssd1 vccd1 vccd1 _14078_/B sky130_fd_sc_hd__or2_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11289_ _11348_/A _11253_/B _11351_/A vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__o21ai_4
X_13028_ _13643_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__nand2_4
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14979_ _15096_/S _14979_/B vssd1 vssd1 vccd1 vccd1 _14979_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16718_ _16715_/Y _16717_/Y _17131_/A vssd1 vssd1 vccd1 vccd1 _16718_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16649_ _16649_/A _16649_/B _16649_/C vssd1 vssd1 vccd1 vccd1 _16649_/X sky130_fd_sc_hd__and3_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09121_ _09015_/X _09017_/Y _09119_/A _09119_/Y vssd1 vssd1 vccd1 vccd1 _09122_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap263 _15141_/B vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__buf_4
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09954_ _10078_/A _10078_/B _09936_/A vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08905_ _08905_/A _08905_/B _08905_/C vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__nand3_4
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09885_/A _09885_/B _09885_/C vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__and3_2
XFILLER_106_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _12275_/A _12107_/B _12088_/C _12088_/D vssd1 vssd1 vccd1 vccd1 _08862_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08767_ _09025_/C _12166_/B _08754_/C _08754_/D vssd1 vssd1 vccd1 vccd1 _08768_/B
+ sky130_fd_sc_hd__a22oi_2
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10660_ _10660_/A _10757_/A vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__nor2_4
XFILLER_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09319_ _12592_/A _09748_/B _10311_/D _10308_/B vssd1 vssd1 vccd1 vccd1 _09328_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10591_ _10694_/A _10694_/B _17468_/D _17467_/D vssd1 vssd1 vccd1 vccd1 _10592_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12330_ _12498_/B _12330_/B vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__nand2_2
XFILLER_182_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__xnor2_4
XFILLER_108_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14000_ _14001_/A _14001_/B vssd1 vssd1 vccd1 vccd1 _14092_/A sky130_fd_sc_hd__nand2_1
X_11212_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__xnor2_4
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _12192_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12193_/C sky130_fd_sc_hd__xnor2_4
XFILLER_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11143_ _11144_/A _11146_/B _11143_/C _11143_/D vssd1 vssd1 vccd1 vccd1 _11237_/A
+ sky130_fd_sc_hd__nand4_4
Xoutput75 _17468_/Q vssd1 vssd1 vccd1 vccd1 leds[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput86 _17445_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[11] sky130_fd_sc_hd__clkbuf_2
Xoutput97 _17455_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[21] sky130_fd_sc_hd__clkbuf_2
X_15951_ _16165_/A _16355_/B vssd1 vssd1 vccd1 vccd1 _15953_/B sky130_fd_sc_hd__nand2_1
X_11074_ _11074_/A _11074_/B vssd1 vssd1 vccd1 vccd1 _11075_/C sky130_fd_sc_hd__nand2_2
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14902_ _15204_/A _16880_/A _16807_/A _17613_/Q vssd1 vssd1 vccd1 vccd1 _14967_/D
+ sky130_fd_sc_hd__or4b_2
X_10025_ _09865_/B _09975_/X _09991_/Y _10005_/X vssd1 vssd1 vccd1 vccd1 _10025_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15882_ _15883_/A _15883_/B _15881_/Y vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__o21bai_4
XFILLER_48_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14833_ _17476_/D _17477_/D vssd1 vssd1 vccd1 vccd1 _14933_/B sky130_fd_sc_hd__or2_4
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14764_ _14765_/A _17065_/A vssd1 vssd1 vccd1 vccd1 _14764_/Y sky130_fd_sc_hd__nor2_1
X_17552_ fanout934/X _17552_/D vssd1 vssd1 vccd1 vccd1 _17552_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11976_ _12174_/B _12174_/D _12129_/B _12174_/A vssd1 vssd1 vccd1 vccd1 _11978_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16503_ _16503_/A _16670_/A vssd1 vssd1 vccd1 vccd1 _16503_/Y sky130_fd_sc_hd__nand2_1
X_13715_ _13601_/A _13604_/A _13818_/A _13714_/Y vssd1 vssd1 vccd1 vccd1 _13818_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ _11074_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _10927_/X sky130_fd_sc_hd__or2_2
XFILLER_60_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17483_ fanout927/X _17483_/D vssd1 vssd1 vccd1 vccd1 _17483_/Q sky130_fd_sc_hd__dfxtp_4
X_14695_ _14723_/B _14695_/B vssd1 vssd1 vccd1 vccd1 _14699_/A sky130_fd_sc_hd__or2_2
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13646_ _13749_/A _13645_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__a21o_1
X_16434_ _16511_/B _16434_/B vssd1 vssd1 vccd1 vccd1 _16436_/B sky130_fd_sc_hd__or2_4
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10859_/B _10859_/C _10859_/A vssd1 vssd1 vccd1 vccd1 _10861_/A sky130_fd_sc_hd__a21o_1
XFILLER_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _16365_/A _16365_/B vssd1 vssd1 vccd1 vccd1 _16367_/B sky130_fd_sc_hd__or2_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A _13577_/B vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__nor2_1
X_10789_ _10899_/C _10897_/B _10901_/A _10787_/Y vssd1 vssd1 vccd1 vccd1 _10796_/B
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15316_ _15314_/A _15713_/B1 _14929_/X _14801_/B vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_185_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12528_ _12528_/A _12528_/B _12528_/C vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__nor3_4
X_16296_ _16389_/A _16296_/B vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__nand2_2
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _14848_/B _15116_/B _15110_/B _14848_/A vssd1 vssd1 vccd1 vccd1 _15248_/B
+ sky130_fd_sc_hd__a31o_1
X_12459_ _12267_/Y _12290_/X _12457_/X _12458_/Y vssd1 vssd1 vccd1 vccd1 _12481_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15178_ _15174_/Y _15175_/X _15176_/Y _15177_/Y _15309_/B vssd1 vssd1 vccd1 vccd1
+ _15178_/X sky130_fd_sc_hd__a311o_1
XFILLER_119_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ _08718_/A _14127_/X _14128_/X vssd1 vssd1 vccd1 vccd1 _14129_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_98_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout309 _08731_/A vssd1 vssd1 vccd1 vccd1 _15143_/A sky130_fd_sc_hd__buf_6
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09670_ _09530_/X _09541_/X _09668_/A _09668_/Y vssd1 vssd1 vccd1 vccd1 _09670_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09104_ _11920_/B _09172_/B _17466_/D _12770_/A vssd1 vssd1 vccd1 vccd1 _09106_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ _09048_/B _09048_/C _09048_/A vssd1 vssd1 vccd1 vccd1 _09050_/A sky130_fd_sc_hd__a21o_2
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout810 _12923_/D vssd1 vssd1 vccd1 vccd1 _12338_/C sky130_fd_sc_hd__buf_12
XFILLER_120_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout821 _10920_/B vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__buf_8
Xfanout832 _17485_/Q vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__buf_12
X_09937_ _10560_/B _09937_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__nand2_2
Xfanout843 _10963_/C vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__buf_8
XFILLER_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout854 _14906_/B vssd1 vssd1 vccd1 vccd1 _11561_/C sky130_fd_sc_hd__buf_8
XFILLER_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout865 _17306_/A1 vssd1 vssd1 vccd1 vccd1 _11377_/C sky130_fd_sc_hd__buf_8
Xfanout876 _11377_/D vssd1 vssd1 vccd1 vccd1 _11561_/D sky130_fd_sc_hd__buf_6
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09868_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09870_/C sky130_fd_sc_hd__or2_2
Xfanout887 _10321_/C vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__buf_8
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout898 _10559_/B vssd1 vssd1 vccd1 vccd1 _10560_/D sky130_fd_sc_hd__buf_8
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _12258_/A _11881_/D _08798_/A _08786_/Y vssd1 vssd1 vccd1 vccd1 _08821_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09801_/B _09798_/Y _10062_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _09941_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_46_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _12923_/D _12770_/D _11839_/S vssd1 vssd1 vccd1 vccd1 _11831_/B sky130_fd_sc_hd__mux2_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11756_/A _11755_/B _11759_/A vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__a21o_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A _13500_/B _13500_/C vssd1 vssd1 vccd1 vccd1 _13501_/B sky130_fd_sc_hd__nor3_1
X_10712_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _10712_/X sky130_fd_sc_hd__or2_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14763_/S _14478_/X _14479_/Y _14423_/Y vssd1 vssd1 vccd1 vccd1 _17598_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _15524_/C _11692_/B _11670_/C vssd1 vssd1 vccd1 vccd1 _11693_/A sky130_fd_sc_hd__or3b_1
XFILLER_186_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ _13431_/A _13431_/B _13431_/C vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__or3_2
XFILLER_186_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10643_ _10644_/A _10644_/C vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__nor2_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16150_ _16667_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16245_/A sky130_fd_sc_hd__nor2_4
XFILLER_167_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13362_ _13363_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__nor2_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10574_ _10458_/X _10472_/Y _10557_/X _10572_/X vssd1 vssd1 vccd1 vccd1 _10574_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15101_ _12077_/C _15101_/A1 _12245_/B _12021_/B _14942_/A _14982_/A vssd1 vssd1
+ vccd1 vccd1 _15102_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _12312_/A _12312_/B _12312_/C vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__a21o_1
XFILLER_182_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16081_ _16081_/A _16081_/B vssd1 vssd1 vccd1 vccd1 _16089_/A sky130_fd_sc_hd__nand2_4
XFILLER_181_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13293_ _13411_/B _13293_/B vssd1 vssd1 vccd1 vccd1 _13295_/C sky130_fd_sc_hd__nand2_1
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15032_ _12700_/C _12032_/Y _15100_/A _15038_/A vssd1 vssd1 vccd1 vccd1 _16011_/C
+ sky130_fd_sc_hd__o211ai_4
X_12244_ _12244_/A _12429_/A vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__or2_1
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12175_ _12175_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12177_/A sky130_fd_sc_hd__nor2_1
XFILLER_111_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11126_ _11126_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11257_/B sky130_fd_sc_hd__xnor2_4
XFILLER_68_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16983_ _16983_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _16984_/C sky130_fd_sc_hd__nand2_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15934_ _16595_/A _16041_/B vssd1 vssd1 vccd1 vccd1 _15935_/B sky130_fd_sc_hd__nor2_1
X_11057_ _11057_/A _11057_/B _11057_/C vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__nand3_4
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__a21o_1
XFILLER_190_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15865_ _15866_/A _15866_/B _15866_/C vssd1 vssd1 vccd1 vccd1 _15867_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17604_ fanout942/X _17604_/D vssd1 vssd1 vccd1 vccd1 _17604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14816_ _16397_/B _16398_/A _12235_/C vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__a21o_1
XFILLER_92_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _15811_/A _15796_/B _16136_/A vssd1 vssd1 vccd1 vccd1 _15797_/B sky130_fd_sc_hd__or3b_1
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17535_ fanout933/X _17535_/D vssd1 vssd1 vccd1 vccd1 _17535_/Q sky130_fd_sc_hd__dfxtp_2
X_14747_ _14747_/A _14747_/B _14747_/C vssd1 vssd1 vccd1 vccd1 _14748_/B sky130_fd_sc_hd__and3_1
X_11959_ _11958_/A _11958_/B _11958_/C vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14678_ _14678_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__nor2_4
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17466_ fanout928/X _17466_/D vssd1 vssd1 vccd1 vccd1 _17466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16417_ _16417_/A _16519_/A vssd1 vssd1 vccd1 vccd1 _16419_/B sky130_fd_sc_hd__nand2_1
X_13629_ _14210_/B _13627_/X _13628_/Y _12401_/A _12854_/Y vssd1 vssd1 vccd1 vccd1
+ _13629_/X sky130_fd_sc_hd__o221a_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17397_ _17397_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17397_/X sky130_fd_sc_hd__or2_1
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16348_ _16462_/A _16348_/B vssd1 vssd1 vccd1 vccd1 _16367_/A sky130_fd_sc_hd__nand2b_4
XFILLER_160_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16279_ _16279_/A _16279_/B _16279_/C vssd1 vssd1 vccd1 vccd1 _16280_/B sky130_fd_sc_hd__nor3_2
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout128 _17288_/A2 vssd1 vssd1 vccd1 vccd1 _17291_/A2 sky130_fd_sc_hd__buf_4
XFILLER_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout139 _16127_/B vssd1 vssd1 vccd1 vccd1 _16226_/C sky130_fd_sc_hd__buf_12
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09722_ _09722_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09653_ _09926_/A _09926_/B _14982_/B vssd1 vssd1 vccd1 vccd1 _09653_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09584_ _09584_/A _11900_/B _09892_/D _10036_/D vssd1 vssd1 vccd1 vccd1 _09587_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_70_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09018_ _08930_/A _08930_/C _08930_/B vssd1 vssd1 vccd1 vccd1 _09018_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_191_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ _14786_/A _10971_/A _10745_/D _10412_/C vssd1 vssd1 vccd1 vccd1 _10293_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout640 _17506_/Q vssd1 vssd1 vccd1 vccd1 _17065_/A sky130_fd_sc_hd__buf_4
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout651 _12025_/B vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__buf_4
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout662 _17503_/Q vssd1 vssd1 vccd1 vccd1 _09654_/D sky130_fd_sc_hd__buf_6
X_13980_ _13980_/A _13980_/B vssd1 vssd1 vccd1 vccd1 _13982_/B sky130_fd_sc_hd__xnor2_4
XFILLER_93_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout673 fanout676/X vssd1 vssd1 vccd1 vccd1 _13895_/C sky130_fd_sc_hd__buf_4
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout684 fanout686/X vssd1 vssd1 vccd1 vccd1 _16789_/A sky130_fd_sc_hd__buf_8
Xfanout695 _12565_/D vssd1 vssd1 vccd1 vccd1 _12088_/D sky130_fd_sc_hd__buf_6
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12931_ _12931_/A _12931_/B vssd1 vssd1 vccd1 vccd1 _12932_/B sky130_fd_sc_hd__or2_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15651_/A _15651_/B vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__and2_2
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _12386_/X _12389_/X _12862_/S vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__mux2_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14601_/A _14601_/B _14601_/C vssd1 vssd1 vccd1 vccd1 _14603_/A sky130_fd_sc_hd__or3_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _17363_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _14981_/B sky130_fd_sc_hd__and2_1
X_15581_ _15662_/A _15581_/B vssd1 vssd1 vccd1 vccd1 _15582_/B sky130_fd_sc_hd__nand2_4
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12792_/A _12792_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12794_/B sky130_fd_sc_hd__o21a_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14585_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__and2_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _13194_/D _17322_/A2 _17319_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17489_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__nand2b_4
XFILLER_109_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14463_/A _14463_/B _14463_/C vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__nand3_2
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17251_ _17451_/Q _17290_/A2 _17249_/X _17250_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17451_/D sky130_fd_sc_hd__o221a_1
X_11675_ _15056_/A _11675_/B _11675_/C vssd1 vssd1 vccd1 vccd1 _15011_/A sky130_fd_sc_hd__or3_1
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13414_ _13658_/A _17389_/A _13948_/C _13745_/D vssd1 vssd1 vccd1 vccd1 _13415_/B
+ sky130_fd_sc_hd__and4_1
X_16202_ _16098_/A _16101_/Y _16203_/B vssd1 vssd1 vccd1 vccd1 _16292_/B sky130_fd_sc_hd__a21oi_4
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10626_ _10626_/A _10626_/B vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__nor2_2
X_17182_ input29/X wire217/X vssd1 vssd1 vccd1 vccd1 _17198_/C sky130_fd_sc_hd__and2b_1
X_14394_ _14394_/A _14394_/B vssd1 vssd1 vccd1 vccd1 _14396_/B sky130_fd_sc_hd__or2_2
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16133_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16142_/A sky130_fd_sc_hd__xnor2_2
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _13346_/A _13346_/B _13346_/C vssd1 vssd1 vccd1 vccd1 _13347_/A sky130_fd_sc_hd__a21oi_1
XFILLER_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_2
X_16064_ _16064_/A _16064_/B vssd1 vssd1 vccd1 vccd1 _16066_/A sky130_fd_sc_hd__nor2_4
X_13276_ _17371_/A _13276_/B vssd1 vssd1 vccd1 vccd1 _13276_/Y sky130_fd_sc_hd__nor2_1
X_10488_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__nand2b_2
XFILLER_29_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15015_ _16012_/S _16583_/A1 _11854_/X _15013_/Y vssd1 vssd1 vccd1 vccd1 _15015_/X
+ sky130_fd_sc_hd__o31a_1
X_12227_ _12219_/X _12226_/X _14421_/S vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12158_ _12487_/A _12487_/B _12158_/C _12340_/B vssd1 vssd1 vccd1 vccd1 _12325_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11109_ _11075_/A _11075_/B _11075_/C vssd1 vssd1 vccd1 vccd1 _11110_/C sky130_fd_sc_hd__o21ai_4
X_16966_ _16966_/A _16966_/B vssd1 vssd1 vccd1 vccd1 _16969_/A sky130_fd_sc_hd__or2_1
X_12089_ _12089_/A _12089_/B vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__nor2_2
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15917_ _16226_/B _17043_/B vssd1 vssd1 vccd1 vccd1 _15917_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16897_ _16897_/A _16897_/B _16897_/C vssd1 vssd1 vccd1 vccd1 _16900_/A sky130_fd_sc_hd__or3_2
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15848_ _15848_/A _15848_/B vssd1 vssd1 vccd1 vccd1 _15850_/A sky130_fd_sc_hd__nor2_4
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15779_ _15690_/A _15779_/B vssd1 vssd1 vccd1 vccd1 _15781_/B sky130_fd_sc_hd__nand2b_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17518_ fanout927/X _17518_/D vssd1 vssd1 vccd1 vccd1 _17518_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_75_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17449_ fanout938/X _17449_/D vssd1 vssd1 vccd1 vccd1 _17449_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09705_ _09718_/B _09718_/C _09718_/A vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__a21o_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwb_buttons_leds_947 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_947/HI led_enb[0] sky130_fd_sc_hd__conb_1
Xwb_buttons_leds_958 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_958/HI led_enb[11] sky130_fd_sc_hd__conb_1
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09567_ _16933_/A _16982_/B vssd1 vssd1 vccd1 vccd1 _09567_/Y sky130_fd_sc_hd__nor2_2
XFILLER_82_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ _09498_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__or2_2
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _11460_/A _11460_/B _11460_/C vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__or3_4
XFILLER_184_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10427_/A sky130_fd_sc_hd__xnor2_4
XFILLER_165_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ _11630_/A _11391_/B _11436_/B vssd1 vssd1 vccd1 vccd1 _11393_/C sky130_fd_sc_hd__and3_1
XFILLER_164_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13130_ _13127_/X _13128_/Y _12987_/X _12993_/A vssd1 vssd1 vccd1 vccd1 _13130_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ _10342_/A _10342_/B _10342_/C vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__and3_2
XFILLER_192_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _13061_/A _13061_/B _13061_/C vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__nand3_4
XFILLER_151_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10273_ _15707_/A _15622_/A _10272_/X vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__o21a_2
XFILLER_133_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12375_/A sky130_fd_sc_hd__nor2_2
XFILLER_105_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _16750_/A _16750_/B _16883_/C _16670_/C vssd1 vssd1 vccd1 vccd1 _16822_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout470 _12578_/A vssd1 vssd1 vccd1 vccd1 _10904_/B sky130_fd_sc_hd__buf_6
XFILLER_120_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout481 _17521_/Q vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__buf_4
XFILLER_19_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16751_ _16751_/A _16751_/B _16751_/C vssd1 vssd1 vccd1 vccd1 _16753_/A sky130_fd_sc_hd__and3_1
Xfanout492 _17519_/Q vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__clkbuf_16
X_13963_ _13964_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__nand2b_1
XFILLER_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15702_ _15262_/A _16108_/B _15206_/A vssd1 vssd1 vccd1 vccd1 _15705_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12914_ _12915_/A _12915_/B _12915_/C vssd1 vssd1 vccd1 vccd1 _13072_/B sky130_fd_sc_hd__a21oi_2
XFILLER_185_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13894_ _13895_/A _13789_/C _16864_/A vssd1 vssd1 vccd1 vccd1 _13896_/A sky130_fd_sc_hd__a21boi_1
X_16682_ _16680_/X _16682_/B vssd1 vssd1 vccd1 vccd1 _16684_/A sky130_fd_sc_hd__nand2b_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12845_ _12211_/X _12224_/X _12845_/S vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__mux2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15633_ _16304_/A _15623_/X _15632_/X vssd1 vssd1 vccd1 vccd1 _15633_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_185_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _15564_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__xor2_4
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12931_/A _12776_/B vssd1 vssd1 vccd1 vccd1 _12778_/C sky130_fd_sc_hd__or2_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ input61/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17303_/X sky130_fd_sc_hd__or3_1
X_14515_ _14569_/B _14515_/B vssd1 vssd1 vccd1 vccd1 _14518_/C sky130_fd_sc_hd__nand2_1
X_11727_ _11732_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__nand2_2
X_15495_ _15660_/A _15581_/B _15213_/C vssd1 vssd1 vccd1 vccd1 _15496_/B sky130_fd_sc_hd__a21oi_2
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17234_ _17587_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__a21o_1
X_14446_ _14446_/A _14508_/A _14446_/C vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__nand3_4
X_11658_ _14791_/A _15008_/B _11681_/A _11658_/D vssd1 vssd1 vccd1 vccd1 _11678_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10609_ _10610_/B _10610_/A vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__nand2b_2
X_14377_ _14378_/A _14378_/B _14378_/C vssd1 vssd1 vccd1 vccd1 _14446_/A sky130_fd_sc_hd__a21oi_4
XFILLER_128_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17165_ _17165_/A1 _14758_/B _17163_/X _17164_/X vssd1 vssd1 vccd1 vccd1 _17166_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11589_ _11630_/A _11563_/D _11564_/A _11562_/Y vssd1 vssd1 vccd1 vccd1 _11590_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13328_ _13329_/A _13329_/B _13329_/C vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__a21o_1
X_16116_ _15097_/X _15100_/Y _15102_/Y _15123_/Y _15130_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _16116_/X sky130_fd_sc_hd__mux4_1
XFILLER_182_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17096_ _17096_/A _17096_/B _17096_/C vssd1 vssd1 vccd1 vccd1 _17096_/Y sky130_fd_sc_hd__nor3_1
XFILLER_143_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16047_ _16048_/A _16048_/B vssd1 vssd1 vccd1 vccd1 _16047_/X sky130_fd_sc_hd__and2b_1
X_13259_ _13093_/B _13095_/B _13093_/A vssd1 vssd1 vccd1 vccd1 _13260_/A sky130_fd_sc_hd__o21ba_1
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16949_ _16950_/B _16950_/A vssd1 vssd1 vccd1 vccd1 _17003_/B sky130_fd_sc_hd__nand2b_1
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__xnor2_4
X_09352_ _09353_/A _09351_/Y _09928_/C _11813_/B vssd1 vssd1 vccd1 vccd1 _09491_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09283_ _10254_/A _10791_/C vssd1 vssd1 vccd1 vccd1 _17119_/B sky130_fd_sc_hd__nand2_8
XFILLER_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08998_ _17373_/A _11930_/B _12270_/C _12270_/D vssd1 vssd1 vccd1 vccd1 _08999_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_88_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ _10907_/B _10909_/B _10907_/A vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__o21ba_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _09619_/A _09619_/B _09656_/A vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__or3_1
XFILLER_55_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _10891_/A _10891_/B _10891_/C vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__or3_1
XFILLER_188_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12630_ _12631_/A _12631_/B _12631_/C vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__o21a_2
XFILLER_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12561_ _12561_/A _12561_/B _12561_/C vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__or3_1
XFILLER_169_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14300_ _14680_/A _14428_/B vssd1 vssd1 vccd1 vccd1 _14367_/A sky130_fd_sc_hd__nand2_1
X_11512_ _11512_/A _11512_/B _11512_/C vssd1 vssd1 vccd1 vccd1 _11558_/A sky130_fd_sc_hd__nand3_4
XFILLER_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15280_ _15281_/A _15281_/B vssd1 vssd1 vccd1 vccd1 _15428_/A sky130_fd_sc_hd__nor2_4
X_12492_ _12492_/A _12492_/B _12492_/C vssd1 vssd1 vccd1 vccd1 _12494_/A sky130_fd_sc_hd__nor3_1
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14231_ _14154_/A _14156_/B _14154_/B vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__o21ba_1
XFILLER_184_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11443_ _11435_/A _11435_/B _11435_/C vssd1 vssd1 vccd1 vccd1 _11444_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14162_ _14162_/A _14162_/B vssd1 vssd1 vccd1 vccd1 _14237_/B sky130_fd_sc_hd__nor2_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11374_ _11423_/B _15402_/A _11373_/B _11370_/X vssd1 vssd1 vccd1 vccd1 _11376_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13113_ _13114_/A _13114_/B vssd1 vssd1 vccd1 vccd1 _13248_/B sky130_fd_sc_hd__and2_2
X_10325_ _10325_/A _10325_/B vssd1 vssd1 vccd1 vccd1 _10326_/C sky130_fd_sc_hd__and2_2
X_14093_ _14200_/A _14093_/B vssd1 vssd1 vccd1 vccd1 _14094_/C sky130_fd_sc_hd__nor2_1
XFILLER_140_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13181_/B _13044_/B vssd1 vssd1 vccd1 vccd1 _13046_/C sky130_fd_sc_hd__and2_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _10254_/B _10377_/B _10491_/B _10254_/A vssd1 vssd1 vccd1 vccd1 _10257_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_79_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10187_/X sky130_fd_sc_hd__and3_2
XFILLER_182_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16803_ _17140_/A _14864_/B _16798_/Y _16802_/X vssd1 vssd1 vccd1 vccd1 _16803_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_120_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14995_ _14992_/Y _14994_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _14995_/X sky130_fd_sc_hd__mux2_1
XFILLER_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16734_ _13459_/A _17075_/A2 _16733_/X vssd1 vssd1 vccd1 vccd1 _16734_/X sky130_fd_sc_hd__a21o_1
X_13946_ _13948_/B _13948_/C _13948_/D _13948_/A vssd1 vssd1 vccd1 vccd1 _13949_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_75_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16665_ _16665_/A _16665_/B vssd1 vssd1 vccd1 vccd1 _16673_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _14599_/A _14153_/B _14213_/D _14141_/D vssd1 vssd1 vccd1 vccd1 _13878_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_35_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15616_ _15262_/B _16108_/B _15617_/A vssd1 vssd1 vccd1 vccd1 _15616_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_50_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12828_ _12676_/A _12677_/Y _12826_/A _12827_/Y vssd1 vssd1 vccd1 vccd1 _12991_/A
+ sky130_fd_sc_hd__o211a_2
X_16596_ _16748_/C _16596_/B vssd1 vssd1 vccd1 vccd1 _16597_/B sky130_fd_sc_hd__xnor2_2
XFILLER_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15547_ _15530_/A _16008_/C1 _15523_/X _15546_/X vssd1 vssd1 vccd1 vccd1 _15548_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12759_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _12761_/C sky130_fd_sc_hd__xnor2_1
XFILLER_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15478_ _16226_/C _15667_/B _15473_/X _15476_/Y vssd1 vssd1 vccd1 vccd1 _15479_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17217_ _17549_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17217_/X sky130_fd_sc_hd__and2_1
X_14429_ _14430_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _14497_/B sky130_fd_sc_hd__nor2_2
XFILLER_163_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17148_ _17134_/B _16977_/A _17131_/X _17147_/X vssd1 vssd1 vccd1 vccd1 _17573_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__or2_1
X_17079_ _16917_/A _17067_/Y _17068_/X _17078_/X vssd1 vssd1 vccd1 vccd1 _17079_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08921_ _11895_/A _12592_/B _12576_/D _12090_/B vssd1 vssd1 vccd1 vccd1 _08922_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_115_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08852_ _12270_/B _12734_/C _12734_/D _11895_/A vssd1 vssd1 vccd1 vccd1 _08854_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_111_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08783_ _08783_/A _08783_/B _08783_/C vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__or3_2
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _09404_/A _09404_/B vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__xnor2_2
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _09335_/A vssd1 vssd1 vccd1 vccd1 _09335_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09266_ _09407_/B _09509_/B _09791_/B _09838_/A vssd1 vssd1 vccd1 vccd1 _09266_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_193_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _09227_/A _09197_/B vssd1 vssd1 vccd1 vccd1 _09198_/C sky130_fd_sc_hd__and2_1
XFILLER_181_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10110_ _10235_/A _17469_/D _17467_/D _10236_/A vssd1 vssd1 vccd1 vccd1 _10110_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11090_ _11090_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__nor2_2
XFILLER_121_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10041_ _10042_/A _10042_/C vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13800_ _13800_/A _13800_/B _13800_/C vssd1 vssd1 vccd1 vccd1 _13801_/B sky130_fd_sc_hd__and3_1
XFILLER_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11992_ _12155_/A _11991_/B _11971_/X vssd1 vssd1 vccd1 vccd1 _11993_/C sky130_fd_sc_hd__o21ba_2
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14780_ _16317_/A _16014_/A vssd1 vssd1 vccd1 vccd1 _16005_/B sky130_fd_sc_hd__or2_2
XFILLER_95_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13731_ _13936_/A _13732_/B vssd1 vssd1 vccd1 vccd1 _13731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10943_ _10943_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10946_/B sky130_fd_sc_hd__nand3_2
XFILLER_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16450_ _16450_/A _16450_/B vssd1 vssd1 vccd1 vccd1 _16453_/A sky130_fd_sc_hd__xor2_4
XFILLER_44_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13662_ _13662_/A _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__or3_4
X_10874_ _10874_/A _10879_/A _10874_/C vssd1 vssd1 vccd1 vccd1 _10883_/B sky130_fd_sc_hd__or3_4
XFILLER_182_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15401_/A _15402_/B _16533_/A vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__and3_1
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12613_ _12458_/A _12458_/Y _12611_/X _12612_/Y vssd1 vssd1 vccd1 vccd1 _12631_/A
+ sky130_fd_sc_hd__a211oi_4
X_16381_ _16381_/A _16381_/B vssd1 vssd1 vccd1 vccd1 _16385_/A sky130_fd_sc_hd__xor2_4
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _13688_/A _13593_/B vssd1 vssd1 vccd1 vccd1 _13595_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15332_ _15821_/A _16536_/A vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__nand2_2
X_12544_ _11805_/X _11843_/X _12845_/S vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__mux2_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15263_ _15143_/X _15262_/X _15305_/C vssd1 vssd1 vccd1 vccd1 _15263_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_32_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ _12476_/A _12476_/B _12476_/C vssd1 vssd1 vccd1 vccd1 _12477_/A sky130_fd_sc_hd__a21oi_4
XFILLER_184_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17002_ _17003_/A _17003_/B _17003_/C vssd1 vssd1 vccd1 vccd1 _17090_/A sky130_fd_sc_hd__a21o_2
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14214_ _14214_/A _14214_/B vssd1 vssd1 vccd1 vccd1 _14216_/A sky130_fd_sc_hd__nor2_1
XFILLER_184_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11426_ _11426_/A _11426_/B _11426_/C vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__nand3_2
XFILLER_137_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_6 _17558_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _14924_/A _12401_/A _12401_/B _15178_/X _15193_/X vssd1 vssd1 vccd1 vccd1
+ _15194_/X sky130_fd_sc_hd__o311a_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14145_ _14145_/A _14145_/B vssd1 vssd1 vccd1 vccd1 _14146_/B sky130_fd_sc_hd__and2_1
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11357_ _11357_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11359_/B sky130_fd_sc_hd__xor2_2
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ _10542_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10309_/C sky130_fd_sc_hd__and2_2
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ _14077_/A _14077_/B vssd1 vssd1 vccd1 vccd1 _14188_/A sky130_fd_sc_hd__nand2_2
XFILLER_152_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11288_ _11288_/A _11291_/B _11288_/C vssd1 vssd1 vccd1 vccd1 _11351_/A sky130_fd_sc_hd__nand3_4
XFILLER_112_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13027_ _13027_/A _13027_/B vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__nor2_2
X_10239_ _09981_/C _17467_/D _10365_/B _10236_/X vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_39_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ _14978_/A _14978_/B vssd1 vssd1 vccd1 vccd1 _14978_/Y sky130_fd_sc_hd__nor2_1
X_16717_ _16566_/Y _16854_/C _16716_/Y vssd1 vssd1 vccd1 vccd1 _16717_/Y sky130_fd_sc_hd__a21oi_2
X_13929_ _13929_/A _13929_/B vssd1 vssd1 vccd1 vccd1 _13932_/A sky130_fd_sc_hd__xor2_4
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16648_ _17156_/B _16648_/B _16648_/C vssd1 vssd1 vccd1 vccd1 _16648_/X sky130_fd_sc_hd__or3_1
XFILLER_35_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16579_ _17140_/A _16651_/B _16579_/C vssd1 vssd1 vccd1 vccd1 _16579_/X sky130_fd_sc_hd__or3_2
XFILLER_31_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ _09119_/A _09119_/Y _09015_/X _09017_/Y vssd1 vssd1 vccd1 vccd1 _09122_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_31_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09051_ _09051_/A _09051_/B _09051_/C vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__and3_4
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09953_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__xnor2_4
X_08904_ _08904_/A _08904_/B _08904_/C vssd1 vssd1 vccd1 vccd1 _08905_/C sky130_fd_sc_hd__nand3_2
X_09884_ _09884_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09885_/C sky130_fd_sc_hd__xnor2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _12107_/B _12088_/C _12088_/D _12275_/A vssd1 vssd1 vccd1 vccd1 _08835_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__xnor2_4
XFILLER_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _09318_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__nand2_2
XFILLER_178_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10590_ _10694_/B _17468_/D _17467_/D _10694_/A vssd1 vssd1 vccd1 vccd1 _10593_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09249_ _09248_/B _09248_/C _09248_/A vssd1 vssd1 vccd1 vccd1 _09249_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _12261_/A _12261_/B vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__nand2b_1
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11211_ _11719_/B _11211_/B vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__nand2_4
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12191_ _12192_/A _12192_/B vssd1 vssd1 vccd1 vccd1 _12191_/X sky130_fd_sc_hd__and2b_1
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ _11110_/A _11110_/C _11110_/B vssd1 vssd1 vccd1 vccd1 _11143_/D sky130_fd_sc_hd__a21o_2
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput76 _17469_/Q vssd1 vssd1 vccd1 vccd1 leds[3] sky130_fd_sc_hd__clkbuf_2
Xoutput87 _17446_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[12] sky130_fd_sc_hd__clkbuf_2
X_15950_ _15577_/Y _16361_/A _15949_/X vssd1 vssd1 vccd1 vccd1 _15953_/A sky130_fd_sc_hd__o21ai_1
XFILLER_163_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11073_ _11107_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11074_/B sky130_fd_sc_hd__or2_1
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput98 _17456_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14901_ _16807_/A _14901_/B vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__or2_1
X_10024_ _10023_/B _10023_/C _10023_/A vssd1 vssd1 vccd1 vccd1 _10027_/C sky130_fd_sc_hd__a21o_2
XFILLER_62_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15881_ _15881_/A _15881_/B vssd1 vssd1 vccd1 vccd1 _15881_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_76_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14832_ _14832_/A _17153_/A vssd1 vssd1 vccd1 vccd1 _17151_/B sky130_fd_sc_hd__or2_1
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17551_ fanout946/X _17551_/D vssd1 vssd1 vccd1 vccd1 _17551_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14763_ _14758_/Y _14762_/Y _14763_/S vssd1 vssd1 vccd1 vccd1 _17606_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11975_ _08989_/A _08991_/B _08989_/B vssd1 vssd1 vccd1 vccd1 _11982_/A sky130_fd_sc_hd__o21ba_1
XTAP_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16502_ _16595_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__nor2_2
X_13714_ _13814_/B _13713_/B _13713_/C vssd1 vssd1 vccd1 vccd1 _13714_/Y sky130_fd_sc_hd__o21ai_4
X_10926_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10928_/B sky130_fd_sc_hd__xnor2_4
X_17482_ fanout927/X _17482_/D vssd1 vssd1 vccd1 vccd1 _17482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_186_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14694_ _14693_/A _14693_/B _14693_/C vssd1 vssd1 vccd1 vccd1 _14695_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16433_ _16760_/B _16809_/C _16432_/C vssd1 vssd1 vccd1 vccd1 _16434_/B sky130_fd_sc_hd__a21oi_1
X_13645_ _13749_/A _13645_/B _13645_/C vssd1 vssd1 vccd1 vccd1 _13749_/B sky130_fd_sc_hd__nand3_2
XFILLER_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10857_ _10859_/B _10859_/C _10859_/A vssd1 vssd1 vccd1 vccd1 _10857_/Y sky130_fd_sc_hd__a21oi_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16363_/B _16364_/B vssd1 vssd1 vccd1 vccd1 _16365_/B sky130_fd_sc_hd__and2b_1
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13576_ _13576_/A _13576_/B _13576_/C vssd1 vssd1 vccd1 vccd1 _13577_/B sky130_fd_sc_hd__and3_1
X_10788_ _10901_/A _10787_/Y _10899_/C _10897_/B vssd1 vssd1 vccd1 vccd1 _10901_/B
+ sky130_fd_sc_hd__and4bb_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15315_ _16115_/A _15381_/B _15315_/C vssd1 vssd1 vccd1 vccd1 _15315_/X sky130_fd_sc_hd__or3_1
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12527_ _12355_/A _12355_/B _12356_/X vssd1 vssd1 vccd1 vccd1 _12528_/C sky130_fd_sc_hd__o21ba_2
X_16295_ _16295_/A _16295_/B vssd1 vssd1 vccd1 vccd1 _16296_/B sky130_fd_sc_hd__xnor2_1
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15246_ _12858_/Y _15252_/B _15245_/X _15537_/A vssd1 vssd1 vccd1 vccd1 _15246_/X
+ sky130_fd_sc_hd__o22a_1
X_12458_ _12458_/A _12458_/B _12626_/B _12458_/D vssd1 vssd1 vccd1 vccd1 _12458_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_173_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11409_ _11408_/A _11458_/A vssd1 vssd1 vccd1 vccd1 _11411_/B sky130_fd_sc_hd__and2b_2
X_12389_ _12022_/Y _12024_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15177_ _15174_/Y _15175_/X _15176_/Y vssd1 vssd1 vccd1 vccd1 _15177_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_126_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14128_ _12219_/X _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__o21a_1
XFILLER_180_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14059_ _14058_/A _14058_/B _14060_/A vssd1 vssd1 vccd1 vccd1 _14192_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1070 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09103_ _09103_/A _09103_/B vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__xnor2_1
XFILLER_176_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09034_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09048_/C sky130_fd_sc_hd__nand2_1
XFILLER_190_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout800 _12340_/B vssd1 vssd1 vccd1 vccd1 _09555_/C sky130_fd_sc_hd__buf_8
XFILLER_132_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout811 _12502_/B1 vssd1 vssd1 vccd1 vccd1 _12923_/D sky130_fd_sc_hd__buf_12
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__nor2_2
Xfanout822 _12465_/B vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__clkbuf_16
Xfanout833 _11268_/B vssd1 vssd1 vccd1 vccd1 _15381_/A sky130_fd_sc_hd__clkbuf_8
Xfanout844 _14899_/A vssd1 vssd1 vccd1 vccd1 _11518_/C sky130_fd_sc_hd__buf_6
XFILLER_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout855 _10963_/D vssd1 vssd1 vccd1 vccd1 _14906_/B sky130_fd_sc_hd__buf_8
Xfanout866 _17482_/Q vssd1 vssd1 vccd1 vccd1 _17306_/A1 sky130_fd_sc_hd__buf_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__nor2_1
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout877 _17481_/Q vssd1 vssd1 vccd1 vccd1 _11377_/D sky130_fd_sc_hd__clkbuf_16
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout888 _17479_/Q vssd1 vssd1 vccd1 vccd1 _10321_/C sky130_fd_sc_hd__buf_8
Xfanout899 _11553_/D vssd1 vssd1 vccd1 vccd1 _15008_/B sky130_fd_sc_hd__buf_6
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08812_/A _08814_/B _08812_/B vssd1 vssd1 vccd1 vccd1 _08822_/A sky130_fd_sc_hd__o21ba_1
XFILLER_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _11953_/B _09944_/D _09172_/B _09942_/A vssd1 vssd1 vccd1 vccd1 _09798_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08749_ _12237_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__nand2_2
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _16727_/B _16795_/A _16568_/B _16641_/A vssd1 vssd1 vccd1 vccd1 _11760_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_92_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10711_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__xnor2_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _15303_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13430_ _13430_/A _13430_/B vssd1 vssd1 vccd1 vccd1 _13431_/C sky130_fd_sc_hd__and2_2
X_10642_ _10647_/C _10534_/D _10535_/A _10533_/Y vssd1 vssd1 vccd1 vccd1 _10644_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13361_ _13361_/A _13361_/B vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10573_ _10557_/X _10572_/X _10458_/X _10472_/Y vssd1 vssd1 vccd1 vccd1 _10573_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15100_ _15100_/A _15100_/B vssd1 vssd1 vccd1 vccd1 _15100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_181_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12312_/A _12312_/B _12312_/C vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__nand3_2
X_16080_ _16080_/A _16080_/B _16080_/C vssd1 vssd1 vccd1 vccd1 _16081_/B sky130_fd_sc_hd__or3_2
X_13292_ _13292_/A _13292_/B vssd1 vssd1 vccd1 vccd1 _13293_/B sky130_fd_sc_hd__or2_1
XFILLER_181_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12243_ _12243_/A _12243_/B _13094_/B _13088_/B vssd1 vssd1 vccd1 vccd1 _12429_/A
+ sky130_fd_sc_hd__and4_1
X_15031_ _15030_/A _15089_/S _15093_/A _15030_/D vssd1 vssd1 vccd1 vccd1 _15031_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ _12174_/A _12174_/B _12338_/D _12174_/D vssd1 vssd1 vccd1 vccd1 _12175_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_123_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11125_ _11125_/A _11264_/A vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__or2_4
XFILLER_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16982_ _16982_/A _16982_/B _17038_/C vssd1 vssd1 vccd1 vccd1 _17040_/A sky130_fd_sc_hd__or3_2
XFILLER_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15933_ _15933_/A _15933_/B vssd1 vssd1 vccd1 vccd1 _15935_/A sky130_fd_sc_hd__nand2_1
X_11056_ _11157_/B _11055_/B _11055_/C _11055_/D vssd1 vssd1 vccd1 vccd1 _11056_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_95_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10007_ _10007_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _10009_/C sky130_fd_sc_hd__xnor2_2
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15864_ _15864_/A _15864_/B vssd1 vssd1 vccd1 vccd1 _15866_/C sky130_fd_sc_hd__xnor2_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17603_ fanout942/X _17603_/D vssd1 vssd1 vccd1 vccd1 _17603_/Q sky130_fd_sc_hd__dfxtp_1
X_14815_ _16302_/B _16302_/C _16302_/A vssd1 vssd1 vccd1 vccd1 _16398_/A sky130_fd_sc_hd__a21bo_1
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15795_ _16136_/A _15373_/B _15811_/A vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__a21bo_1
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17534_ fanout932/X _17534_/D vssd1 vssd1 vccd1 vccd1 _17534_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14747_/A _14747_/B _14747_/C vssd1 vssd1 vccd1 vccd1 _14748_/A sky130_fd_sc_hd__a21oi_1
X_11958_ _11958_/A _11958_/B _11958_/C vssd1 vssd1 vccd1 vccd1 _11960_/A sky130_fd_sc_hd__or3_1
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17465_ fanout942/X _17465_/D vssd1 vssd1 vccd1 vccd1 _17465_/Q sky130_fd_sc_hd__dfxtp_4
X_10909_ _10909_/A _10909_/B vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__xnor2_4
X_14677_ _14677_/A _14677_/B vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__xnor2_1
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ _12118_/B _11889_/B vssd1 vssd1 vccd1 vccd1 _11891_/C sky130_fd_sc_hd__nand2_2
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16416_ _16595_/A _16667_/A _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16519_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _17164_/A _13628_/B vssd1 vssd1 vccd1 vccd1 _13628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_193_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17396_ input43/X _17396_/A2 _17395_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17526_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ _16347_/A _16347_/B _16345_/X vssd1 vssd1 vccd1 vccd1 _16348_/B sky130_fd_sc_hd__or3b_2
XFILLER_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13559_ _13559_/A vssd1 vssd1 vccd1 vccd1 _13559_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16278_ _16279_/B _16279_/C _16279_/A vssd1 vssd1 vccd1 vccd1 _16280_/A sky130_fd_sc_hd__o21a_1
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15229_ _15230_/A _15230_/B vssd1 vssd1 vccd1 vccd1 _15231_/A sky130_fd_sc_hd__or2_1
XFILLER_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout129 _17270_/A2 vssd1 vssd1 vccd1 vccd1 _17288_/A2 sky130_fd_sc_hd__buf_4
X_09721_ _09721_/A _09721_/B _09739_/B vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__and3_1
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09652_ _09780_/A _09652_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__and3_1
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _09583_/A _09583_/B vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_928 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09017_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09017_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_164_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout630 _14867_/A vssd1 vssd1 vccd1 vccd1 _14318_/C sky130_fd_sc_hd__buf_4
XFILLER_144_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout641 _17506_/Q vssd1 vssd1 vccd1 vccd1 _14593_/C sky130_fd_sc_hd__buf_6
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__or2_1
Xfanout652 _12025_/B vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__buf_4
Xfanout663 _14155_/B vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__buf_8
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout674 fanout676/X vssd1 vssd1 vccd1 vccd1 _16859_/A sky130_fd_sc_hd__clkbuf_16
Xfanout685 fanout686/X vssd1 vssd1 vccd1 vccd1 _13789_/C sky130_fd_sc_hd__buf_4
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12930_ _12931_/A _12931_/B vssd1 vssd1 vccd1 vccd1 _13117_/B sky130_fd_sc_hd__nand2_2
Xfanout696 _12245_/B vssd1 vssd1 vccd1 vccd1 _12565_/D sky130_fd_sc_hd__buf_12
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12383_/X _12385_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__mux2_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14600_/A _14600_/B vssd1 vssd1 vccd1 vccd1 _14601_/C sky130_fd_sc_hd__nor2_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11812_ _14978_/A _14979_/B _14912_/B vssd1 vssd1 vccd1 vccd1 _12546_/C sky130_fd_sc_hd__o21a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _15580_/A _15580_/B vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__nor2_2
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12792_/A _12792_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__nor3_2
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14531_ _14531_/A _14531_/B _14531_/C vssd1 vssd1 vccd1 vccd1 _14532_/B sky130_fd_sc_hd__or3_1
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11732_/A _11732_/C _11732_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__o21bai_4
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17250_ _17560_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17250_/X sky130_fd_sc_hd__and2_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14518_/B _14460_/X _14382_/A _14395_/Y vssd1 vssd1 vccd1 vccd1 _14463_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11674_ _11674_/A _11674_/B vssd1 vssd1 vccd1 vccd1 _15235_/A sky130_fd_sc_hd__or2_2
XFILLER_169_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16201_ _16382_/A _16201_/B vssd1 vssd1 vccd1 vccd1 _16203_/B sky130_fd_sc_hd__or2_4
XFILLER_174_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13413_ _17389_/A _13948_/C _13745_/D _13658_/A vssd1 vssd1 vccd1 vccd1 _13415_/A
+ sky130_fd_sc_hd__a22oi_2
X_10625_ _10970_/A _10743_/C _10528_/A _10526_/Y vssd1 vssd1 vccd1 vccd1 _10626_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_17181_ _17191_/A _17181_/B _17181_/C _17181_/D vssd1 vssd1 vccd1 vccd1 wire217/A
+ sky130_fd_sc_hd__nor4_2
X_14393_ _14393_/A _14393_/B _14393_/C vssd1 vssd1 vccd1 vccd1 _14394_/B sky130_fd_sc_hd__and3_1
XFILLER_155_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _16133_/A _16133_/B vssd1 vssd1 vccd1 vccd1 _16241_/A sky130_fd_sc_hd__and2_1
XFILLER_183_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13344_ _13462_/B _13344_/B vssd1 vssd1 vccd1 vccd1 _13346_/C sky130_fd_sc_hd__nand2_1
X_10556_ _10555_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__and2b_2
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _15955_/Y _16168_/C vssd1 vssd1 vccd1 vccd1 _16064_/B sky130_fd_sc_hd__and2b_1
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__xnor2_4
X_13275_ _12213_/X _12225_/X _13516_/S vssd1 vssd1 vccd1 vccd1 _13276_/B sky130_fd_sc_hd__mux2_1
XFILLER_182_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _14963_/X _14990_/X _15005_/X vssd1 vssd1 vccd1 vccd1 _15014_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12226_ _12222_/X _12225_/X _17369_/A vssd1 vssd1 vccd1 vccd1 _12226_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ _12487_/B _12158_/C _12340_/B _12487_/A vssd1 vssd1 vccd1 vccd1 _12161_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11110_/B sky130_fd_sc_hd__nor2_2
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16965_ _16974_/A _17134_/C _16965_/C vssd1 vssd1 vccd1 vccd1 _16966_/B sky130_fd_sc_hd__and3b_1
X_12088_ _12088_/A _12088_/B _12088_/C _12088_/D vssd1 vssd1 vccd1 vccd1 _12089_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15916_ _16226_/B _15726_/D _15817_/X _16127_/A vssd1 vssd1 vccd1 vccd1 _15916_/X
+ sky130_fd_sc_hd__a22o_1
X_11039_ _11046_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11039_/Y sky130_fd_sc_hd__nand2b_2
X_16896_ _16952_/B _16896_/B vssd1 vssd1 vccd1 vccd1 _16897_/C sky130_fd_sc_hd__and2_1
XFILLER_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15847_ _16056_/A _16355_/B _15846_/B vssd1 vssd1 vccd1 vccd1 _15848_/B sky130_fd_sc_hd__a21oi_2
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _15877_/B _15778_/B vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__or2_1
XFILLER_75_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17517_ fanout936/X _17517_/D vssd1 vssd1 vccd1 vccd1 _17517_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14729_ _14729_/A _14729_/B vssd1 vssd1 vccd1 vccd1 _14731_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ fanout939/X _17448_/D vssd1 vssd1 vccd1 vccd1 _17448_/Q sky130_fd_sc_hd__dfxtp_4
X_17379_ _17379_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17379_/X sky130_fd_sc_hd__or2_1
XFILLER_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09704_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09718_/C sky130_fd_sc_hd__nand2_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwb_buttons_leds_948 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_948/HI led_enb[1] sky130_fd_sc_hd__conb_1
X_09635_ _10321_/A _09803_/B _09517_/A _09515_/Y vssd1 vssd1 vccd1 vccd1 _09636_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xwb_buttons_leds_959 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_959/HI o_wb_stall sky130_fd_sc_hd__conb_1
XFILLER_16_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ _09566_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _16982_/B sky130_fd_sc_hd__nand2_4
XFILLER_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ _09497_/A _09504_/A _09497_/C vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__nor3_1
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _10315_/X _10408_/Y _10402_/Y _10402_/A vssd1 vssd1 vccd1 vccd1 _10410_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _11387_/C _11389_/X _11393_/B vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__o21ba_2
XFILLER_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10341_ _10352_/A _10340_/B _10337_/X vssd1 vssd1 vccd1 vccd1 _10342_/C sky130_fd_sc_hd__a21o_2
XFILLER_180_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13060_ _13060_/A _13060_/B vssd1 vssd1 vccd1 vccd1 _13061_/C sky130_fd_sc_hd__xnor2_4
X_10272_ _14784_/A _15709_/A _15624_/A _10392_/A vssd1 vssd1 vccd1 vccd1 _10272_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _09538_/A _09538_/B _09536_/A vssd1 vssd1 vccd1 vccd1 _12013_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout460 _17523_/Q vssd1 vssd1 vccd1 vccd1 _13298_/A sky130_fd_sc_hd__buf_4
XFILLER_171_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout471 _12578_/A vssd1 vssd1 vccd1 vccd1 _16136_/A sky130_fd_sc_hd__buf_6
X_16750_ _16750_/A _16750_/B vssd1 vssd1 vccd1 vccd1 _16751_/C sky130_fd_sc_hd__xnor2_2
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout482 _11900_/B vssd1 vssd1 vccd1 vccd1 _12107_/B sky130_fd_sc_hd__buf_6
X_13962_ _14047_/A _13962_/B vssd1 vssd1 vccd1 vccd1 _13964_/B sky130_fd_sc_hd__and2_2
Xfanout493 _14785_/A vssd1 vssd1 vccd1 vccd1 _10508_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15701_ _11700_/A _11700_/C _11700_/B vssd1 vssd1 vccd1 vccd1 _15701_/X sky130_fd_sc_hd__a21o_1
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12913_ _12913_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12915_/C sky130_fd_sc_hd__xnor2_1
X_16681_ _16827_/A _16827_/B _16681_/C _16681_/D vssd1 vssd1 vccd1 vccd1 _16682_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13893_ _14383_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _16864_/A sky130_fd_sc_hd__nand2_4
XFILLER_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _16012_/S _16735_/A _13142_/X _15626_/Y _15631_/X vssd1 vssd1 vccd1 vccd1
+ _15632_/X sky130_fd_sc_hd__o311a_1
X_12844_ _12221_/X _12223_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12844_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _15564_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15563_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12775_/A _12775_/B vssd1 vssd1 vccd1 vccd1 _12776_/B sky130_fd_sc_hd__nor2_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _17302_/A1 _17322_/A2 _17301_/X _17428_/B vssd1 vssd1 vccd1 vccd1 _17480_/D
+ sky130_fd_sc_hd__o211a_1
X_14514_ _14514_/A _14514_/B vssd1 vssd1 vccd1 vccd1 _14515_/B sky130_fd_sc_hd__or2_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11727_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15494_ _15494_/A _15846_/B vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__and2_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17233_ _17445_/Q _17233_/A2 _17231_/X _17232_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17445_/D sky130_fd_sc_hd__o221a_1
X_14445_ _14445_/A _14445_/B _14445_/C vssd1 vssd1 vccd1 vccd1 _14446_/C sky130_fd_sc_hd__nand3_2
X_11657_ _11657_/A _11657_/B _11657_/C vssd1 vssd1 vccd1 vccd1 _11658_/D sky130_fd_sc_hd__or3_2
XFILLER_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _10699_/A _10607_/B _10607_/A vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__o21ba_2
XFILLER_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17164_ _17164_/A _17164_/B _17164_/C _17164_/D vssd1 vssd1 vccd1 vccd1 _17164_/X
+ sky130_fd_sc_hd__or4_1
X_14376_ _14376_/A _14376_/B vssd1 vssd1 vccd1 vccd1 _14378_/C sky130_fd_sc_hd__xor2_4
X_11588_ _11579_/A _11579_/C _11579_/B vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__a21o_1
XFILLER_143_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16115_ _16115_/A _16115_/B _16115_/C vssd1 vssd1 vccd1 vccd1 _16122_/A sky130_fd_sc_hd__or3_1
XFILLER_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _13486_/A _13327_/B vssd1 vssd1 vccd1 vccd1 _13329_/C sky130_fd_sc_hd__nor2_2
X_17095_ _17093_/Y _17095_/B vssd1 vssd1 vccd1 vccd1 _17096_/C sky130_fd_sc_hd__and2b_1
X_10539_ _10540_/B _10540_/C _10540_/A vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__a21o_1
XFILLER_155_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16046_ _16046_/A _16046_/B vssd1 vssd1 vccd1 vccd1 _16048_/B sky130_fd_sc_hd__xnor2_2
X_13258_ _13258_/A _13258_/B _13258_/C vssd1 vssd1 vccd1 vccd1 _13261_/B sky130_fd_sc_hd__or3_2
XFILLER_170_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12209_ _12374_/A _12018_/B _12375_/A vssd1 vssd1 vccd1 vccd1 _12210_/B sky130_fd_sc_hd__a21o_2
X_13189_ _13189_/A _13189_/B _13189_/C vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__nand3_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16948_ _16938_/A _09424_/X _16743_/C _16882_/A vssd1 vssd1 vccd1 vccd1 _16950_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_38_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16879_ _16933_/A _15801_/A _17083_/A _16878_/X vssd1 vssd1 vccd1 vccd1 _16880_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09420_ _16983_/A _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__o21ba_4
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _09926_/A _09652_/B _14981_/A vssd1 vssd1 vccd1 vccd1 _09351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _12256_/B _12171_/B vssd1 vssd1 vccd1 vccd1 _16990_/A sky130_fd_sc_hd__nand2_8
XFILLER_127_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08997_ _11930_/B _12270_/C _12270_/D _17373_/A vssd1 vssd1 vccd1 vccd1 _08999_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_29_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09618_ _09618_/A _09618_/B _09747_/A vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__nand3_2
XFILLER_189_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _10891_/B _10891_/C _10891_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__o21ai_2
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _10236_/A _10235_/A _12174_/D _10490_/D vssd1 vssd1 vccd1 vccd1 _09552_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_58_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12560_ _12560_/A _12560_/B vssd1 vssd1 vccd1 vccd1 _12561_/C sky130_fd_sc_hd__xor2_4
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11468_/Y _11471_/X _11469_/X vssd1 vssd1 vccd1 vccd1 _11512_/C sky130_fd_sc_hd__a21o_1
XFILLER_141_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12491_ _12491_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _12492_/C sky130_fd_sc_hd__nor2_1
XFILLER_156_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14230_ _14230_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ _11442_/A _11442_/B vssd1 vssd1 vccd1 vccd1 _11444_/B sky130_fd_sc_hd__xnor2_4
XFILLER_184_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ _14161_/A _14161_/B vssd1 vssd1 vccd1 vccd1 _14237_/A sky130_fd_sc_hd__xor2_4
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11373_ _11370_/X _11373_/B vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__and2b_2
XFILLER_152_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10324_ _10445_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10325_/B sky130_fd_sc_hd__or2_1
X_13112_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13114_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14092_ _14092_/A _14092_/B _14092_/C vssd1 vssd1 vccd1 vccd1 _14093_/B sky130_fd_sc_hd__and3_1
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13043_ _13043_/A _13043_/B _13043_/C vssd1 vssd1 vccd1 vccd1 _13044_/B sky130_fd_sc_hd__or3_1
X_10255_ _10255_/A _10392_/D vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__nand2_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10186_ _10331_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10188_/C sky130_fd_sc_hd__and2_4
XFILLER_182_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16802_ _11849_/Y _14421_/X _16801_/Y vssd1 vssd1 vccd1 vccd1 _16802_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14994_ _15100_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout290 _12865_/S vssd1 vssd1 vccd1 vccd1 _15312_/S sky130_fd_sc_hd__buf_6
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16733_ _16729_/B _17162_/A2 _16733_/B1 _14863_/B _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16733_/X sky130_fd_sc_hd__a221o_1
X_13945_ _15457_/A _13943_/X _13944_/X vssd1 vssd1 vccd1 vccd1 _13945_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16664_ _16935_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16665_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13876_ _13977_/B _14213_/D _14141_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _13878_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15615_ _15615_/A _16207_/B _15615_/C vssd1 vssd1 vccd1 vccd1 _15615_/X sky130_fd_sc_hd__or3_2
XFILLER_179_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12827_ _12825_/A _12825_/B _12825_/C vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__o21ai_4
X_16595_ _16595_/A _16938_/D _16503_/Y vssd1 vssd1 vccd1 vccd1 _16596_/B sky130_fd_sc_hd__or3b_2
XFILLER_15_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15546_ _15309_/B _15533_/Y _15545_/X _15528_/Y vssd1 vssd1 vccd1 vccd1 _15546_/X
+ sky130_fd_sc_hd__o211a_1
X_12758_ _12759_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__nand2b_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11709_ _11465_/A _11464_/B _11708_/A vssd1 vssd1 vccd1 vccd1 _11709_/Y sky130_fd_sc_hd__o21bai_1
X_15477_ _15816_/A _15559_/A _15752_/A _15473_/X vssd1 vssd1 vccd1 vccd1 _15564_/A
+ sky130_fd_sc_hd__or4b_4
X_12689_ _12689_/A _12689_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12691_/A sky130_fd_sc_hd__nor3_2
XFILLER_175_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ _17581_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17216_/X sky130_fd_sc_hd__a21o_1
X_14428_ _14676_/A _14428_/B vssd1 vssd1 vccd1 vccd1 _14430_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ _17167_/B _16485_/A _17137_/X _17146_/X vssd1 vssd1 vccd1 vccd1 _17147_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14359_ _14708_/B _14360_/C _16789_/A _14290_/A vssd1 vssd1 vccd1 vccd1 _14361_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_155_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17078_ _14826_/X _16485_/A _17069_/Y _17077_/X vssd1 vssd1 vccd1 vccd1 _17078_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16029_ _16315_/C _16662_/C _15917_/Y vssd1 vssd1 vccd1 vccd1 _16032_/A sky130_fd_sc_hd__o21a_1
XFILLER_130_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _12592_/B _12576_/D _12567_/B _11895_/A vssd1 vssd1 vccd1 vccd1 _08922_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_112_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08851_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__and2_2
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08782_ _08783_/B _08783_/C _08783_/A vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__o21ai_4
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09403_ _09437_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__nand2_2
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09334_ _09334_/A _09334_/B _09334_/C vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__and3_4
XFILLER_139_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _09838_/A _09407_/B _09509_/B _09791_/B vssd1 vssd1 vccd1 vccd1 _09268_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_193_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09196_ _09196_/A _09196_/B _09202_/A vssd1 vssd1 vccd1 vccd1 _09197_/B sky130_fd_sc_hd__or3_1
XFILLER_193_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10040_ _15711_/A _10431_/B _10034_/A _09900_/Y vssd1 vssd1 vccd1 vccd1 _10042_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11991_ _12155_/A _11991_/B _11971_/X vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__nor3b_4
XFILLER_57_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13730_ _13514_/B _13935_/A _13728_/Y vssd1 vssd1 vccd1 vccd1 _13732_/B sky130_fd_sc_hd__o21ba_1
XFILLER_16_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10942_ _10943_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__a21o_1
XFILLER_45_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ _13770_/A vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__inv_2
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10873_ _10874_/A _10874_/C vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__nor2_2
X_15400_ _15481_/A _15400_/B vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__or2_4
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12612_/A _12612_/B _12612_/C vssd1 vssd1 vccd1 vccd1 _12612_/Y sky130_fd_sc_hd__nor3_4
X_16380_ _16381_/A _16381_/B vssd1 vssd1 vccd1 vccd1 _16563_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13593_/B sky130_fd_sc_hd__and2_1
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _15331_/A _15331_/B vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__xor2_4
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12543_ _11832_/X _11838_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__mux2_1
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15262_ _15262_/A _15262_/B _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _15262_/X
+ sky130_fd_sc_hd__or4_4
X_12474_ _12474_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12476_/C sky130_fd_sc_hd__xnor2_4
XFILLER_185_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17001_ _17052_/B _17001_/B vssd1 vssd1 vccd1 vccd1 _17003_/C sky130_fd_sc_hd__or2_1
X_14213_ _14213_/A _14213_/B _14213_/C _14213_/D vssd1 vssd1 vccd1 vccd1 _14214_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11425_ _11380_/A _11380_/C _11380_/B vssd1 vssd1 vccd1 vccd1 _11426_/C sky130_fd_sc_hd__o21ai_2
X_15193_ _14963_/X _16582_/B _15192_/X _17164_/C _15188_/Y vssd1 vssd1 vccd1 vccd1
+ _15193_/X sky130_fd_sc_hd__o221a_1
XANTENNA_7 _17528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ _14145_/A _14145_/B vssd1 vssd1 vccd1 vccd1 _14229_/B sky130_fd_sc_hd__nor2_2
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ _11357_/A _11357_/B vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__and2b_1
XFILLER_99_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _10307_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__nor2_4
X_14075_ _14165_/A _14075_/B vssd1 vssd1 vccd1 vccd1 _14077_/B sky130_fd_sc_hd__and2_1
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11287_ _11291_/A _11256_/Y _11272_/Y _11311_/A vssd1 vssd1 vccd1 vccd1 _11288_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_106_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13026_ _17397_/A _17395_/A _13897_/B _14153_/C vssd1 vssd1 vccd1 vccd1 _13027_/B
+ sky130_fd_sc_hd__and4_1
X_10238_ _10366_/A _17467_/D vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10169_ _10170_/A _10170_/C vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__nor2_1
XFILLER_120_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14977_ _17131_/A _15028_/A _14977_/C vssd1 vssd1 vccd1 vccd1 _14977_/X sky130_fd_sc_hd__and3_2
XFILLER_35_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16716_ _16558_/B _16560_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__a21oi_4
X_13928_ _13929_/A _13929_/B vssd1 vssd1 vccd1 vccd1 _14030_/B sky130_fd_sc_hd__nand2b_1
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16647_ _16647_/A vssd1 vssd1 vccd1 vccd1 _16648_/C sky130_fd_sc_hd__inv_2
X_13859_ _13961_/B _13859_/B vssd1 vssd1 vccd1 vccd1 _13861_/C sky130_fd_sc_hd__or2_1
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16578_ _16480_/A _16400_/B _16571_/A vssd1 vssd1 vccd1 vccd1 _16579_/C sky130_fd_sc_hd__a21oi_1
X_15529_ _15472_/A _15373_/B _15530_/A vssd1 vssd1 vccd1 vccd1 _15529_/Y sky130_fd_sc_hd__a21boi_1
X_09050_ _09050_/A _09261_/A vssd1 vssd1 vccd1 vccd1 _09051_/C sky130_fd_sc_hd__nand2_2
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__nor2_4
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08903_ _08903_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _08905_/B sky130_fd_sc_hd__xnor2_4
XFILLER_83_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09869_/X _09870_/Y _09877_/X _09881_/X vssd1 vssd1 vccd1 vccd1 _09885_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08800_/X _08801_/Y _08832_/A _08832_/Y vssd1 vssd1 vccd1 vccd1 _08874_/B
+ sky130_fd_sc_hd__a211oi_2
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _11877_/B sky130_fd_sc_hd__nand2b_2
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09317_ _09317_/A _09323_/A _09317_/C vssd1 vssd1 vccd1 vccd1 _09318_/B sky130_fd_sc_hd__or3_1
XFILLER_178_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _09248_/A _09248_/B _09248_/C vssd1 vssd1 vccd1 vccd1 _09248_/Y sky130_fd_sc_hd__nand3_4
XFILLER_193_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09179_ _09179_/A _09179_/B vssd1 vssd1 vccd1 vccd1 _09345_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11210_ _11719_/A _11208_/Y _11168_/A _11168_/Y vssd1 vssd1 vccd1 vccd1 _11211_/B
+ sky130_fd_sc_hd__a211o_1
X_12190_ _12190_/A _12190_/B vssd1 vssd1 vccd1 vccd1 _12192_/B sky130_fd_sc_hd__xnor2_4
XFILLER_123_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _11146_/A _11113_/Y _11128_/Y _11255_/A vssd1 vssd1 vccd1 vccd1 _11143_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput77 _17470_/Q vssd1 vssd1 vccd1 vccd1 leds[4] sky130_fd_sc_hd__clkbuf_2
X_11072_ _11072_/A _11072_/B _11072_/C vssd1 vssd1 vccd1 vccd1 _11075_/B sky130_fd_sc_hd__and3_2
Xoutput88 _17447_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[13] sky130_fd_sc_hd__clkbuf_2
Xoutput99 _17457_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14900_ _15204_/A _16880_/A _15147_/C vssd1 vssd1 vccd1 vccd1 _14900_/X sky130_fd_sc_hd__o21a_1
X_10023_ _10023_/A _10023_/B _10023_/C vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__nand3_1
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15880_ _15881_/A _15881_/B vssd1 vssd1 vccd1 vccd1 _15992_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14831_ _17167_/A _17151_/A _17167_/B vssd1 vssd1 vccd1 vccd1 _14831_/Y sky130_fd_sc_hd__nand3_1
XTAP_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17550_ fanout946/X _17550_/D vssd1 vssd1 vccd1 vccd1 _17550_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14762_ _14762_/A _14762_/B vssd1 vssd1 vccd1 vccd1 _14762_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11974_ _09234_/A _09236_/B _09234_/B vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__o21ba_1
XFILLER_45_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16501_ _16609_/B _16501_/B vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__and2_2
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13713_ _13814_/B _13713_/B _13713_/C vssd1 vssd1 vccd1 vccd1 _13818_/A sky130_fd_sc_hd__or3_4
XTAP_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10925_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _11049_/B sky130_fd_sc_hd__and2_1
X_17481_ fanout927/X _17481_/D vssd1 vssd1 vccd1 vccd1 _17481_/Q sky130_fd_sc_hd__dfxtp_4
X_14693_ _14693_/A _14693_/B _14693_/C vssd1 vssd1 vccd1 vccd1 _14723_/B sky130_fd_sc_hd__and3_1
XFILLER_44_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16432_ _16760_/B _16809_/C _16432_/C vssd1 vssd1 vccd1 vccd1 _16511_/B sky130_fd_sc_hd__and3_1
X_13644_ _13644_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13645_/C sky130_fd_sc_hd__xnor2_2
XFILLER_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ _10865_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10859_/C sky130_fd_sc_hd__nand2_2
XFILLER_147_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16364_/B _16363_/B vssd1 vssd1 vccd1 vccd1 _16365_/A sky130_fd_sc_hd__and2b_2
XFILLER_169_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13576_/A _13576_/B _13576_/C vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__a21oi_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ _11561_/A _10932_/B _10991_/C vssd1 vssd1 vccd1 vccd1 _10787_/Y sky130_fd_sc_hd__a21oi_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15315_/C sky130_fd_sc_hd__nor2_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12526_ _12526_/A _12526_/B _12526_/C vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__and3_2
XFILLER_184_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16294_ _16294_/A _16294_/B vssd1 vssd1 vccd1 vccd1 _16295_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15245_ _14983_/X _14986_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__mux2_1
X_12457_ _12458_/A _12458_/B _12626_/B _12458_/D vssd1 vssd1 vccd1 vccd1 _12457_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_172_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11408_ _11408_/A _11408_/B _11408_/C vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__or3_4
X_15176_ _15119_/A _15119_/B _15117_/A vssd1 vssd1 vccd1 vccd1 _15176_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_193_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12388_ _12384_/X _12387_/X _13838_/S vssd1 vssd1 vccd1 vccd1 _12388_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14127_ _12226_/X _12230_/B _14421_/S vssd1 vssd1 vccd1 vccd1 _14127_/X sky130_fd_sc_hd__mux2_4
XFILLER_153_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11339_ _11340_/B _11340_/A vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__nand2b_4
XFILLER_193_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14058_ _14058_/A _14058_/B vssd1 vssd1 vccd1 vccd1 _14060_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _13010_/B _13268_/A vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ _09103_/B _09103_/A vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__and2b_1
XFILLER_148_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__xnor2_2
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout801 _10839_/D vssd1 vssd1 vccd1 vccd1 _12340_/B sky130_fd_sc_hd__buf_12
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout812 _12502_/B1 vssd1 vssd1 vccd1 vccd1 _10392_/D sky130_fd_sc_hd__buf_8
X_09935_ _10075_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__and2_1
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout823 _14897_/A vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__buf_4
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout834 _11268_/B vssd1 vssd1 vccd1 vccd1 _14896_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout845 _10963_/C vssd1 vssd1 vccd1 vccd1 _14899_/A sky130_fd_sc_hd__clkbuf_8
Xfanout856 _17483_/Q vssd1 vssd1 vccd1 vccd1 _10963_/D sky130_fd_sc_hd__buf_12
XFILLER_131_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09866_ _09866_/A _09866_/B _09884_/B vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__and3_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout867 _17304_/A1 vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__buf_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout878 _10446_/B vssd1 vssd1 vccd1 vccd1 _09944_/D sky130_fd_sc_hd__buf_4
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout889 _17479_/Q vssd1 vssd1 vccd1 vccd1 _17467_/D sky130_fd_sc_hd__buf_6
XFILLER_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08817_ _08831_/B _08831_/C _08831_/A vssd1 vssd1 vccd1 vccd1 _08832_/A sky130_fd_sc_hd__o21a_4
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _09942_/A _09944_/D _10062_/C vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__and3_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _08748_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__and2_2
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__nand2_4
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A _11690_/B vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10641_ _10641_/A _10724_/A vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__nor2_4
XFILLER_42_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13360_ _13360_/A _13360_/B vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__xor2_2
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10572_ _10572_/A _10572_/B _10586_/B vssd1 vssd1 vccd1 vccd1 _10572_/X sky130_fd_sc_hd__or3_4
XFILLER_182_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12311_ _12311_/A _12311_/B vssd1 vssd1 vccd1 vccd1 _12312_/C sky130_fd_sc_hd__xor2_4
XFILLER_127_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13291_ _13292_/A _13292_/B vssd1 vssd1 vccd1 vccd1 _13411_/B sky130_fd_sc_hd__nand2_2
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _15030_/A _15089_/S _15093_/A _15030_/D vssd1 vssd1 vccd1 vccd1 _15093_/B
+ sky130_fd_sc_hd__nand4_2
X_12242_ _12243_/B _13094_/B _13088_/B _12243_/A vssd1 vssd1 vccd1 vccd1 _12244_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_182_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12173_ _12174_/B _12338_/D _12174_/D _12174_/A vssd1 vssd1 vccd1 vccd1 _12175_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_122_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11124_ _11125_/A _11123_/Y _11124_/C _11391_/B vssd1 vssd1 vccd1 vccd1 _11264_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_122_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _16974_/A _17170_/B1 _16980_/X vssd1 vssd1 vccd1 vccd1 _17569_/D sky130_fd_sc_hd__a21oi_1
XFILLER_110_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15932_ _15932_/A _15932_/B _16039_/B _16150_/B vssd1 vssd1 vccd1 vccd1 _15933_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11055_ _11157_/B _11055_/B _11055_/C _11055_/D vssd1 vssd1 vccd1 vccd1 _11055_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10006_ _09991_/Y _10005_/X _09865_/B _09975_/X vssd1 vssd1 vccd1 vccd1 _10028_/A
+ sky130_fd_sc_hd__o211a_1
X_15863_ _15863_/A _15863_/B vssd1 vssd1 vccd1 vccd1 _15864_/B sky130_fd_sc_hd__xnor2_4
XFILLER_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17602_ fanout940/X _17602_/D vssd1 vssd1 vccd1 vccd1 _17602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14814_ _14778_/X _14813_/X _08776_/C vssd1 vssd1 vccd1 vccd1 _16302_/C sky130_fd_sc_hd__a21o_1
XFILLER_188_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15794_ _15794_/A _15794_/B _15888_/B vssd1 vssd1 vccd1 vccd1 _15794_/X sky130_fd_sc_hd__or3b_4
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _14745_/A _14745_/B vssd1 vssd1 vccd1 vccd1 _14747_/C sky130_fd_sc_hd__xnor2_1
X_17533_ fanout932/X _17533_/D vssd1 vssd1 vccd1 vccd1 _17533_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _11957_/A _12163_/B vssd1 vssd1 vccd1 vccd1 _11958_/C sky130_fd_sc_hd__nor2_1
XFILLER_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17464_ fanout938/X _17464_/D vssd1 vssd1 vccd1 vccd1 _17464_/Q sky130_fd_sc_hd__dfxtp_4
X_10908_ _11005_/A _11097_/D vssd1 vssd1 vccd1 vccd1 _10909_/B sky130_fd_sc_hd__nand2_4
X_14676_ _14676_/A _17153_/A vssd1 vssd1 vccd1 vccd1 _14677_/B sky130_fd_sc_hd__nand2_2
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ _11888_/A _11888_/B vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__or2_1
XFILLER_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16415_ _16667_/A _16662_/C _17043_/B _16505_/A vssd1 vssd1 vccd1 vccd1 _16417_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_13627_ _12702_/X _12704_/X _13627_/S vssd1 vssd1 vccd1 vccd1 _13627_/X sky130_fd_sc_hd__mux2_1
X_10839_ _10933_/A _10933_/B _10933_/D _10839_/D vssd1 vssd1 vccd1 vccd1 _10841_/A
+ sky130_fd_sc_hd__and4_2
X_17395_ _17395_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17395_/X sky130_fd_sc_hd__or2_1
XFILLER_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16346_ _16347_/A _16347_/B _16345_/X vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__o21ba_1
XFILLER_186_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ _13558_/A _13558_/B _13558_/C vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__and3_2
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ _12509_/A _12509_/B vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__nor2_4
X_16277_ _16277_/A _16277_/B vssd1 vssd1 vccd1 vccd1 _16283_/A sky130_fd_sc_hd__nand2_4
XFILLER_157_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13489_ _13486_/X _13487_/Y _13365_/Y _13369_/B vssd1 vssd1 vccd1 vccd1 _13490_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15228_ _15228_/A _15228_/B vssd1 vssd1 vccd1 vccd1 _15230_/B sky130_fd_sc_hd__xnor2_1
XFILLER_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15159_ _15159_/A _15159_/B vssd1 vssd1 vccd1 vccd1 _15161_/B sky130_fd_sc_hd__xnor2_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09720_ _09720_/A _09866_/A vssd1 vssd1 vccd1 vccd1 _09739_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09651_ _09779_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09652_/C sky130_fd_sc_hd__and2_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09582_ _11902_/A _10753_/B _09447_/A _09445_/Y vssd1 vssd1 vccd1 vccd1 _09583_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09016_/Y sky130_fd_sc_hd__nand3_4
XFILLER_164_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout620 _14829_/B vssd1 vssd1 vccd1 vccd1 _13300_/C sky130_fd_sc_hd__buf_6
Xfanout631 _08968_/B vssd1 vssd1 vccd1 vccd1 _14867_/A sky130_fd_sc_hd__buf_6
X_09918_ _09912_/B _09912_/C _09912_/A vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__o21bai_4
Xfanout642 _11813_/B vssd1 vssd1 vccd1 vccd1 _12102_/D sky130_fd_sc_hd__buf_6
XFILLER_120_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout653 _17504_/Q vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__buf_6
XFILLER_101_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout664 _14769_/B vssd1 vssd1 vccd1 vccd1 _14865_/B sky130_fd_sc_hd__buf_6
XFILLER_101_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout675 fanout676/X vssd1 vssd1 vccd1 vccd1 _14360_/C sky130_fd_sc_hd__clkbuf_4
Xfanout686 _17501_/Q vssd1 vssd1 vccd1 vccd1 fanout686/X sky130_fd_sc_hd__buf_12
XFILLER_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09849_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09863_/C sky130_fd_sc_hd__nand2_1
Xfanout697 _10311_/D vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__buf_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12860_ _15457_/B _15457_/C _17165_/A1 vssd1 vssd1 vccd1 vccd1 _12860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _17363_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _14979_/B sky130_fd_sc_hd__and2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12791_/A _12947_/B vssd1 vssd1 vccd1 vccd1 _12792_/C sky130_fd_sc_hd__nor2_2
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14531_/A _14531_/B _14531_/C vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__o21ai_2
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A _11742_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__or2_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14382_/A _14395_/Y _14518_/B _14460_/X vssd1 vssd1 vccd1 vccd1 _14463_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_169_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11674_/B sky130_fd_sc_hd__nor2_1
X_16200_ _16200_/A _16200_/B _16200_/C vssd1 vssd1 vccd1 vccd1 _16201_/B sky130_fd_sc_hd__and3_1
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ _13301_/A _13303_/B _13301_/B vssd1 vssd1 vccd1 vccd1 _13420_/A sky130_fd_sc_hd__o21ba_4
XFILLER_169_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17180_ _17180_/A _17180_/B _17180_/C _17180_/D vssd1 vssd1 vccd1 vccd1 _17181_/D
+ sky130_fd_sc_hd__or4_2
X_10624_ _10624_/A _10624_/B vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__xnor2_2
X_14392_ _14394_/A vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__inv_2
XFILLER_155_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16131_ _15913_/A _16023_/Y _16026_/B _16022_/X vssd1 vssd1 vccd1 vccd1 _16133_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_13343_ _17407_/A _16651_/A _13342_/C vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__a21o_1
XFILLER_155_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10555_ _10555_/A _10555_/B _10555_/C vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__or3_4
XFILLER_183_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16062_ _16695_/A _16589_/B _16062_/C vssd1 vssd1 vccd1 vccd1 _16064_/A sky130_fd_sc_hd__and3_2
X_13274_ _15457_/B _13273_/X _17165_/A1 vssd1 vssd1 vccd1 vccd1 _13274_/Y sky130_fd_sc_hd__o21ai_1
X_10486_ _10478_/A _10480_/B _10478_/B vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__o21ba_2
XFILLER_170_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15013_ _11655_/A _15804_/A2 _15007_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _15013_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12225_ _12223_/X _12224_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12156_ _12156_/A _12156_/B vssd1 vssd1 vccd1 vccd1 _12190_/A sky130_fd_sc_hd__nand2_4
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11107_ _11107_/A _11107_/B vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__or2_4
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16964_ _16965_/C _17134_/C _16974_/A vssd1 vssd1 vccd1 vccd1 _16966_/A sky130_fd_sc_hd__a21boi_1
X_12087_ _12256_/B _12088_/C _12088_/D _12088_/A vssd1 vssd1 vccd1 vccd1 _12089_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15915_ _16028_/A _15915_/B vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__or2_2
X_11038_ _11038_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11040_/B sky130_fd_sc_hd__xnor2_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16895_ _16895_/A _16895_/B vssd1 vssd1 vccd1 vccd1 _16896_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15846_ _16056_/A _15846_/B _16355_/B vssd1 vssd1 vccd1 vccd1 _15848_/A sky130_fd_sc_hd__and3_2
XTAP_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ _15877_/A _15776_/B _15776_/C vssd1 vssd1 vccd1 vccd1 _15778_/B sky130_fd_sc_hd__o21a_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12989_ _12819_/X _12824_/A _12987_/X _12988_/Y vssd1 vssd1 vccd1 vccd1 _12993_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17516_ fanout927/X _17516_/D vssd1 vssd1 vccd1 vccd1 _17516_/Q sky130_fd_sc_hd__dfxtp_1
X_14728_ _14726_/X _14728_/B vssd1 vssd1 vccd1 vccd1 _14731_/A sky130_fd_sc_hd__nand2b_1
XFILLER_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14659_ _14698_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14662_/A sky130_fd_sc_hd__and2_4
X_17447_ fanout939/X _17447_/D vssd1 vssd1 vccd1 vccd1 _17447_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17378_ input65/X _17384_/A2 _17377_/Y _17428_/B vssd1 vssd1 vccd1 vccd1 _17517_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16329_ _16329_/A _16425_/B vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__nor2_2
XFILLER_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__xnor2_4
XFILLER_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09645_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwb_buttons_leds_949 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_949/HI led_enb[2] sky130_fd_sc_hd__conb_1
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09565_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__xnor2_4
XFILLER_130_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _09619_/B _09656_/A _09619_/A vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__o21ai_4
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _10337_/X _10340_/B vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__and2b_1
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _14785_/A _10791_/D vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__nand2_2
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12010_ _12010_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__xnor2_2
XFILLER_79_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout450 _11791_/B vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__buf_8
Xfanout461 _11791_/C vssd1 vssd1 vccd1 vccd1 _10254_/B sky130_fd_sc_hd__buf_6
Xfanout472 _17522_/Q vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__buf_12
X_13961_ _13961_/A _13961_/B _13961_/C vssd1 vssd1 vccd1 vccd1 _13962_/B sky130_fd_sc_hd__or3_1
XFILLER_4_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout483 _12595_/B vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__buf_8
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout494 _14785_/A vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__buf_12
XFILLER_46_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12912_ _12913_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__and2_1
X_15700_ _15700_/A _15700_/B vssd1 vssd1 vccd1 vccd1 _15700_/Y sky130_fd_sc_hd__xnor2_2
X_16680_ _16827_/B _16681_/C _16681_/D _16827_/A vssd1 vssd1 vccd1 vccd1 _16680_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13892_ _14013_/A _13892_/B vssd1 vssd1 vccd1 vccd1 _13912_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12843_ _16922_/A _12843_/B vssd1 vssd1 vccd1 vccd1 _12856_/A sky130_fd_sc_hd__nand2_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15631_ _16115_/A _15709_/B _15624_/Y _15628_/X _15630_/X vssd1 vssd1 vccd1 vccd1
+ _15631_/X sky130_fd_sc_hd__o32a_1
XFILLER_104_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15562_ _15655_/A _15655_/B vssd1 vssd1 vccd1 vccd1 _15564_/B sky130_fd_sc_hd__xnor2_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12775_/A _12775_/B vssd1 vssd1 vccd1 vccd1 _12931_/A sky130_fd_sc_hd__and2_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14514_/A _14514_/B vssd1 vssd1 vccd1 vccd1 _14569_/B sky130_fd_sc_hd__nand2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ input58/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17301_/X sky130_fd_sc_hd__or3_1
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11725_/A _11725_/B _11725_/C vssd1 vssd1 vccd1 vccd1 _11731_/B sky130_fd_sc_hd__and3_4
X_15493_ _15948_/A _15687_/B vssd1 vssd1 vccd1 vccd1 _15846_/B sky130_fd_sc_hd__nor2_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14444_ _14445_/A _14445_/B _14445_/C vssd1 vssd1 vccd1 vccd1 _14508_/A sky130_fd_sc_hd__a21o_2
XFILLER_159_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17232_ _17554_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__and2_1
XFILLER_175_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11656_ _11657_/B _11657_/C _11657_/A vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__o21ai_4
XFILLER_174_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _10607_/A _10607_/B vssd1 vssd1 vccd1 vccd1 _10699_/B sky130_fd_sc_hd__nor2_2
X_17163_ _17151_/A _17163_/A2 _17162_/X vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__o21ba_1
X_14375_ _14376_/B _14376_/A vssd1 vssd1 vccd1 vccd1 _14445_/B sky130_fd_sc_hd__nand2b_1
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _11583_/A _11582_/C _11582_/A vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16114_ _16114_/A _16114_/B vssd1 vssd1 vccd1 vccd1 _16115_/C sky130_fd_sc_hd__nor2_1
X_13326_ _13326_/A _13326_/B _13326_/C vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__nor3_1
XFILLER_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17094_ _17093_/A _17093_/B _17093_/C vssd1 vssd1 vccd1 vccd1 _17095_/B sky130_fd_sc_hd__o21ai_1
XFILLER_127_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10538_ _10540_/B _10540_/C _10540_/A vssd1 vssd1 vccd1 vccd1 _10538_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_171_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16045_ _16046_/A _16046_/B vssd1 vssd1 vccd1 vccd1 _16045_/X sky130_fd_sc_hd__and2b_1
XFILLER_143_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _13258_/A _13258_/B _13258_/C vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__o21ai_4
X_10469_ _10469_/A _10469_/B _10469_/C vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__nor3_1
X_12208_ _12375_/B _12208_/B vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__nor2_4
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13188_ _13189_/A _13189_/B _13189_/C vssd1 vssd1 vccd1 vccd1 _13188_/X sky130_fd_sc_hd__and3_2
XFILLER_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12139_ _12305_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__and2_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _16947_/A _16947_/B vssd1 vssd1 vccd1 vccd1 _16950_/A sky130_fd_sc_hd__xnor2_4
XFILLER_65_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16878_ _10254_/B _10013_/B _09711_/X vssd1 vssd1 vccd1 vccd1 _16878_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15829_ _15932_/A _16039_/B _16150_/B _15734_/B vssd1 vssd1 vccd1 vccd1 _15829_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09350_ _09926_/A _09350_/B _14982_/B vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__and3_2
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__xnor2_4
XFILLER_178_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08996_ _08996_/A _08996_/B vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__nor2_4
XFILLER_130_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09617_ _09618_/B _09747_/A _09618_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__a21o_1
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ _09548_/A _09548_/B vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__nor2_2
XFILLER_93_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09479_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09480_/C sky130_fd_sc_hd__xnor2_4
XFILLER_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11553_/B _14792_/B _11509_/B _11506_/X vssd1 vssd1 vccd1 vccd1 _11512_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12490_ _12490_/A _12642_/A _12490_/C vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__nor3_4
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _11442_/B _11442_/A vssd1 vssd1 vccd1 vccd1 _11496_/A sky130_fd_sc_hd__nand2b_1
XFILLER_11_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _14064_/A _14066_/B _14064_/B vssd1 vssd1 vccd1 vccd1 _14161_/B sky130_fd_sc_hd__o21ba_4
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11372_ _11423_/A _11423_/C _11370_/D _15396_/A vssd1 vssd1 vccd1 vccd1 _11373_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__and2b_2
X_10323_ _10445_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__nand2_2
X_14091_ _14092_/A _14092_/B _14092_/C vssd1 vssd1 vccd1 vccd1 _14200_/A sky130_fd_sc_hd__a21oi_2
XFILLER_153_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13042_ _13043_/A _13043_/B _13043_/C vssd1 vssd1 vccd1 vccd1 _13181_/B sky130_fd_sc_hd__o21ai_1
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10254_ _10254_/A _10254_/B _10377_/B _10962_/B vssd1 vssd1 vccd1 vccd1 _10257_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10185_ _10184_/A _10184_/B _10184_/C vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__o21ai_1
XFILLER_67_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16801_ _14925_/Y _15386_/B _16800_/X vssd1 vssd1 vccd1 vccd1 _16801_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14993_ _10321_/C _17302_/A1 _17304_/A1 _17306_/A1 _10430_/A _14982_/A vssd1 vssd1
+ vccd1 vccd1 _14994_/B sky130_fd_sc_hd__mux4_1
Xfanout280 _08723_/Y vssd1 vssd1 vccd1 vccd1 _12054_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout291 _12862_/S vssd1 vssd1 vccd1 vccd1 _12865_/S sky130_fd_sc_hd__buf_6
XFILLER_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16732_ _14863_/B _16652_/B _16731_/Y vssd1 vssd1 vccd1 vccd1 _16732_/X sky130_fd_sc_hd__o21a_1
X_13944_ _11822_/X _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _13944_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16663_ _16661_/X _16663_/B vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__nand2b_1
X_13875_ _13765_/A _13767_/B _13765_/B vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__o21ba_4
XFILLER_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12826_ _12826_/A vssd1 vssd1 vccd1 vccd1 _12826_/Y sky130_fd_sc_hd__clkinv_2
X_15614_ _15614_/A _15614_/B vssd1 vssd1 vccd1 vccd1 _15615_/C sky130_fd_sc_hd__and2_1
X_16594_ _16667_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16748_/C sky130_fd_sc_hd__nor2_2
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15545_ _10419_/A _12401_/A _13012_/X _15536_/X _15544_/X vssd1 vssd1 vccd1 vccd1
+ _15545_/X sky130_fd_sc_hd__o311a_1
X_12757_ _12757_/A _12915_/A vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__and2_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A _11708_/B vssd1 vssd1 vccd1 vccd1 _16105_/A sky130_fd_sc_hd__xor2_4
X_15476_ _15559_/A vssd1 vssd1 vccd1 vccd1 _15476_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ _12499_/B _12501_/B _12499_/A vssd1 vssd1 vccd1 vccd1 _12689_/C sky130_fd_sc_hd__o21ba_2
X_14427_ _14427_/A _14497_/A vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__or2_1
X_17215_ _17439_/Q _17266_/A2 _17213_/X _17214_/X _17372_/C1 vssd1 vssd1 vccd1 vccd1
+ _17439_/D sky130_fd_sc_hd__o221a_1
XFILLER_175_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__xnor2_4
X_17146_ _16917_/A _17135_/Y _17136_/X _17145_/Y vssd1 vssd1 vccd1 vccd1 _17146_/X
+ sky130_fd_sc_hd__a31o_1
X_14358_ _15457_/A _16735_/B _14357_/X vssd1 vssd1 vccd1 vccd1 _14358_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_129_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _13309_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13312_/C sky130_fd_sc_hd__and2_2
X_17077_ _17077_/A _17077_/B _17077_/C _17076_/X vssd1 vssd1 vccd1 vccd1 _17077_/X
+ sky130_fd_sc_hd__or4b_1
X_14289_ _14708_/B _13789_/C _16722_/A _14290_/A vssd1 vssd1 vccd1 vccd1 _14291_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_144_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16028_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16035_/A sky130_fd_sc_hd__xnor2_4
XFILLER_143_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08850_ _08996_/B _08850_/B vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08783_/C sky130_fd_sc_hd__and2b_1
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09402_ _09292_/A _09291_/C _09291_/B vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__a21o_1
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09333_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09334_/C sky130_fd_sc_hd__xnor2_4
XFILLER_179_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _09269_/A _09269_/B vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _09196_/B _09202_/A _09196_/A vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__o21ai_4
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08979_ _12772_/A _11920_/D _08978_/C vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11990_ _11990_/A _11990_/B _11990_/C vssd1 vssd1 vccd1 vccd1 _11991_/B sky130_fd_sc_hd__and3_2
XFILLER_60_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10941_ _10943_/A _10943_/B _10943_/C vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ _13662_/A _13662_/B _13662_/C vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__o21a_2
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10872_ _11124_/C _11334_/C _10854_/A _10852_/Y vssd1 vssd1 vccd1 vccd1 _10874_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_182_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _12612_/A _12612_/B _12612_/C vssd1 vssd1 vccd1 vccd1 _12611_/X sky130_fd_sc_hd__o21a_2
XFILLER_188_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__nor2_2
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15331_/A _15331_/B vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__nor2_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12542_ _12372_/X _12380_/B _12696_/B _12541_/Y _17070_/B vssd1 vssd1 vccd1 vccd1
+ _12542_/Y sky130_fd_sc_hd__a311oi_4
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15261_ _16226_/C _15647_/A vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__nand2_4
X_12473_ _12473_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__xnor2_4
X_14212_ _14213_/B _14213_/C _14213_/D _14213_/A vssd1 vssd1 vccd1 vccd1 _14214_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_172_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17000_ _17000_/A _17000_/B vssd1 vssd1 vccd1 vccd1 _17001_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11424_ _11426_/B vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__clkinv_2
XFILLER_137_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15192_ _15901_/S _15805_/B _15190_/X vssd1 vssd1 vccd1 vccd1 _15192_/X sky130_fd_sc_hd__o21a_1
XANTENNA_8 _17529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14215_/A _14213_/C vssd1 vssd1 vccd1 vccd1 _14145_/B sky130_fd_sc_hd__nand2_1
X_11355_ _11354_/A _11361_/A vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__nand2b_2
XFILLER_152_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10306_ _12398_/S _10309_/B _10183_/A _10181_/Y vssd1 vssd1 vccd1 vccd1 _10307_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14074_ _14074_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _14075_/B sky130_fd_sc_hd__nand2_1
X_11286_ _11272_/Y _11311_/A _11291_/A _11256_/Y vssd1 vssd1 vccd1 vccd1 _11291_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_193_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13025_ _17395_/A _13897_/B _14153_/C _17397_/A vssd1 vssd1 vccd1 vccd1 _13027_/A
+ sky130_fd_sc_hd__a22oi_4
X_10237_ _10236_/B _17468_/D _11027_/D _10236_/A vssd1 vssd1 vccd1 vccd1 _10365_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _15711_/A _10543_/B _10162_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _10170_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10099_ _10094_/A _10092_/X _09806_/A _09807_/Y vssd1 vssd1 vccd1 vccd1 _10348_/B
+ sky130_fd_sc_hd__o211a_2
X_14976_ _15660_/A _15918_/A _15278_/A _15726_/A vssd1 vssd1 vccd1 vccd1 _14977_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16715_ _16853_/A _16853_/B vssd1 vssd1 vccd1 vccd1 _16715_/Y sky130_fd_sc_hd__nand2_2
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ _14254_/A _13903_/B _13803_/A _13801_/A vssd1 vssd1 vccd1 vccd1 _13929_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16646_ _16572_/A _16574_/B _16643_/A _16644_/X vssd1 vssd1 vccd1 vccd1 _16647_/A
+ sky130_fd_sc_hd__a211o_1
X_13858_ _13858_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13859_/B sky130_fd_sc_hd__nor2_1
XFILLER_179_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12812_/A sky130_fd_sc_hd__xnor2_4
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16577_ _16577_/A _16577_/B vssd1 vssd1 vccd1 vccd1 _16577_/X sky130_fd_sc_hd__xor2_1
X_13789_ _13895_/A _13895_/B _13789_/C _14213_/C vssd1 vssd1 vccd1 vccd1 _13790_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15528_ _15525_/X _15526_/X _15527_/Y vssd1 vssd1 vccd1 vccd1 _15528_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15459_ _16011_/A _14919_/X _15806_/B1 vssd1 vssd1 vccd1 vccd1 _15459_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_129_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17129_ _17130_/A _17130_/B vssd1 vssd1 vccd1 vccd1 _17131_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09951_ _09951_/A _09951_/B _09951_/C vssd1 vssd1 vccd1 vccd1 _09952_/B sky130_fd_sc_hd__nor3_2
XFILLER_103_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08902_ _08903_/B _08903_/A vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__nand2b_1
XFILLER_48_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09877_/X _09881_/X _09869_/X _09870_/Y vssd1 vssd1 vccd1 vccd1 _09885_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08832_/A _08832_/Y _08800_/X _08801_/Y vssd1 vssd1 vccd1 vccd1 _08874_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__xor2_4
XFILLER_122_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09316_ _09316_/A _09316_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__and3_2
XFILLER_179_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09247_ _11990_/B _09245_/Y _09152_/Y _09155_/A vssd1 vssd1 vccd1 vccd1 _09248_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09178_/A _09178_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__and3_1
XFILLER_182_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11140_ _11128_/Y _11255_/A _11146_/A _11113_/Y vssd1 vssd1 vccd1 vccd1 _11146_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_190_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput78 _17471_/Q vssd1 vssd1 vccd1 vccd1 leds[5] sky130_fd_sc_hd__clkbuf_2
X_11071_ _11065_/A _11065_/C _11065_/D _11065_/B vssd1 vssd1 vccd1 vccd1 _11071_/Y
+ sky130_fd_sc_hd__a22oi_4
Xoutput89 _17448_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[14] sky130_fd_sc_hd__clkbuf_2
X_10022_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10023_/C sky130_fd_sc_hd__nand2_1
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14830_ _14597_/B _14828_/Y _14829_/X _17167_/A vssd1 vssd1 vccd1 vccd1 _17167_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14761_ _14738_/A _14708_/C _14739_/Y _14748_/A _14760_/Y vssd1 vssd1 vccd1 vccd1
+ _14762_/B sky130_fd_sc_hd__a311o_1
X_11973_ _08993_/C _08992_/Y _08965_/Y vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__a21o_2
XTAP_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16500_ _16747_/A _16499_/B _16499_/C vssd1 vssd1 vccd1 vccd1 _16501_/B sky130_fd_sc_hd__o21ai_1
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13712_ _13605_/A _13605_/B _13562_/A vssd1 vssd1 vccd1 vccd1 _13713_/C sky130_fd_sc_hd__a21oi_2
X_10924_ _10924_/A _10924_/B vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__xnor2_4
XTAP_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14692_ _14723_/A _14692_/B vssd1 vssd1 vccd1 vccd1 _14693_/C sky130_fd_sc_hd__nor2_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17480_ fanout926/X _17480_/D vssd1 vssd1 vccd1 vccd1 _17480_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_186_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _16431_/A _16511_/A vssd1 vssd1 vccd1 vccd1 _16432_/C sky130_fd_sc_hd__nor2_1
XFILLER_16_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13643_ _13643_/A _13948_/C vssd1 vssd1 vccd1 vccd1 _13644_/B sky130_fd_sc_hd__nand2_2
X_10855_ _10855_/A _10855_/B vssd1 vssd1 vccd1 vccd1 _10865_/B sky130_fd_sc_hd__xnor2_4
XFILLER_188_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16362_ _16362_/A _16362_/B vssd1 vssd1 vccd1 vccd1 _16364_/B sky130_fd_sc_hd__xnor2_1
XFILLER_158_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13574_ _13702_/B _13574_/B vssd1 vssd1 vccd1 vccd1 _13576_/C sky130_fd_sc_hd__nand2_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _11561_/A _10932_/B _10991_/C vssd1 vssd1 vccd1 vccd1 _10901_/A sky130_fd_sc_hd__and3_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _12526_/A _12526_/B _12526_/C vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__a21oi_4
X_15313_ _12858_/Y _16011_/C _15312_/X _16011_/A vssd1 vssd1 vccd1 vccd1 _15313_/Y
+ sky130_fd_sc_hd__o22ai_4
X_16293_ _16293_/A _16293_/B vssd1 vssd1 vccd1 vccd1 _16293_/Y sky130_fd_sc_hd__xnor2_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12456_ _12626_/A _12454_/Y _12280_/X _12284_/A vssd1 vssd1 vccd1 vccd1 _12458_/D
+ sky130_fd_sc_hd__a211o_2
X_15244_ _15244_/A _15244_/B _15244_/C vssd1 vssd1 vccd1 vccd1 _15244_/X sky130_fd_sc_hd__or3_1
XFILLER_184_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ _11402_/A _11402_/B _11451_/A vssd1 vssd1 vccd1 vccd1 _11408_/C sky130_fd_sc_hd__o21ba_2
X_15175_ _15175_/A _15175_/B _15796_/B vssd1 vssd1 vccd1 vccd1 _15175_/X sky130_fd_sc_hd__or3_2
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12387_ _12385_/X _12386_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12387_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14126_ _14763_/S _14124_/Y _14205_/B _14038_/Y vssd1 vssd1 vccd1 vccd1 _17593_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _11386_/A _11337_/B _11337_/A vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__o21ba_2
XFILLER_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14057_ _14057_/A _14057_/B vssd1 vssd1 vccd1 vccd1 _14060_/A sky130_fd_sc_hd__xor2_2
XFILLER_113_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11269_ _11122_/B _11518_/C _15244_/A _11320_/A vssd1 vssd1 vccd1 vccd1 _11313_/A
+ sky130_fd_sc_hd__a31o_4
X_13008_ _11781_/B _12377_/Y _13005_/B _13005_/X _13007_/Y vssd1 vssd1 vccd1 vccd1
+ _13010_/B sky130_fd_sc_hd__a311o_4
XFILLER_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14959_ _14958_/A _14956_/Y _14958_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16629_ _16630_/A _16630_/B _16630_/C vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__a21oi_4
XFILLER_165_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09101_ _09101_/A _09165_/A vssd1 vssd1 vccd1 vccd1 _09103_/B sky130_fd_sc_hd__nor2_4
X_09032_ _17081_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__xnor2_2
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout802 _10839_/D vssd1 vssd1 vccd1 vccd1 _13067_/D sky130_fd_sc_hd__buf_6
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _10075_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__nor2_1
XFILLER_132_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout813 _12502_/B1 vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__buf_8
Xfanout824 _14897_/A vssd1 vssd1 vccd1 vccd1 _15450_/A sky130_fd_sc_hd__buf_4
XFILLER_58_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout835 _11268_/B vssd1 vssd1 vccd1 vccd1 _11480_/C sky130_fd_sc_hd__buf_4
Xfanout846 _17484_/Q vssd1 vssd1 vccd1 vccd1 _10963_/C sky130_fd_sc_hd__buf_12
X_09865_ _09865_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__nand2_1
Xfanout857 _17306_/A1 vssd1 vssd1 vccd1 vccd1 _12127_/D sky130_fd_sc_hd__buf_8
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout868 _17304_/A1 vssd1 vssd1 vccd1 vccd1 _11920_/D sky130_fd_sc_hd__buf_6
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout879 _17302_/A1 vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__buf_8
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08831_/C sky130_fd_sc_hd__and2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _11953_/B _10321_/C vssd1 vssd1 vccd1 vccd1 _10062_/C sky130_fd_sc_hd__and2_1
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08747_ _08747_/A vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__inv_2
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _10641_/A _10639_/Y _10640_/C _10640_/D vssd1 vssd1 vccd1 vccd1 _10724_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10586_/B sky130_fd_sc_hd__xnor2_4
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12311_/B sky130_fd_sc_hd__nor2_4
XFILLER_182_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13290_ _13417_/B _13290_/B vssd1 vssd1 vccd1 vccd1 _13292_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12241_ _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12250_/A sky130_fd_sc_hd__xor2_4
XFILLER_163_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12172_ _12172_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__xnor2_1
XFILLER_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11123_ _11122_/B _11480_/C _11518_/C _11266_/A vssd1 vssd1 vccd1 vccd1 _11123_/Y
+ sky130_fd_sc_hd__a22oi_2
X_16980_ _17156_/B _16969_/Y _16979_/X _16963_/X vssd1 vssd1 vccd1 vccd1 _16980_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ _16410_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16040_/A sky130_fd_sc_hd__nor2_1
X_11054_ _11041_/Y _11042_/X _11047_/Y _11050_/X vssd1 vssd1 vccd1 vccd1 _11055_/D
+ sky130_fd_sc_hd__a211o_2
XFILLER_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10005_ _10005_/A _10005_/B _10005_/C vssd1 vssd1 vccd1 vccd1 _10005_/X sky130_fd_sc_hd__and3_4
XFILLER_77_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15862_ _15863_/B _15863_/A vssd1 vssd1 vccd1 vccd1 _15980_/B sky130_fd_sc_hd__and2b_1
XFILLER_92_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17601_ fanout943/X _17601_/D vssd1 vssd1 vccd1 vccd1 _17601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14813_ _16112_/B _16112_/C _16315_/A vssd1 vssd1 vccd1 vccd1 _14813_/X sky130_fd_sc_hd__a21bo_1
XFILLER_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15793_ _15793_/A _15793_/B vssd1 vssd1 vccd1 vccd1 _15794_/B sky130_fd_sc_hd__nor2_1
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17532_ fanout933/X _17532_/D vssd1 vssd1 vccd1 vccd1 _17532_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _14744_/A _14744_/B vssd1 vssd1 vccd1 vccd1 _14745_/B sky130_fd_sc_hd__nand2_1
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _11956_/A _12163_/A _11956_/C vssd1 vssd1 vccd1 vccd1 _12163_/B sky130_fd_sc_hd__nor3_2
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17463_ fanout941/X _17463_/D vssd1 vssd1 vccd1 vccd1 _17463_/Q sky130_fd_sc_hd__dfxtp_4
X_10907_ _10907_/A _10907_/B vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__nor2_2
XFILLER_178_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14675_ _14675_/A _17167_/A vssd1 vssd1 vccd1 vccd1 _14677_/A sky130_fd_sc_hd__xnor2_4
X_11887_ _11888_/A _11888_/B vssd1 vssd1 vccd1 vccd1 _12118_/B sky130_fd_sc_hd__nand2_2
XFILLER_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16414_ _16414_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16422_/A sky130_fd_sc_hd__xor2_2
XFILLER_60_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10838_ _11124_/C _11132_/C vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__nand2_2
X_13626_ _14839_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _13841_/A sky130_fd_sc_hd__nand2_1
X_17394_ input42/X _17396_/A2 _17393_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17525_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _16345_/A _16345_/B vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__or2_1
X_13557_ _13558_/A _13558_/B _13558_/C vssd1 vssd1 vccd1 vccd1 _13557_/Y sky130_fd_sc_hd__a21oi_4
X_10769_ _10769_/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10771_/C sky130_fd_sc_hd__and2_2
XFILLER_121_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _12508_/A _12508_/B _12508_/C vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__nor3_2
XFILLER_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16276_ _16276_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16277_/B sky130_fd_sc_hd__nand2_1
X_13488_ _13365_/Y _13369_/B _13486_/X _13487_/Y vssd1 vssd1 vccd1 vccd1 _13490_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12439_ _12592_/A _12592_/B _17139_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _12616_/A
+ sky130_fd_sc_hd__and4_1
X_15227_ _15166_/A _15166_/B _15162_/A vssd1 vssd1 vccd1 vccd1 _15228_/B sky130_fd_sc_hd__o21a_1
XFILLER_154_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15158_ _15159_/A _15159_/B vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__nand2_2
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14109_ _14013_/A _14013_/B _14013_/C _14110_/B vssd1 vssd1 vccd1 vccd1 _14197_/B
+ sky130_fd_sc_hd__a211o_2
X_15089_ _15774_/A _15088_/Y _15089_/S vssd1 vssd1 vccd1 vccd1 _15091_/B sky130_fd_sc_hd__mux2_1
XFILLER_113_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09650_ _09928_/C _09652_/B _09619_/B _09494_/Y vssd1 vssd1 vccd1 vccd1 _09656_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ _09581_/A _09581_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09581_/Y sky130_fd_sc_hd__nand3_2
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09015_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__and3_2
XFILLER_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout610 _08969_/B vssd1 vssd1 vccd1 vccd1 _13948_/C sky130_fd_sc_hd__buf_4
Xfanout621 _14599_/D vssd1 vssd1 vccd1 vccd1 _14708_/D sky130_fd_sc_hd__buf_4
XFILLER_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout632 _17507_/Q vssd1 vssd1 vccd1 vccd1 _08968_/B sky130_fd_sc_hd__clkbuf_16
X_09917_ _09915_/A _10059_/A _09770_/Y _09830_/X vssd1 vssd1 vccd1 vccd1 _09960_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_99_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout643 _11813_/B vssd1 vssd1 vccd1 vccd1 _12736_/B sky130_fd_sc_hd__buf_4
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout654 _14428_/B vssd1 vssd1 vccd1 vccd1 _13903_/B sky130_fd_sc_hd__clkbuf_16
Xfanout665 _14769_/B vssd1 vssd1 vccd1 vccd1 _14485_/D sky130_fd_sc_hd__buf_6
Xfanout676 _17502_/Q vssd1 vssd1 vccd1 vccd1 fanout676/X sky130_fd_sc_hd__buf_12
X_09848_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__xnor2_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout687 _12565_/C vssd1 vssd1 vccd1 vccd1 _12088_/C sky130_fd_sc_hd__buf_6
XFILLER_101_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout698 _12245_/B vssd1 vssd1 vccd1 vccd1 _10311_/D sky130_fd_sc_hd__buf_4
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09779_/A _09928_/D vssd1 vssd1 vccd1 vccd1 _14952_/A sky130_fd_sc_hd__and2_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11807_/Y _11809_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A _12947_/A _12790_/C vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__nor3_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11741_ _10778_/A _10777_/C _10777_/A vssd1 vssd1 vccd1 vccd1 _11742_/B sky130_fd_sc_hd__o21a_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14518_/A _14459_/B _14459_/C vssd1 vssd1 vccd1 vccd1 _14460_/X sky130_fd_sc_hd__a21o_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11672_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__nand3_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13411_ _13411_/A _13411_/B _13411_/C vssd1 vssd1 vccd1 vccd1 _13423_/B sky130_fd_sc_hd__nand3_4
X_10623_ _10624_/B _10624_/A vssd1 vssd1 vccd1 vccd1 _10623_/X sky130_fd_sc_hd__and2b_2
X_14391_ _14393_/A _14393_/B _14393_/C vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__a21oi_2
X_16130_ _16130_/A _16130_/B vssd1 vssd1 vccd1 vccd1 _16133_/A sky130_fd_sc_hd__xor2_4
X_13342_ _17407_/A _13564_/C _13342_/C vssd1 vssd1 vccd1 vccd1 _13462_/B sky130_fd_sc_hd__nand3_2
XFILLER_183_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10554_ _10406_/B _10474_/Y _10519_/A _10519_/Y vssd1 vssd1 vccd1 vccd1 _10555_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_167_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16061_ _16352_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _16168_/C sky130_fd_sc_hd__nand2_1
X_13273_ _13627_/S _12222_/X _12229_/C _12858_/Y vssd1 vssd1 vccd1 vccd1 _13273_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_143_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10485_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__or2_2
XFILLER_154_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12224_ _11802_/Y _11842_/Y _12546_/B vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__mux2_1
X_15012_ _14796_/C _15899_/A2 _15009_/X _15011_/X _16218_/C1 vssd1 vssd1 vccd1 vccd1
+ _15012_/X sky130_fd_sc_hd__a2111o_1
XFILLER_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12155_ _12155_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _12192_/A sky130_fd_sc_hd__nor2_4
XFILLER_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11106_ _10904_/B _11423_/C _11605_/B _10905_/B vssd1 vssd1 vccd1 vccd1 _11107_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16963_ _16931_/X _16932_/X _16960_/X _16962_/Y vssd1 vssd1 vccd1 vccd1 _16963_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12086_ _11882_/A _11884_/B _11882_/B vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__o21ba_4
XFILLER_96_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15914_ _16315_/B _15658_/Y _16813_/B _15820_/A vssd1 vssd1 vccd1 vccd1 _15915_/B
+ sky130_fd_sc_hd__o22a_1
X_11037_ _11038_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__and2b_4
X_16894_ _16895_/A _16895_/B vssd1 vssd1 vccd1 vccd1 _16952_/B sky130_fd_sc_hd__or2_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _16055_/A _16681_/D vssd1 vssd1 vccd1 vccd1 _16268_/A sky130_fd_sc_hd__or2_1
XTAP_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _15877_/A _15776_/B _15776_/C vssd1 vssd1 vccd1 vccd1 _15877_/B sky130_fd_sc_hd__nor3_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _13125_/B _12986_/Y _12825_/A _12826_/Y vssd1 vssd1 vccd1 vccd1 _12988_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_75_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17515_ fanout927/X _17515_/D vssd1 vssd1 vccd1 vccd1 _17515_/Q sky130_fd_sc_hd__dfxtp_4
X_14727_ _14727_/A _14727_/B vssd1 vssd1 vccd1 vccd1 _14728_/B sky130_fd_sc_hd__or2_1
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__xor2_1
XFILLER_162_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17446_ fanout939/X _17446_/D vssd1 vssd1 vccd1 vccd1 _17446_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_178_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14658_ _14658_/A _14658_/B _14658_/C vssd1 vssd1 vccd1 vccd1 _14659_/B sky130_fd_sc_hd__or3_1
XFILLER_162_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ _13718_/A _13607_/X _13486_/X _13490_/C vssd1 vssd1 vccd1 vccd1 _13609_/X
+ sky130_fd_sc_hd__a211o_2
X_17377_ _17377_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14589_ _13142_/X _13145_/B _17371_/A vssd1 vssd1 vccd1 vccd1 _14590_/B sky130_fd_sc_hd__mux2_2
X_16328_ _16328_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _16425_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16259_ _16352_/A _16352_/B _16259_/C vssd1 vssd1 vccd1 vccd1 _16358_/A sky130_fd_sc_hd__and3_1
XFILLER_173_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09702_ _09702_/A _09706_/B vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__nor2_2
XFILLER_110_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09633_ _10067_/A _09791_/B _09520_/C vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09564_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09581_/A sky130_fd_sc_hd__nand2b_2
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _09619_/B _09494_/Y _09928_/C _09652_/B vssd1 vssd1 vccd1 vccd1 _09656_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_51_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ _14784_/A _15624_/A vssd1 vssd1 vccd1 vccd1 _15622_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout440 _17393_/A vssd1 vssd1 vccd1 vccd1 _13643_/A sky130_fd_sc_hd__buf_6
Xfanout451 _09566_/A vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout462 _10905_/B vssd1 vssd1 vccd1 vccd1 _11006_/B sky130_fd_sc_hd__buf_6
XFILLER_120_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13960_ _13961_/A _13961_/B _13961_/C vssd1 vssd1 vccd1 vccd1 _14047_/A sky130_fd_sc_hd__o21ai_2
Xfanout473 _12107_/A vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__buf_8
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout484 _12595_/B vssd1 vssd1 vccd1 vccd1 _17383_/A sky130_fd_sc_hd__buf_6
Xfanout495 _15472_/A vssd1 vssd1 vccd1 vccd1 _14785_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_101_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _13060_/A _12911_/B vssd1 vssd1 vccd1 vccd1 _12913_/B sky130_fd_sc_hd__and2_1
X_13891_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13892_/B sky130_fd_sc_hd__or2_1
XFILLER_171_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15630_ _15175_/A _15629_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15630_/X sky130_fd_sc_hd__a21o_1
X_12842_ _13003_/B _12842_/B vssd1 vssd1 vccd1 vccd1 _12843_/B sky130_fd_sc_hd__xnor2_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15655_/A _15655_/B vssd1 vssd1 vccd1 vccd1 _15656_/A sky130_fd_sc_hd__nand2_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12775_/B sky130_fd_sc_hd__xnor2_1
XFILLER_187_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _10321_/C _17322_/A2 _17299_/X _17428_/B vssd1 vssd1 vccd1 vccd1 _17479_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A _14512_/B vssd1 vssd1 vccd1 vccd1 _14514_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11217_/A _11215_/Y _11214_/Y vssd1 vssd1 vccd1 vccd1 _11725_/C sky130_fd_sc_hd__o21ai_4
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _15551_/A _15492_/B vssd1 vssd1 vccd1 vccd1 _15687_/B sky130_fd_sc_hd__or2_4
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17586_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__a21o_1
X_14443_ _14443_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14445_/C sky130_fd_sc_hd__xor2_2
X_11655_ _11655_/A _11676_/A vssd1 vssd1 vccd1 vccd1 _11657_/C sky130_fd_sc_hd__and2_1
XFILLER_156_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10606_ _11006_/B _10963_/D _11005_/B _11006_/A vssd1 vssd1 vccd1 vccd1 _10607_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17162_ _17151_/B _17162_/A2 _16974_/B _17153_/A _17170_/B1 vssd1 vssd1 vccd1 vccd1
+ _17162_/X sky130_fd_sc_hd__a221o_1
X_14374_ _14302_/A _14304_/B _14302_/B vssd1 vssd1 vccd1 vccd1 _14376_/B sky130_fd_sc_hd__o21ba_2
X_11586_ _11586_/A _11620_/A _11586_/C vssd1 vssd1 vccd1 vccd1 _11700_/A sky130_fd_sc_hd__nand3_1
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ _16315_/A _16112_/B _16112_/C vssd1 vssd1 vccd1 vccd1 _16113_/Y sky130_fd_sc_hd__a21oi_1
X_13325_ _13326_/A _13326_/B _13326_/C vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__o21a_2
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10537_ _10637_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10540_/C sky130_fd_sc_hd__nand2_2
X_17093_ _17093_/A _17093_/B _17093_/C vssd1 vssd1 vccd1 vccd1 _17093_/Y sky130_fd_sc_hd__nor3_1
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16044_ _16044_/A _16044_/B vssd1 vssd1 vccd1 vccd1 _16046_/B sky130_fd_sc_hd__xor2_4
XFILLER_155_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10468_ _10581_/A _10581_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _11771_/A sky130_fd_sc_hd__o21ai_2
X_13256_ _13256_/A _13256_/B vssd1 vssd1 vccd1 vccd1 _13258_/C sky130_fd_sc_hd__and2_2
X_12207_ _12371_/B _12206_/B _12206_/C vssd1 vssd1 vccd1 vccd1 _12208_/B sky130_fd_sc_hd__o21a_4
X_13187_ _13326_/B _13187_/B vssd1 vssd1 vccd1 vccd1 _13189_/C sky130_fd_sc_hd__nor2_4
X_10399_ _10399_/A _10399_/B vssd1 vssd1 vccd1 vccd1 _10501_/B sky130_fd_sc_hd__nor2_2
XFILLER_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12139_/B sky130_fd_sc_hd__or3_1
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16946_ _16947_/A _16947_/B vssd1 vssd1 vccd1 vccd1 _17003_/A sky130_fd_sc_hd__nand2b_1
X_12069_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12070_/D sky130_fd_sc_hd__inv_2
XFILLER_96_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16877_ _16931_/A _16931_/B _16851_/A vssd1 vssd1 vccd1 vccd1 _16910_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15828_ _15737_/A _15737_/B _15735_/B vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__o21ai_4
XFILLER_18_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15759_ _15759_/A _15759_/B vssd1 vssd1 vccd1 vccd1 _15760_/B sky130_fd_sc_hd__xnor2_4
X_09280_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__nand2b_2
XFILLER_166_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ input70/X _17429_/B _17429_/C vssd1 vssd1 vccd1 vccd1 _17433_/S sky130_fd_sc_hd__or3_4
XFILLER_193_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08995_ _11932_/A _12270_/C _08943_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _09004_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_141_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09616_ _09618_/B _09747_/A _09618_/A vssd1 vssd1 vccd1 vccd1 _09616_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_44_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09547_ _09409_/C _09791_/B _09410_/A _09408_/Y vssd1 vssd1 vccd1 vccd1 _09548_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09478_ _09478_/A _09478_/B _09603_/A vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__nand3_2
XFILLER_180_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11440_ _11440_/A _11479_/A vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__nor2_4
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11371_ _11423_/B _15402_/A vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__nand2_2
XFILLER_165_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10322_ _10322_/A _10322_/B vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__xnor2_2
X_13110_ _13241_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__and2_1
X_14090_ _14090_/A _14090_/B vssd1 vssd1 vccd1 vccd1 _14092_/C sky130_fd_sc_hd__xnor2_2
XFILLER_164_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13041_ _13181_/A _13041_/B vssd1 vssd1 vccd1 vccd1 _13043_/C sky130_fd_sc_hd__and2_1
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__xnor2_4
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10184_ _10184_/A _10184_/B _10184_/C vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__or3_4
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16800_ _14771_/A _14863_/A _17075_/A2 _16799_/X vssd1 vssd1 vccd1 vccd1 _16800_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14992_ _15100_/A _14992_/B vssd1 vssd1 vccd1 vccd1 _14992_/Y sky130_fd_sc_hd__nand2_1
Xfanout270 _16209_/B vssd1 vssd1 vccd1 vccd1 _16644_/B sky130_fd_sc_hd__buf_6
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout281 _08723_/Y vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__buf_8
XFILLER_75_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout292 _12862_/S vssd1 vssd1 vccd1 vccd1 _15130_/S sky130_fd_sc_hd__buf_6
X_16731_ _14863_/B _16652_/B _17140_/A vssd1 vssd1 vccd1 vccd1 _16731_/Y sky130_fd_sc_hd__a21oi_1
X_13943_ _11844_/X _11854_/X _14421_/S vssd1 vssd1 vccd1 vccd1 _13943_/X sky130_fd_sc_hd__mux2_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16662_ _16747_/A _16938_/B _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16663_/B
+ sky130_fd_sc_hd__or4_2
X_13874_ _14018_/A _13874_/B vssd1 vssd1 vccd1 vccd1 _13918_/A sky130_fd_sc_hd__and2_1
XFILLER_90_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15613_ _15610_/Y _15611_/X _15612_/X vssd1 vssd1 vccd1 vccd1 _15613_/Y sky130_fd_sc_hd__a21boi_4
X_12825_ _12825_/A _12825_/B _12825_/C vssd1 vssd1 vccd1 vccd1 _12826_/A sky130_fd_sc_hd__or3_4
X_16593_ _16686_/B _16593_/B vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__nor2_2
XFILLER_188_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15544_ _16115_/A _15624_/B _15541_/Y _15543_/X _15540_/X vssd1 vssd1 vccd1 vccd1
+ _15544_/X sky130_fd_sc_hd__o311a_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12915_/A sky130_fd_sc_hd__o21ai_2
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _15997_/A _15997_/B vssd1 vssd1 vccd1 vccd1 _11707_/Y sky130_fd_sc_hd__nand2_2
XFILLER_175_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15475_ _15475_/A _15918_/A _16246_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _15559_/A
+ sky130_fd_sc_hd__and4_2
X_12687_ _12684_/X _12685_/Y _12528_/A _12530_/A vssd1 vssd1 vccd1 vccd1 _12689_/B
+ sky130_fd_sc_hd__a211oi_4
X_17214_ _17548_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__and2_1
X_14426_ _14593_/A _14593_/B _14769_/B _16859_/A vssd1 vssd1 vccd1 vccd1 _14497_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11638_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__nand2_2
XFILLER_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17145_ _17070_/B _17138_/Y _17144_/X vssd1 vssd1 vccd1 vccd1 _17145_/Y sky130_fd_sc_hd__o21ai_2
X_14357_ _12703_/X _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _14357_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _11557_/X _11603_/A _11526_/B _11552_/X vssd1 vssd1 vccd1 vccd1 _11576_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13308_ _13308_/A _13308_/B _13308_/C vssd1 vssd1 vccd1 vccd1 _13309_/B sky130_fd_sc_hd__nand3_4
XFILLER_170_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17076_ _17164_/A _16582_/A _15180_/X _11849_/Y _14667_/B vssd1 vssd1 vccd1 vccd1
+ _17076_/X sky130_fd_sc_hd__o32a_1
X_14288_ _08718_/A _16653_/B _14287_/X vssd1 vssd1 vccd1 vccd1 _14288_/Y sky130_fd_sc_hd__a21oi_4
X_16027_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16027_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13239_ _13366_/A _13239_/B vssd1 vssd1 vccd1 vccd1 _13241_/B sky130_fd_sc_hd__and2_2
XFILLER_170_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08780_ _08780_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08802_/B sky130_fd_sc_hd__xnor2_2
XFILLER_85_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16929_ _17169_/A1 _16918_/X _16919_/Y _16922_/Y _16928_/X vssd1 vssd1 vccd1 vccd1
+ _16929_/X sky130_fd_sc_hd__o311a_2
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09401_ _09401_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__nor2_4
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _09332_/A _09332_/B _09463_/A vssd1 vssd1 vccd1 vccd1 _09334_/B sky130_fd_sc_hd__nand3_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _09025_/C _09509_/B _09026_/A _09024_/Y vssd1 vssd1 vccd1 vccd1 _09269_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _09196_/B _09194_/B _12488_/A _12338_/D vssd1 vssd1 vccd1 vccd1 _09202_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_159_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08978_ _12772_/A _11920_/D _08978_/C vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__and3_1
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _10940_/A _10940_/B vssd1 vssd1 vccd1 vccd1 _10943_/C sky130_fd_sc_hd__xnor2_4
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10871_ _14801_/A _11100_/B _10870_/A vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__a21oi_4
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12610_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12612_/C sky130_fd_sc_hd__xnor2_4
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13590_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13592_/B sky130_fd_sc_hd__nor2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12541_ _12372_/X _12380_/B _12696_/B vssd1 vssd1 vccd1 vccd1 _12541_/Y sky130_fd_sc_hd__a21oi_2
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15260_ _15238_/A _16008_/C1 _15259_/Y vssd1 vssd1 vccd1 vccd1 _17548_/D sky130_fd_sc_hd__a21oi_1
XFILLER_184_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12472_ _12473_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _12472_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14211_ _14734_/A _14209_/X _14210_/X _14758_/A vssd1 vssd1 vccd1 vccd1 _14211_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_137_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11423_ _11423_/A _11423_/B _11423_/C _11605_/B vssd1 vssd1 vccd1 vccd1 _11426_/B
+ sky130_fd_sc_hd__and4_2
X_15191_ _14916_/X _14959_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15805_/B sky130_fd_sc_hd__mux2_1
XFILLER_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_9 _17532_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _14142_/A _14229_/A vssd1 vssd1 vccd1 vccd1 _14145_/A sky130_fd_sc_hd__or2_1
X_11354_ _11354_/A _11354_/B _11354_/C vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__or3_4
XFILLER_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10305_ _10305_/A _10305_/B _10305_/C vssd1 vssd1 vccd1 vccd1 _10315_/B sky130_fd_sc_hd__nand3_2
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14073_ _14074_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _14165_/A sky130_fd_sc_hd__or2_2
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11285_ _11285_/A _11285_/B _11285_/C vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__and3_4
X_13024_ _13024_/A _13024_/B vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__xor2_4
X_10236_ _10236_/A _10236_/B _17468_/D _11027_/D vssd1 vssd1 vccd1 vccd1 _10236_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_193_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10167_ _10167_/A _10278_/A vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__nor2_2
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14975_ _15081_/A _15820_/A _16025_/A _15415_/A vssd1 vssd1 vccd1 vccd1 _15028_/A
+ sky130_fd_sc_hd__or4_2
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _17138_/A sky130_fd_sc_hd__and2_4
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16714_ _16714_/A _16714_/B vssd1 vssd1 vccd1 vccd1 _16853_/B sky130_fd_sc_hd__or2_1
X_13926_ _14030_/A _13926_/B vssd1 vssd1 vccd1 vccd1 _13929_/A sky130_fd_sc_hd__nand2_4
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16645_ _16643_/A _16644_/X _16572_/A _16574_/B vssd1 vssd1 vccd1 vccd1 _16648_/B
+ sky130_fd_sc_hd__o211a_1
X_13857_ _13858_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13961_/B sky130_fd_sc_hd__and2_1
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12808_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__and2b_1
X_16576_ _12869_/C _16576_/B vssd1 vssd1 vccd1 vccd1 _16577_/B sky130_fd_sc_hd__nand2b_1
X_13788_ _13895_/B _13789_/C _16722_/A _13895_/A vssd1 vssd1 vccd1 vccd1 _13790_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15527_ _15525_/X _15526_/X _15794_/A vssd1 vssd1 vccd1 vccd1 _15527_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_163_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _12739_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__xnor2_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15458_ _15458_/A _15458_/B vssd1 vssd1 vccd1 vccd1 _15458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14409_ _14409_/A _14473_/A _14409_/C vssd1 vssd1 vccd1 vccd1 _14473_/B sky130_fd_sc_hd__nand3_4
XFILLER_117_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15389_ _14790_/A _16583_/A1 _12852_/X _15377_/Y _15388_/X vssd1 vssd1 vccd1 vccd1
+ _15390_/B sky130_fd_sc_hd__o311a_1
XFILLER_128_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17128_ _17128_/A _17128_/B vssd1 vssd1 vccd1 vccd1 _17130_/B sky130_fd_sc_hd__and2_1
XFILLER_7_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17059_ _17037_/B _17009_/B _17014_/B _17014_/C vssd1 vssd1 vccd1 vccd1 _17060_/B
+ sky130_fd_sc_hd__o22ai_4
XFILLER_131_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09950_ _09951_/B _09951_/C _09951_/A vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__o21a_2
X_08901_ _09037_/A _08900_/B _08900_/A vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__o21ba_4
XFILLER_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _10007_/A _10007_/B vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__and2_2
XFILLER_97_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08832_ _08832_/A _08832_/B _08832_/C vssd1 vssd1 vccd1 vccd1 _08832_/Y sky130_fd_sc_hd__nor3_4
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08763_ _11026_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__nand2_4
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ _09316_/A _09316_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__a21oi_4
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _09152_/Y _09155_/A _11990_/B _09245_/Y vssd1 vssd1 vccd1 vccd1 _09248_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09177_ _09357_/A _09364_/A _09357_/C vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__o21a_1
XFILLER_193_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ _11069_/B _11069_/C _11069_/A vssd1 vssd1 vccd1 vccd1 _11070_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput79 _17472_/Q vssd1 vssd1 vccd1 vccd1 leds[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10021_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760_ _14745_/A _14745_/B _14743_/A vssd1 vssd1 vccd1 vccd1 _14760_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11972_ _09240_/A _09240_/B _09239_/A vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__a21o_2
XTAP_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13711_ _13814_/A _13710_/B _13817_/A _13710_/D vssd1 vssd1 vccd1 vccd1 _13713_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_189_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10923_ _10799_/Y _14805_/A _10922_/X vssd1 vssd1 vccd1 vccd1 _10924_/B sky130_fd_sc_hd__o21a_2
XTAP_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14691_ _14691_/A _14691_/B vssd1 vssd1 vccd1 vccd1 _14692_/B sky130_fd_sc_hd__and2_1
XFILLER_71_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16430_ _16604_/B _16589_/B _16758_/B _16814_/B vssd1 vssd1 vccd1 vccd1 _16511_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13642_ _13642_/A _13642_/B vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10854_ _10854_/A _10874_/A vssd1 vssd1 vccd1 vccd1 _10865_/A sky130_fd_sc_hd__or2_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _16361_/A _16361_/B vssd1 vssd1 vccd1 vccd1 _16362_/B sky130_fd_sc_hd__xnor2_4
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13573_ _14248_/A _16789_/A _13572_/C vssd1 vssd1 vccd1 vccd1 _13574_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _11629_/B _10899_/D vssd1 vssd1 vccd1 vccd1 _10991_/C sky130_fd_sc_hd__and2_4
XFILLER_157_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15034_/Y _15037_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15312_/X sky130_fd_sc_hd__mux2_2
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12524_ _12524_/A _12524_/B vssd1 vssd1 vccd1 vccd1 _12526_/C sky130_fd_sc_hd__nand2_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16292_ _16382_/A _16292_/B vssd1 vssd1 vccd1 vccd1 _16293_/B sky130_fd_sc_hd__nor2_2
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ _15244_/A _15244_/B _15244_/C vssd1 vssd1 vccd1 vccd1 _15243_/Y sky130_fd_sc_hd__o21ai_1
X_12455_ _12280_/X _12284_/A _12626_/A _12454_/Y vssd1 vssd1 vccd1 vccd1 _12626_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_172_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11406_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11408_/B sky130_fd_sc_hd__xnor2_4
XFILLER_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15174_ _15175_/A _15796_/B _11377_/C vssd1 vssd1 vccd1 vccd1 _15174_/Y sky130_fd_sc_hd__o21ai_2
X_12386_ _12020_/Y _12055_/Y _15095_/B vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _14278_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14205_/B sky130_fd_sc_hd__or2_1
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11386_/B sky130_fd_sc_hd__nor2_1
XFILLER_153_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14056_ _14057_/A _14057_/B vssd1 vssd1 vccd1 vccd1 _14150_/B sky130_fd_sc_hd__and2b_1
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11268_ _11268_/A _11268_/B _11268_/C _11268_/D vssd1 vssd1 vccd1 vccd1 _11320_/A
+ sky130_fd_sc_hd__and4_2
X_13007_ _12695_/X _13004_/B _13006_/Y vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10219_ _10219_/A _10219_/B _10219_/C vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__or3_4
X_11199_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__and2b_1
XFILLER_95_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14958_ _14958_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _14958_/Y sky130_fd_sc_hd__nor2_1
X_13909_ _14008_/A _13908_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _13910_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14889_ _15305_/C _14924_/A _16012_/S _15025_/B vssd1 vssd1 vccd1 vccd1 _14889_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16628_ _16628_/A _16628_/B vssd1 vssd1 vccd1 vccd1 _16630_/C sky130_fd_sc_hd__xnor2_4
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16559_ _16558_/B _16558_/C _16558_/A vssd1 vssd1 vccd1 vccd1 _16560_/B sky130_fd_sc_hd__a21o_1
XFILLER_149_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09100_ _09101_/A _09099_/Y _12546_/B _12597_/B vssd1 vssd1 vccd1 vccd1 _09165_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_176_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__nor2_1
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__nand2_1
Xfanout803 _10736_/C vssd1 vssd1 vccd1 vccd1 _10970_/B sky130_fd_sc_hd__buf_8
Xfanout814 _15530_/A vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__buf_6
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout825 _14897_/A vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__buf_6
Xfanout836 _17485_/Q vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__buf_6
X_09864_ _09865_/A _09864_/B _09864_/C vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__nand3_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout847 _12127_/C vssd1 vssd1 vccd1 vccd1 _09803_/B sky130_fd_sc_hd__buf_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout858 _17306_/A1 vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__buf_4
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout869 _17481_/Q vssd1 vssd1 vccd1 vccd1 _17304_/A1 sky130_fd_sc_hd__clkbuf_16
XFILLER_86_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08815_ _08815_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__xnor2_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__nor2_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _12068_/A _12068_/B _12068_/D _12637_/D vssd1 vssd1 vccd1 vccd1 _08747_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_100_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__nor2_2
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09229_ _12800_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__nand2_2
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ _12241_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__nand2b_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _12800_/A _12171_/B vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11122_ _11266_/A _11122_/B _11480_/C _14899_/A vssd1 vssd1 vccd1 vccd1 _11125_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15930_ _15209_/Y _16604_/B _16758_/B _16317_/B vssd1 vssd1 vccd1 vccd1 _15933_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11053_ _11055_/C vssd1 vssd1 vccd1 vccd1 _11053_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10004_/A _10004_/B _10004_/C vssd1 vssd1 vccd1 vccd1 _10005_/C sky130_fd_sc_hd__nand3_2
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15861_ _15861_/A _15861_/B vssd1 vssd1 vccd1 vccd1 _15863_/B sky130_fd_sc_hd__xnor2_4
XFILLER_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17600_ fanout941/X _17600_/D vssd1 vssd1 vccd1 vccd1 _17600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14812_ _16005_/B _16005_/C _17119_/B vssd1 vssd1 vccd1 vccd1 _16112_/C sky130_fd_sc_hd__a21bo_1
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15788_/Y _15790_/X _15791_/Y vssd1 vssd1 vccd1 vccd1 _15792_/X sky130_fd_sc_hd__a21o_2
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17531_ fanout933/X _17531_/D vssd1 vssd1 vccd1 vccd1 _17531_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _14743_/A _14743_/B vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__nand2_1
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11955_ _11956_/A _12163_/A _11956_/C vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17462_ fanout941/X _17462_/D vssd1 vssd1 vccd1 vccd1 _17462_/Q sky130_fd_sc_hd__dfxtp_4
X_10906_ _10905_/B _11027_/C _11027_/D _10905_/A vssd1 vssd1 vccd1 vccd1 _10907_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14674_ _14675_/A _17167_/A vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__or2_2
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11886_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11888_/B sky130_fd_sc_hd__xor2_2
XFILLER_60_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16413_ _16414_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16509_/A sky130_fd_sc_hd__nand2_2
X_13625_ _14666_/S _13625_/B vssd1 vssd1 vccd1 vccd1 _13625_/Y sky130_fd_sc_hd__nor2_2
XFILLER_189_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10837_ _10803_/A _10802_/B _10802_/A vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__o21ba_4
X_17393_ _17393_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17393_/X sky130_fd_sc_hd__or2_1
X_16344_ _16344_/A _16344_/B vssd1 vssd1 vccd1 vccd1 _16345_/B sky130_fd_sc_hd__nor2_1
XFILLER_157_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ _13680_/B _13556_/B vssd1 vssd1 vccd1 vccd1 _13558_/C sky130_fd_sc_hd__nor2_2
X_10768_ _10655_/A _10655_/B _10669_/B _10669_/A vssd1 vssd1 vccd1 vccd1 _10769_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _12508_/A _12508_/B _12508_/C vssd1 vssd1 vccd1 vccd1 _12509_/A sky130_fd_sc_hd__o21a_1
X_16275_ _16276_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__or2_2
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _13603_/B _13486_/C _13486_/A vssd1 vssd1 vccd1 vccd1 _13487_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_145_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10699_ _10699_/A _10699_/B vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__xnor2_4
X_15226_ _15226_/A _15226_/B vssd1 vssd1 vccd1 vccd1 _15228_/A sky130_fd_sc_hd__xnor2_2
XFILLER_138_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12438_ _12592_/B _17139_/A _12597_/B _12592_/A vssd1 vssd1 vccd1 vccd1 _12440_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15157_ _15157_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15159_/B sky130_fd_sc_hd__xnor2_4
X_12369_ _12170_/B _12172_/B _12170_/A vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__o21ba_4
XFILLER_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14108_ _14108_/A _14108_/B vssd1 vssd1 vccd1 vccd1 _14110_/B sky130_fd_sc_hd__xor2_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15088_ _15918_/A _15774_/A vssd1 vssd1 vccd1 vccd1 _15088_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _13950_/A _14181_/B _13951_/A _13949_/B vssd1 vssd1 vccd1 vccd1 _14043_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ _09581_/A _09581_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__a21o_4
XFILLER_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09016_/C sky130_fd_sc_hd__xnor2_4
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout600 _15062_/S0 vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__buf_4
Xfanout611 _08969_/B vssd1 vssd1 vccd1 vccd1 _13947_/B sky130_fd_sc_hd__buf_8
Xfanout622 _14829_/B vssd1 vssd1 vccd1 vccd1 _14599_/D sky130_fd_sc_hd__buf_4
X_09916_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__nor2_4
Xfanout633 _12595_/C vssd1 vssd1 vccd1 vccd1 _12270_/D sky130_fd_sc_hd__buf_6
Xfanout644 _17505_/Q vssd1 vssd1 vccd1 vccd1 _11813_/B sky130_fd_sc_hd__clkbuf_16
Xfanout655 _14428_/B vssd1 vssd1 vccd1 vccd1 _13523_/B sky130_fd_sc_hd__buf_4
Xfanout666 _14155_/B vssd1 vssd1 vccd1 vccd1 _14769_/B sky130_fd_sc_hd__buf_6
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__xnor2_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout677 _12567_/B vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__buf_8
XFILLER_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout688 _12021_/B vssd1 vssd1 vccd1 vccd1 _12565_/C sky130_fd_sc_hd__buf_12
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout699 _17499_/Q vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__buf_8
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09778_ _09928_/C _11808_/B _09655_/A _09653_/Y vssd1 vssd1 vccd1 vccd1 _09784_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08729_ input28/X vssd1 vssd1 vccd1 vccd1 _17362_/A sky130_fd_sc_hd__inv_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11737_/Y _11753_/A _11732_/Y _11733_/X vssd1 vssd1 vccd1 vccd1 _11758_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _15524_/C _11671_/B vssd1 vssd1 vccd1 vccd1 _11672_/C sky130_fd_sc_hd__or2_1
XFILLER_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _13411_/A _13411_/B _13411_/C vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__a21o_4
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10622_ _10716_/A _10621_/B _10621_/A vssd1 vssd1 vccd1 vccd1 _10624_/B sky130_fd_sc_hd__o21ba_2
XFILLER_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14390_ _14456_/A _14456_/B vssd1 vssd1 vccd1 vccd1 _14393_/C sky130_fd_sc_hd__xnor2_2
XFILLER_139_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _13341_/A _13462_/A vssd1 vssd1 vccd1 vccd1 _13342_/C sky130_fd_sc_hd__and2_1
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10566_/B _10553_/B vssd1 vssd1 vccd1 vccd1 _10555_/B sky130_fd_sc_hd__nand2_2
XFILLER_182_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16060_ _16060_/A _16060_/B vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__xor2_2
XFILLER_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13272_ _16922_/A _13270_/Y _13386_/B _13143_/Y _13146_/X vssd1 vssd1 vccd1 vccd1
+ _17585_/D sky130_fd_sc_hd__a32o_1
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__xor2_2
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15011_ _15011_/A _15011_/B _15011_/C vssd1 vssd1 vccd1 vccd1 _15011_/X sky130_fd_sc_hd__and3_1
X_12223_ _11837_/Y _11840_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12154_ _12316_/B _12152_/X _11917_/X _11947_/X vssd1 vssd1 vccd1 vccd1 _12193_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_190_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11105_ _11112_/B _11105_/B vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__nand2_4
XFILLER_151_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16962_ _17131_/A _17014_/A vssd1 vssd1 vccd1 vccd1 _16962_/Y sky130_fd_sc_hd__nand2_1
X_12085_ _12085_/A _12085_/B _12085_/C vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__nand3_2
XFILLER_104_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15913_ _15913_/A _16939_/B vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__nor2_4
X_11036_ _11036_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11038_/B sky130_fd_sc_hd__xnor2_4
X_16893_ _16893_/A _16893_/B vssd1 vssd1 vccd1 vccd1 _16895_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15844_ _16758_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16681_/D sky130_fd_sc_hd__nand2_4
XTAP_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15775_ _15775_/A _15775_/B vssd1 vssd1 vccd1 vccd1 _15776_/C sky130_fd_sc_hd__xor2_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12987_ _12825_/A _12826_/Y _13125_/B _12986_/Y vssd1 vssd1 vccd1 vccd1 _12987_/X
+ sky130_fd_sc_hd__o211a_4
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14727_/A _14750_/A _14726_/C vssd1 vssd1 vccd1 vccd1 _14726_/X sky130_fd_sc_hd__and3_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17514_ fanout926/X _17514_/D vssd1 vssd1 vccd1 vccd1 _17514_/Q sky130_fd_sc_hd__dfxtp_1
X_11938_ _09004_/A _09004_/B _09002_/X vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__a21oi_2
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17445_ fanout935/X _17445_/D vssd1 vssd1 vccd1 vccd1 _17445_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14657_ _14658_/A _14658_/B _14658_/C vssd1 vssd1 vccd1 vccd1 _14698_/A sky130_fd_sc_hd__o21ai_2
XFILLER_33_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11869_ _12245_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _11871_/B sky130_fd_sc_hd__nand2_1
X_13608_ _13486_/X _13490_/C _13718_/A _13607_/X vssd1 vssd1 vccd1 vccd1 _13718_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17376_ input64/X _17396_/A2 _17375_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17516_/D
+ sky130_fd_sc_hd__o211a_1
X_14588_ _14763_/S _14586_/X _14587_/Y _14541_/X _14543_/Y vssd1 vssd1 vccd1 vccd1
+ _17600_/D sky130_fd_sc_hd__a32o_1
XFILLER_20_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16327_ _16328_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _16329_/A sky130_fd_sc_hd__and2_1
XFILLER_174_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ _13643_/A _13948_/D _13408_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13541_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_145_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _16174_/A _16174_/B _16175_/B _16175_/A vssd1 vssd1 vccd1 vccd1 _16272_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15209_ _15203_/X _15208_/X _15238_/A vssd1 vssd1 vccd1 vccd1 _15209_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _16189_/A _16189_/B vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__nor2_1
XFILLER_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09701_ _11026_/A _10736_/C _09701_/C vssd1 vssd1 vccd1 vccd1 _09706_/B sky130_fd_sc_hd__and3_2
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _09632_/A _09632_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09563_ _16990_/B _09563_/B vssd1 vssd1 vccd1 vccd1 _09565_/B sky130_fd_sc_hd__xnor2_4
XFILLER_70_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09494_ _09926_/A _09654_/D _14948_/B vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_934 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout430 _11867_/B vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__buf_6
Xfanout441 _12079_/A vssd1 vssd1 vccd1 vccd1 _17393_/A sky130_fd_sc_hd__buf_6
XFILLER_150_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout452 _10905_/A vssd1 vssd1 vccd1 vccd1 _11006_/A sky130_fd_sc_hd__buf_6
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout463 _11791_/C vssd1 vssd1 vccd1 vccd1 _10905_/B sky130_fd_sc_hd__buf_6
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout474 _12595_/A vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__buf_8
XFILLER_86_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout485 _17520_/Q vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__buf_8
XFILLER_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout496 _17519_/Q vssd1 vssd1 vccd1 vccd1 _15472_/A sky130_fd_sc_hd__buf_8
X_12910_ _12910_/A _12910_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _12911_/B sky130_fd_sc_hd__or3_1
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12841_ _13003_/A _12698_/B _12693_/X vssd1 vssd1 vccd1 vccd1 _12842_/B sky130_fd_sc_hd__o21ai_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15558_/Y _15675_/A vssd1 vssd1 vccd1 vccd1 _15655_/B sky130_fd_sc_hd__and2b_4
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12772_/A _13067_/D vssd1 vssd1 vccd1 vccd1 _12773_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14509_/A _14509_/B _14509_/C vssd1 vssd1 vccd1 vccd1 _14512_/B sky130_fd_sc_hd__o21a_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _10766_/C _10766_/B _10764_/X vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__a21bo_2
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15551_/A _15492_/B vssd1 vssd1 vccd1 vccd1 _15581_/B sky130_fd_sc_hd__nor2_8
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17444_/Q _17233_/A2 _17228_/X _17229_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17444_/D sky130_fd_sc_hd__o221a_1
X_14442_ _14367_/A _17023_/A _14370_/A vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__o21ba_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11654_ _14796_/A _11675_/C _11650_/X vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__o21a_1
XFILLER_168_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10605_ _11005_/A _10963_/C vssd1 vssd1 vccd1 vccd1 _10699_/A sky130_fd_sc_hd__nand2_4
X_17161_ _12442_/B _17140_/B _17160_/Y vssd1 vssd1 vccd1 vccd1 _17166_/B sky130_fd_sc_hd__o21ai_1
X_14373_ _14445_/A _14373_/B vssd1 vssd1 vccd1 vccd1 _14376_/A sky130_fd_sc_hd__and2_2
XFILLER_168_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ _11543_/A _11543_/B _11542_/X vssd1 vssd1 vccd1 vccd1 _11586_/C sky130_fd_sc_hd__o21bai_2
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16112_ _16315_/A _16112_/B _16112_/C vssd1 vssd1 vccd1 vccd1 _16112_/X sky130_fd_sc_hd__and3_1
X_13324_ _13324_/A _13324_/B vssd1 vssd1 vccd1 vccd1 _13326_/C sky130_fd_sc_hd__xnor2_1
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17092_ _17118_/A _17092_/B vssd1 vssd1 vccd1 vccd1 _17093_/C sky130_fd_sc_hd__xnor2_1
X_10536_ _10536_/A _10536_/B vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__xnor2_4
XFILLER_182_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16043_ _16043_/A _16043_/B vssd1 vssd1 vccd1 vccd1 _16044_/B sky130_fd_sc_hd__and2_2
XFILLER_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ _13252_/A _13253_/Y _13118_/A _13119_/Y vssd1 vssd1 vccd1 vccd1 _13256_/B
+ sky130_fd_sc_hd__o211ai_1
X_10467_ _10467_/A _10470_/A vssd1 vssd1 vccd1 vccd1 _10581_/C sky130_fd_sc_hd__nor2_1
XFILLER_170_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _12371_/B _12206_/B _12206_/C vssd1 vssd1 vccd1 vccd1 _12375_/B sky130_fd_sc_hd__nor3_4
XFILLER_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _13186_/A _13186_/B vssd1 vssd1 vccd1 vccd1 _13187_/B sky130_fd_sc_hd__and2_1
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _10970_/A _10899_/D _10293_/A _10291_/Y vssd1 vssd1 vccd1 vccd1 _10399_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_123_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12137_ _12138_/A _12138_/B _12138_/C vssd1 vssd1 vccd1 vccd1 _12305_/A sky130_fd_sc_hd__o21ai_4
XFILLER_151_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16945_ _16814_/B _15658_/Y _17119_/C _16883_/C _16887_/A vssd1 vssd1 vccd1 vccd1
+ _16947_/B sky130_fd_sc_hd__a41o_4
X_12068_ _12068_/A _12068_/B _12068_/C _12068_/D vssd1 vssd1 vccd1 vccd1 _12239_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11019_ _11020_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__and2_2
X_16876_ _16859_/A _16806_/A2 _16857_/Y _16875_/X vssd1 vssd1 vccd1 vccd1 _17567_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15827_ _15827_/A _15827_/B vssd1 vssd1 vccd1 vccd1 _15837_/A sky130_fd_sc_hd__xor2_4
XTAP_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758_ _15759_/A _15759_/B vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__or2_2
XFILLER_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14709_ _14677_/A _14677_/B _14674_/X vssd1 vssd1 vccd1 vccd1 _14744_/A sky130_fd_sc_hd__o21ai_4
X_15689_ _15782_/B _15689_/B vssd1 vssd1 vccd1 vccd1 _15690_/C sky130_fd_sc_hd__nand2_2
XFILLER_33_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17428_ input68/X _17428_/B _17428_/C _17428_/D vssd1 vssd1 vccd1 vccd1 _17542_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_178_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17359_ input60/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17359_/X sky130_fd_sc_hd__or3_1
XFILLER_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08994_ _08994_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09615_ _09746_/A _09754_/A _09746_/C vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__o21ai_4
XFILLER_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09546_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__xor2_2
XFILLER_36_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09477_ _09478_/B _09603_/A _09478_/A vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__a21o_1
XFILLER_145_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11370_ _15396_/A _11423_/A _11370_/C _11370_/D vssd1 vssd1 vccd1 vccd1 _11370_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_180_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10321_ _10321_/A _10560_/A _10321_/C _10560_/D vssd1 vssd1 vccd1 vccd1 _10445_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_30_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _13040_/A _13040_/B _13040_/C vssd1 vssd1 vccd1 vccd1 _13041_/B sky130_fd_sc_hd__or3_1
XFILLER_140_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10252_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__nand2b_2
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10183_ _10183_/A _10307_/A vssd1 vssd1 vccd1 vccd1 _10184_/C sky130_fd_sc_hd__nor2_1
XFILLER_65_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14991_ _12295_/D _12463_/D _12618_/D _12770_/D _10430_/A _14982_/A vssd1 vssd1 vccd1
+ vccd1 _14992_/B sky130_fd_sc_hd__mux4_1
Xfanout260 _17295_/X vssd1 vssd1 vccd1 vccd1 _17355_/C sky130_fd_sc_hd__buf_2
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout271 _14939_/X vssd1 vssd1 vccd1 vccd1 _16209_/B sky130_fd_sc_hd__buf_4
XFILLER_8_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout282 _15096_/S vssd1 vssd1 vccd1 vccd1 _17365_/A sky130_fd_sc_hd__clkbuf_8
X_13942_ _17070_/B _13940_/X _14032_/B _13842_/X vssd1 vssd1 vccd1 vccd1 _17591_/D
+ sky130_fd_sc_hd__o31ai_1
XFILLER_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16730_ _16730_/A _16730_/B vssd1 vssd1 vccd1 vccd1 _16730_/Y sky130_fd_sc_hd__xnor2_1
Xfanout293 _12862_/S vssd1 vssd1 vccd1 vccd1 _15035_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16661_ _16938_/B _16662_/C _16662_/D _16747_/A vssd1 vssd1 vccd1 vccd1 _16661_/X
+ sky130_fd_sc_hd__o22a_1
X_13873_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _13874_/B sky130_fd_sc_hd__or2_1
XFILLER_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15612_ _15610_/Y _15611_/X _16911_/A vssd1 vssd1 vccd1 vccd1 _15612_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12824_ _12824_/A _12824_/B vssd1 vssd1 vccd1 vccd1 _12825_/C sky130_fd_sc_hd__nand2_2
X_16592_ _16814_/B _16935_/B _16591_/C vssd1 vssd1 vccd1 vccd1 _16593_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15543_ _10716_/A _17163_/A2 _15542_/X vssd1 vssd1 vccd1 vccd1 _15543_/X sky130_fd_sc_hd__o21ba_1
XFILLER_187_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12755_ _12755_/A _12755_/B _12755_/C vssd1 vssd1 vccd1 vccd1 _12757_/A sky130_fd_sc_hd__or3_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _15793_/A _15793_/B _15889_/A _11705_/Y _11704_/B vssd1 vssd1 vccd1 vccd1
+ _15997_/B sky130_fd_sc_hd__a32o_4
X_15474_ _14899_/X _14968_/X _16827_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15645_/B
+ sky130_fd_sc_hd__a211o_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12528_/A _12530_/A _12684_/X _12685_/Y vssd1 vssd1 vccd1 vccd1 _12689_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_175_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14425_ _14593_/B _14769_/B _16859_/A _14593_/A vssd1 vssd1 vccd1 vccd1 _14427_/A
+ sky130_fd_sc_hd__a22oi_1
X_17213_ _17580_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17213_/X sky130_fd_sc_hd__a21o_1
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__nor2_2
XFILLER_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17144_ _16582_/A _16011_/X _17140_/X _17143_/X vssd1 vssd1 vccd1 vccd1 _17144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14356_ _12706_/X _12710_/B _14356_/S vssd1 vssd1 vccd1 vccd1 _16735_/B sky130_fd_sc_hd__mux2_4
XFILLER_156_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11568_ _11568_/A _11568_/B _11568_/C vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__and3_2
XFILLER_183_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13307_ _13308_/A _13308_/B _13308_/C vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__a21o_1
XFILLER_171_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ _10519_/A _10519_/B _10519_/C vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__nor3_4
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17075_ _14434_/Y _17075_/A2 _17074_/X vssd1 vssd1 vccd1 vccd1 _17077_/C sky130_fd_sc_hd__a21o_1
XFILLER_128_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14287_ _12549_/X _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _14287_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11499_ _11499_/A _11499_/B _11499_/C vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__nor3_4
XFILLER_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16026_ _16026_/A _16026_/B vssd1 vssd1 vccd1 vccd1 _16028_/B sky130_fd_sc_hd__xnor2_4
X_13238_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13239_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _17391_/A _13298_/A _13300_/D _13169_/D vssd1 vssd1 vccd1 vccd1 _13170_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_151_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16928_ _14667_/A _14543_/B _16924_/Y _16927_/X vssd1 vssd1 vccd1 vccd1 _16928_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16859_ _16859_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _16859_/Y sky130_fd_sc_hd__nor2_2
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09400_ _09311_/A _09316_/B _09311_/C vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__a21oi_2
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _09332_/B _09463_/A _09332_/A vssd1 vssd1 vccd1 vccd1 _09334_/A sky130_fd_sc_hd__a21o_4
XFILLER_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__xnor2_1
XFILLER_166_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ _09194_/B vssd1 vssd1 vccd1 vccd1 _09193_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08977_ _08977_/A _09238_/A vssd1 vssd1 vccd1 vccd1 _08978_/C sky130_fd_sc_hd__nor2_1
XFILLER_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10870_ _10870_/A _10870_/B vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__nor2_4
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09391_/C _09399_/Y _09458_/X _09628_/A vssd1 vssd1 vccd1 vccd1 _09530_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__xnor2_4
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _17373_/A _12592_/C _12471_/C vssd1 vssd1 vccd1 vccd1 _12473_/B sky130_fd_sc_hd__and3_4
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14210_ _14210_/A _14210_/B vssd1 vssd1 vccd1 vccd1 _14210_/X sky130_fd_sc_hd__or2_1
XFILLER_184_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11422_ _11395_/B _11383_/C _11383_/B vssd1 vssd1 vccd1 vccd1 _11435_/B sky130_fd_sc_hd__a21o_1
X_15190_ _15254_/S _14918_/Y _15189_/Y _15711_/A vssd1 vssd1 vccd1 vccd1 _15190_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14141_ _14290_/A _14213_/B _14213_/D _14141_/D vssd1 vssd1 vccd1 vccd1 _14229_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_165_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11353_ _11351_/A _11351_/C _11402_/A vssd1 vssd1 vccd1 vccd1 _11354_/C sky130_fd_sc_hd__a21oi_2
XFILLER_180_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _10305_/B _10305_/C _10305_/A vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__a21o_1
X_14072_ _14072_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11284_ _11352_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11285_/C sky130_fd_sc_hd__and2_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13023_ _13024_/A _13024_/B vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__nand2_2
X_10235_ _10235_/A _11027_/D vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__nand2_8
XFILLER_133_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10166_ _10167_/A _10165_/Y _14788_/A _10534_/D vssd1 vssd1 vccd1 vccd1 _10278_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10097_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__nand2_2
X_14974_ _15278_/A vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__inv_2
X_16713_ _16714_/A _16714_/B vssd1 vssd1 vccd1 vccd1 _16853_/A sky130_fd_sc_hd__nand2_2
X_13925_ _13925_/A _13925_/B _13925_/C vssd1 vssd1 vccd1 vccd1 _13926_/B sky130_fd_sc_hd__nand3_2
XFILLER_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13856_ _13856_/A _13856_/B vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__xnor2_1
X_16644_ _16651_/A _16644_/B _16644_/C vssd1 vssd1 vccd1 vccd1 _16644_/X sky130_fd_sc_hd__and3b_1
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ _12807_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13787_ _13787_/A _13787_/B vssd1 vssd1 vccd1 vccd1 _13805_/A sky130_fd_sc_hd__xnor2_1
X_16575_ _16481_/A _16482_/Y _16572_/Y _16574_/Y vssd1 vssd1 vccd1 vccd1 _16575_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10999_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__and3_4
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _15524_/B _11671_/B _15447_/A vssd1 vssd1 vccd1 vccd1 _15526_/X sky130_fd_sc_hd__a21o_1
X_12738_ _12739_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12903_/A sky130_fd_sc_hd__and2b_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15457_ _15457_/A _15457_/B _15457_/C vssd1 vssd1 vccd1 vccd1 _15467_/C sky130_fd_sc_hd__or3_2
XFILLER_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ _12816_/A _12669_/B vssd1 vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__and2_2
X_14408_ _14424_/B _14406_/Y _14340_/B _14342_/A vssd1 vssd1 vccd1 vccd1 _14409_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_175_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15388_ _17164_/C _15380_/X _15387_/X _15379_/X vssd1 vssd1 vccd1 vccd1 _15388_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14339_ _14336_/X _14337_/Y _14222_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14340_/C
+ sky130_fd_sc_hd__o211ai_4
X_17127_ _17127_/A _17127_/B vssd1 vssd1 vccd1 vccd1 _17128_/B sky130_fd_sc_hd__nand2_1
XFILLER_128_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17058_ _17096_/A _17058_/B vssd1 vssd1 vccd1 vccd1 _17062_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08900_ _08900_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__nor2_2
XFILLER_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16009_ _17119_/B _17163_/A2 _16008_/X vssd1 vssd1 vccd1 vccd1 _16017_/A sky130_fd_sc_hd__o21ba_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__nor2_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08831_ _08831_/A _08831_/B _08831_/C vssd1 vssd1 vccd1 vccd1 _08832_/C sky130_fd_sc_hd__nor3_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08760_/Y _16302_/A _08758_/X vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__o21ai_4
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09314_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09316_/C sky130_fd_sc_hd__xnor2_4
XFILLER_55_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09245_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _09245_/Y sky130_fd_sc_hd__nand3_2
XFILLER_166_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09176_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09357_/C sky130_fd_sc_hd__xnor2_1
XFILLER_147_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ _10970_/A _10659_/D _09895_/A _09893_/Y vssd1 vssd1 vccd1 vccd1 _10021_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11971_ _11971_/A _11971_/B vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__and2_1
XFILLER_5_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13710_ _13814_/A _13710_/B _13817_/A _13710_/D vssd1 vssd1 vccd1 vccd1 _13814_/B
+ sky130_fd_sc_hd__nor4_4
XTAP_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10922_ _14787_/A _15463_/A _15381_/A _14786_/A vssd1 vssd1 vccd1 vccd1 _10922_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14690_ _14691_/A _14691_/B vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__nor2_1
XTAP_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13641_ _13641_/A _13745_/B _13745_/D _14175_/B vssd1 vssd1 vccd1 vccd1 _13642_/B
+ sky130_fd_sc_hd__and4_1
X_10853_ _10854_/A _10852_/Y _11124_/C _11334_/C vssd1 vssd1 vccd1 vccd1 _10874_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_188_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _16361_/A _16361_/B vssd1 vssd1 vccd1 vccd1 _16443_/B sky130_fd_sc_hd__nand2b_1
XFILLER_169_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13572_ _14248_/A _16789_/A _13572_/C vssd1 vssd1 vccd1 vccd1 _13702_/B sky130_fd_sc_hd__nand3_2
XFILLER_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10784_ _10784_/A _10784_/B vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__xnor2_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15311_ _16304_/A _15311_/B _14801_/X vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__or3b_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12522_/A _12522_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12524_/B sky130_fd_sc_hd__o21ai_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16382_/B _16562_/C vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__nand2b_4
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _15454_/A _15242_/B _15242_/C vssd1 vssd1 vccd1 vccd1 _15257_/A sky130_fd_sc_hd__and3_1
X_12454_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12454_/Y sky130_fd_sc_hd__nand3_2
XFILLER_138_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _11405_/A vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__inv_2
X_15173_ _15235_/C _15173_/B vssd1 vssd1 vccd1 vccd1 _15173_/Y sky130_fd_sc_hd__nand2_1
X_12385_ _12051_/Y _12053_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14124_ _14278_/A _14125_/B vssd1 vssd1 vccd1 vccd1 _14124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ _11437_/B _11334_/C _11391_/B _11629_/A vssd1 vssd1 vccd1 vccd1 _11337_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_141_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14055_ _14158_/B _14055_/B vssd1 vssd1 vccd1 vccd1 _14057_/B sky130_fd_sc_hd__nor2_2
X_11267_ _11377_/B _14899_/A _14906_/B _11266_/A vssd1 vssd1 vccd1 vccd1 _11268_/D
+ sky130_fd_sc_hd__a22o_1
X_13006_ _12693_/X _12840_/B _12838_/Y vssd1 vssd1 vccd1 vccd1 _13006_/Y sky130_fd_sc_hd__a21oi_1
X_10218_ _10216_/A _10216_/B _10216_/C vssd1 vssd1 vccd1 vccd1 _10219_/C sky130_fd_sc_hd__a21oi_2
X_11198_ _11198_/A _11198_/B vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__xnor2_4
XFILLER_67_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__nor2_2
XFILLER_153_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14957_ _12054_/A _09892_/D _10657_/C vssd1 vssd1 vccd1 vccd1 _15056_/B sky130_fd_sc_hd__a21o_1
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13908_ _14008_/A _13908_/B _13908_/C vssd1 vssd1 vccd1 vccd1 _14027_/B sky130_fd_sc_hd__and3_1
X_14888_ _14888_/A _14888_/B _14888_/C _14888_/D vssd1 vssd1 vccd1 vccd1 _15025_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16627_ _16627_/A _16627_/B vssd1 vssd1 vccd1 vccd1 _16628_/B sky130_fd_sc_hd__xnor2_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13839_ _14841_/B _14840_/B _14666_/S vssd1 vssd1 vccd1 vccd1 _13839_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16558_ _16558_/A _16558_/B _16558_/C vssd1 vssd1 vccd1 vccd1 _16560_/A sky130_fd_sc_hd__nand3_4
X_15509_ _15510_/A _15510_/B vssd1 vssd1 vccd1 vccd1 _15509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16489_ _14775_/X _16580_/A2 _16733_/B1 _16480_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16489_/X sky130_fd_sc_hd__a221o_1
X_09030_ _09030_/A _11867_/B _12166_/B _09030_/D vssd1 vssd1 vccd1 vccd1 _09031_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_191_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__nand2_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout804 _10839_/D vssd1 vssd1 vccd1 vccd1 _10736_/C sky130_fd_sc_hd__clkbuf_16
Xfanout815 _12502_/B1 vssd1 vssd1 vccd1 vccd1 _15530_/A sky130_fd_sc_hd__buf_6
Xfanout826 _12465_/B vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__buf_6
X_09863_ _09863_/A _09863_/B _09863_/C vssd1 vssd1 vccd1 vccd1 _09864_/C sky130_fd_sc_hd__nand3_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout837 _12463_/D vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__buf_8
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout848 _12295_/D vssd1 vssd1 vccd1 vccd1 _12127_/C sky130_fd_sc_hd__buf_8
XFILLER_140_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout859 _10805_/C vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__buf_6
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08814_ _08814_/A _08814_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__xnor2_4
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _10062_/A _09947_/B _09640_/A _09638_/Y vssd1 vssd1 vccd1 vccd1 _09795_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08745_ _12068_/B _12068_/D _12637_/D _12068_/A vssd1 vssd1 vccd1 vccd1 _08748_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09228_ _09228_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__nor2_4
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09159_ _10542_/A _11813_/B vssd1 vssd1 vccd1 vccd1 _14948_/B sky130_fd_sc_hd__and2_2
XFILLER_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12170_ _12170_/A _12170_/B vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11121_/A _11126_/A _11121_/C vssd1 vssd1 vccd1 vccd1 _11130_/B sky130_fd_sc_hd__or3_4
XFILLER_104_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _11047_/Y _11050_/X _11041_/Y _11042_/X vssd1 vssd1 vccd1 vccd1 _11055_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10005_/B sky130_fd_sc_hd__xnor2_4
XFILLER_27_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15860_ _15861_/A _15861_/B vssd1 vssd1 vccd1 vccd1 _15980_/A sky130_fd_sc_hd__and2_1
XFILLER_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14811_ _15895_/B _15895_/C _09424_/X vssd1 vssd1 vccd1 vccd1 _16005_/C sky130_fd_sc_hd__a21o_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15791_ _15788_/Y _15790_/X _16911_/A vssd1 vssd1 vccd1 vccd1 _15791_/Y sky130_fd_sc_hd__o21ai_1
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17530_ fanout932/X _17530_/D vssd1 vssd1 vccd1 vccd1 _17530_/Q sky130_fd_sc_hd__dfxtp_4
X_14742_ _14742_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14743_/B sky130_fd_sc_hd__nand2_1
X_11954_ _12488_/A _12158_/C vssd1 vssd1 vccd1 vccd1 _11956_/C sky130_fd_sc_hd__nand2_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10905_ _10905_/A _10905_/B _11027_/C _11027_/D vssd1 vssd1 vccd1 vccd1 _10907_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_189_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14673_ _14708_/B _14829_/B vssd1 vssd1 vccd1 vccd1 _17167_/A sky130_fd_sc_hd__nand2_8
X_17461_ fanout938/X _17461_/D vssd1 vssd1 vccd1 vccd1 _17461_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_83_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11885_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _12118_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16412_ _16318_/A _16504_/B _16316_/B vssd1 vssd1 vccd1 vccd1 _16414_/B sky130_fd_sc_hd__o21ai_4
X_13624_ _14839_/A _13624_/B vssd1 vssd1 vccd1 vccd1 _13624_/X sky130_fd_sc_hd__or2_2
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10836_ _10836_/A _10850_/A vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__or2_4
X_17392_ input41/X _17396_/A2 _17391_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17524_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16343_ _16344_/A _16344_/B vssd1 vssd1 vccd1 vccd1 _16345_/A sky130_fd_sc_hd__and2_1
X_13555_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _13556_/B sky130_fd_sc_hd__and2_1
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10767_ _10766_/C _11725_/A _10667_/Y _10692_/X vssd1 vssd1 vccd1 vccd1 _10774_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_157_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12508_/C sky130_fd_sc_hd__xnor2_2
X_16274_ _16181_/A _16279_/C _16180_/B _16160_/X vssd1 vssd1 vccd1 vccd1 _16276_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _13486_/A _13603_/B _13486_/C vssd1 vssd1 vccd1 vccd1 _13486_/X sky130_fd_sc_hd__and3_4
XFILLER_139_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10698_ _11027_/B _10809_/D _10697_/B _10694_/X vssd1 vssd1 vccd1 vccd1 _10701_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_157_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15225_ _15225_/A _15225_/B vssd1 vssd1 vccd1 vccd1 _15226_/B sky130_fd_sc_hd__xnor2_4
XFILLER_32_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12437_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__nand3_2
XFILLER_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15156_ _15157_/A _15157_/B vssd1 vssd1 vccd1 vccd1 _15222_/B sky130_fd_sc_hd__nand2b_2
X_12368_ _12368_/A _12368_/B vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__xnor2_4
XFILLER_114_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14108_/A _14108_/B vssd1 vssd1 vccd1 vccd1 _14197_/A sky130_fd_sc_hd__nand2b_1
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11319_ _11268_/A _11268_/B _11268_/C _11268_/D vssd1 vssd1 vccd1 vccd1 _11320_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15087_ _15161_/A _15087_/B vssd1 vssd1 vccd1 vccd1 _15091_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12299_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12300_/B sky130_fd_sc_hd__and2_1
X_14038_ _15457_/A _14036_/X _14037_/X vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_45_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15989_ _15989_/A _15989_/B _15987_/X vssd1 vssd1 vccd1 vccd1 _15990_/B sky130_fd_sc_hd__or3b_1
XFILLER_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09013_ _09013_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _09014_/B sky130_fd_sc_hd__nor2_2
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout601 _15062_/S0 vssd1 vssd1 vccd1 vccd1 _12060_/S sky130_fd_sc_hd__buf_6
Xfanout612 _14554_/B vssd1 vssd1 vccd1 vccd1 _14708_/C sky130_fd_sc_hd__buf_6
XFILLER_59_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09915_ _09915_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__or2_2
XFILLER_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout623 _17508_/Q vssd1 vssd1 vccd1 vccd1 _14829_/B sky130_fd_sc_hd__buf_8
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout634 _09350_/B vssd1 vssd1 vccd1 vccd1 _12595_/C sky130_fd_sc_hd__buf_6
Xfanout645 _13908_/B vssd1 vssd1 vccd1 vccd1 _14002_/B sky130_fd_sc_hd__buf_8
Xfanout656 _16974_/A vssd1 vssd1 vccd1 vccd1 _14545_/D sky130_fd_sc_hd__buf_8
Xfanout667 _17503_/Q vssd1 vssd1 vccd1 vccd1 _14155_/B sky130_fd_sc_hd__buf_6
X_09846_ _11026_/A _10392_/D vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__nand2_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout678 fanout686/X vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__buf_12
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout689 _14863_/B vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__nor2_4
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _15008_/B vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__inv_6
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11670_ _15524_/C _11690_/A _11670_/C vssd1 vssd1 vccd1 vccd1 _11671_/B sky130_fd_sc_hd__and3b_1
XFILLER_187_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10621_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__nor2_2
XFILLER_168_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _13339_/A _13339_/B _13339_/C vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__o21ai_2
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10552_ _10566_/A _10523_/Y _10538_/Y _10550_/X vssd1 vssd1 vccd1 vccd1 _10553_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ _13271_/A _13271_/B vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__or2_1
XFILLER_108_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ _10597_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__nand2_1
XFILLER_185_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15010_ _11651_/A _14794_/B _15008_/B _14794_/A vssd1 vssd1 vccd1 vccd1 _15011_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12222_ _12220_/X _12221_/X _17367_/A vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12153_ _11917_/X _11947_/X _12316_/B _12152_/X vssd1 vssd1 vccd1 vccd1 _12360_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _11104_/A _11104_/B _11104_/C vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__nand3_2
XFILLER_190_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16961_ _16931_/X _16932_/X _16960_/X vssd1 vssd1 vccd1 vccd1 _17014_/A sky130_fd_sc_hd__a21o_1
X_12084_ _12085_/A _12085_/B _12085_/C vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__a21o_4
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15912_ _16352_/B _16129_/B vssd1 vssd1 vccd1 vccd1 _16939_/B sky130_fd_sc_hd__nand2_4
X_11035_ _11035_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11038_/A sky130_fd_sc_hd__xor2_4
X_16892_ _16827_/A _16827_/C _16758_/B _16935_/A vssd1 vssd1 vccd1 vccd1 _16893_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _16758_/A _16020_/B vssd1 vssd1 vccd1 vccd1 _16355_/B sky130_fd_sc_hd__and2_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15774_ _15774_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15775_/B sky130_fd_sc_hd__nand2_1
X_12986_ _12985_/A _12985_/B _12985_/C vssd1 vssd1 vccd1 vccd1 _12986_/Y sky130_fd_sc_hd__o21ai_4
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ fanout925/X _17513_/D vssd1 vssd1 vccd1 vccd1 _17513_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _14727_/B vssd1 vssd1 vccd1 vccd1 _14725_/Y sky130_fd_sc_hd__inv_2
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _11937_/A _11937_/B vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__xnor2_4
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ fanout934/X _17444_/D vssd1 vssd1 vccd1 vccd1 _17444_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14656_ _14691_/A _14656_/B vssd1 vssd1 vccd1 vccd1 _14658_/C sky130_fd_sc_hd__and2_1
X_11868_ _11868_/A _12093_/A vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__nor2_1
XFILLER_162_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13607_ _13607_/A _13607_/B _13607_/C vssd1 vssd1 vccd1 vccd1 _13607_/X sky130_fd_sc_hd__or3_2
X_10819_ _11095_/A _11240_/A _11097_/D _11423_/C vssd1 vssd1 vccd1 vccd1 _10822_/A
+ sky130_fd_sc_hd__and4_2
X_17375_ _17375_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__or2_1
X_14587_ _14629_/C _14587_/B vssd1 vssd1 vccd1 vccd1 _14587_/Y sky130_fd_sc_hd__nand2_1
X_11799_ _14888_/C _11799_/B vssd1 vssd1 vccd1 vccd1 _11800_/D sky130_fd_sc_hd__or2_2
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16326_ _16326_/A _16326_/B vssd1 vssd1 vccd1 vccd1 _16328_/B sky130_fd_sc_hd__xor2_1
XFILLER_146_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13538_ _13538_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__xnor2_4
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16257_ _16257_/A _16257_/B vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__xor2_2
XFILLER_174_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13469_ _13469_/A _13469_/B vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15530_/A _15262_/C _15208_/C _15208_/D vssd1 vssd1 vccd1 vccd1 _15208_/X
+ sky130_fd_sc_hd__or4_4
X_16188_ _16188_/A _16188_/B _16188_/C vssd1 vssd1 vccd1 vccd1 _16189_/B sky130_fd_sc_hd__nor3_1
XFILLER_160_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15139_ _15147_/A _17614_/Q _15147_/C vssd1 vssd1 vccd1 vccd1 _15141_/B sky130_fd_sc_hd__nor3_2
XFILLER_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _11026_/A _10736_/C _09701_/C vssd1 vssd1 vccd1 vccd1 _09702_/A sky130_fd_sc_hd__a21oi_1
XFILLER_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _09632_/B _09632_/A vssd1 vssd1 vccd1 vccd1 _09631_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09562_ _09556_/A _09558_/B _09556_/B vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__o21ba_4
XFILLER_64_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _09926_/A _11813_/B _14949_/A vssd1 vssd1 vccd1 vccd1 _09619_/B sky130_fd_sc_hd__and3_2
XFILLER_169_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout420 _17528_/Q vssd1 vssd1 vccd1 vccd1 _14776_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_28_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout431 _11027_/A vssd1 vssd1 vccd1 vccd1 _11867_/B sky130_fd_sc_hd__buf_12
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout442 _12079_/A vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__buf_12
Xfanout453 _09566_/A vssd1 vssd1 vccd1 vccd1 _10905_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout464 _11791_/C vssd1 vssd1 vccd1 vccd1 _16809_/A sky130_fd_sc_hd__buf_6
Xfanout475 _12595_/A vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__clkbuf_4
Xfanout486 _15262_/B vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__buf_6
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _09813_/A _09813_/C _09813_/B vssd1 vssd1 vccd1 vccd1 _09829_/Y sky130_fd_sc_hd__a21oi_4
Xfanout497 _09748_/A vssd1 vssd1 vccd1 vccd1 _11895_/A sky130_fd_sc_hd__buf_6
XFILLER_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12840_ _12838_/Y _12840_/B vssd1 vssd1 vccd1 vccd1 _13003_/B sky130_fd_sc_hd__nand2b_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12771_/A _12771_/B vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__nor2_1
XFILLER_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _14512_/A vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__inv_2
X_11722_ _11722_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11731_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _15143_/A _15208_/C _15541_/A vssd1 vssd1 vccd1 vccd1 _15492_/B sky130_fd_sc_hd__a21bo_4
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14441_ _14441_/A _14441_/B vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _15056_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__nor2_2
XFILLER_187_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _11006_/A _11006_/B _10963_/D _11005_/B vssd1 vssd1 vccd1 vccd1 _10607_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14372_ _14372_/A _14372_/B _14372_/C vssd1 vssd1 vccd1 vccd1 _14373_/B sky130_fd_sc_hd__or3_1
XFILLER_167_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17160_ _12442_/B _17140_/B _17140_/A vssd1 vssd1 vccd1 vccd1 _17160_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _11584_/A _11584_/B _11583_/Y vssd1 vssd1 vccd1 vccd1 _11620_/A sky130_fd_sc_hd__nor3b_4
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13323_ _17421_/A _13434_/C vssd1 vssd1 vccd1 vccd1 _13324_/B sky130_fd_sc_hd__nand2_1
X_16111_ _17156_/B _16111_/B _16111_/C vssd1 vssd1 vccd1 vccd1 _16111_/X sky130_fd_sc_hd__or3_1
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ _10535_/A _10644_/A vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__or2_4
XFILLER_156_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17091_ _17091_/A _17118_/B vssd1 vssd1 vccd1 vccd1 _17092_/B sky130_fd_sc_hd__or2_1
XFILLER_127_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16042_ _16041_/A _16041_/B _16041_/C vssd1 vssd1 vccd1 vccd1 _16043_/B sky130_fd_sc_hd__o21ai_1
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13254_ _13118_/A _13119_/Y _13252_/A _13253_/Y vssd1 vssd1 vccd1 vccd1 _13256_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_170_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10466_ _10469_/A _10469_/B _10469_/C vssd1 vssd1 vccd1 vccd1 _10470_/A sky130_fd_sc_hd__o21a_1
XFILLER_89_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ _12010_/A _12010_/B _12006_/X vssd1 vssd1 vccd1 vccd1 _12206_/C sky130_fd_sc_hd__a21oi_4
XFILLER_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ _13186_/A _13186_/B vssd1 vssd1 vccd1 vccd1 _13326_/B sky130_fd_sc_hd__nor2_2
XFILLER_123_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__xnor2_4
XFILLER_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12136_ _12136_/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12138_/C sky130_fd_sc_hd__nor2_4
XFILLER_123_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16944_ _16994_/B _16944_/B vssd1 vssd1 vccd1 vccd1 _16947_/A sky130_fd_sc_hd__nand2_4
X_12067_ _12068_/B _12068_/C _12068_/D _12068_/A vssd1 vssd1 vccd1 vccd1 _12070_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ _11018_/A _11018_/B vssd1 vssd1 vccd1 vccd1 _11020_/B sky130_fd_sc_hd__nor2_4
X_16875_ _16917_/A _16862_/X _16863_/Y _16874_/X vssd1 vssd1 vccd1 vccd1 _16875_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15826_ _15827_/A _15827_/B vssd1 vssd1 vccd1 vccd1 _15826_/Y sky130_fd_sc_hd__nor2_1
XTAP_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15757_ _15668_/A _15668_/B _15665_/Y vssd1 vssd1 vccd1 vccd1 _15759_/B sky130_fd_sc_hd__o21a_2
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12805_/A _12807_/B _12805_/B vssd1 vssd1 vccd1 vccd1 _12971_/B sky130_fd_sc_hd__o21ba_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14708_ _14738_/A _14708_/B _14708_/C _14708_/D vssd1 vssd1 vccd1 vccd1 _14713_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_166_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15688_ _16281_/A _16589_/B _15686_/Y vssd1 vssd1 vccd1 vccd1 _15689_/B sky130_fd_sc_hd__a21o_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ input28/X input29/X wire217/X vssd1 vssd1 vccd1 vccd1 _17428_/D sky130_fd_sc_hd__a21boi_1
X_14639_ _14593_/B _14641_/C _14641_/D _14593_/A vssd1 vssd1 vccd1 vccd1 _14642_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_119_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17358_ _13300_/C _17360_/A2 _17357_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17508_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _16735_/A _13943_/X _14926_/X _14990_/X vssd1 vssd1 vccd1 vccd1 _16310_/D
+ sky130_fd_sc_hd__o22a_1
X_17289_ _17573_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17289_/X sky130_fd_sc_hd__and2_1
XFILLER_161_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08993_ _12845_/S _12592_/C _08993_/C vssd1 vssd1 vccd1 vccd1 _08994_/B sky130_fd_sc_hd__and3_2
XFILLER_173_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09614_ _09614_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09746_/C sky130_fd_sc_hd__xnor2_4
XFILLER_141_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09476_ _09478_/B _09603_/A _09478_/A vssd1 vssd1 vccd1 vccd1 _09476_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_180_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10319_/A _10319_/Y _10193_/B _10229_/X vssd1 vssd1 vccd1 vccd1 _10336_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10251_ _10251_/A _10251_/B vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__xnor2_4
XFILLER_152_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _10183_/A _10181_/Y _12398_/S _10309_/B vssd1 vssd1 vccd1 vccd1 _10307_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14990_ _15537_/B _14989_/X _15901_/S vssd1 vssd1 vccd1 vccd1 _14990_/X sky130_fd_sc_hd__mux2_2
Xfanout250 _15794_/A vssd1 vssd1 vccd1 vccd1 _17070_/B sky130_fd_sc_hd__buf_12
XFILLER_182_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout261 _15147_/Y vssd1 vssd1 vccd1 vccd1 _17038_/C sky130_fd_sc_hd__clkbuf_8
Xfanout272 _17063_/A vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__buf_6
X_13941_ _14122_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _14032_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout283 _15038_/A vssd1 vssd1 vccd1 vccd1 _15096_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout294 _08721_/Y vssd1 vssd1 vccd1 vccd1 _12862_/S sky130_fd_sc_hd__buf_6
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16660_ _16651_/A _16806_/A2 _16659_/X vssd1 vssd1 vccd1 vccd1 _17564_/D sky130_fd_sc_hd__a21oi_1
X_13872_ _13873_/A _13873_/B vssd1 vssd1 vccd1 vccd1 _14018_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15611_ _15522_/A _15521_/B _15519_/X vssd1 vssd1 vccd1 vccd1 _15611_/X sky130_fd_sc_hd__a21o_2
X_12823_ _12822_/B _12823_/B vssd1 vssd1 vccd1 vccd1 _12824_/B sky130_fd_sc_hd__nand2b_1
X_16591_ _16814_/B _16935_/B _16591_/C vssd1 vssd1 vccd1 vccd1 _16686_/B sky130_fd_sc_hd__and3_2
XFILLER_90_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15542_ _14785_/X _15899_/A2 _16008_/B1 _15541_/A _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15542_/X sky130_fd_sc_hd__a221o_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12754_ _12754_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12755_/C sky130_fd_sc_hd__xnor2_2
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11705_/A _15888_/A vssd1 vssd1 vccd1 vccd1 _11705_/Y sky130_fd_sc_hd__nand2_1
X_15473_ _16127_/A _16246_/A _16604_/B _15475_/A vssd1 vssd1 vccd1 vccd1 _15473_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12685_/Y sky130_fd_sc_hd__nand2_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17212_ _17438_/Q _17266_/A2 _17210_/X _17211_/X _17322_/C1 vssd1 vssd1 vccd1 vccd1
+ _17438_/D sky130_fd_sc_hd__o221a_1
X_14424_ _14424_/A _14424_/B vssd1 vssd1 vccd1 vccd1 _14469_/A sky130_fd_sc_hd__nor2_1
X_11636_ _15116_/A _11675_/B _15553_/A _15175_/A vssd1 vssd1 vccd1 vccd1 _11637_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17143_ _16653_/A _14734_/B _17142_/X vssd1 vssd1 vccd1 vccd1 _17143_/X sky130_fd_sc_hd__o21a_1
X_14355_ _14763_/S _14353_/Y _14354_/X _14288_/Y vssd1 vssd1 vccd1 vccd1 _17596_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11558_/A _11558_/C _11558_/B vssd1 vssd1 vccd1 vccd1 _11568_/C sky130_fd_sc_hd__a21o_1
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _13308_/C sky130_fd_sc_hd__xnor2_4
X_10518_ _10384_/X _10475_/Y _10485_/X _10499_/A vssd1 vssd1 vccd1 vccd1 _10519_/C
+ sky130_fd_sc_hd__o211a_2
X_14286_ _12545_/X _12553_/B _14421_/S vssd1 vssd1 vccd1 vccd1 _16653_/B sky130_fd_sc_hd__mux2_4
X_17074_ _14765_/X _17162_/A2 _16974_/B _17065_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _17074_/X sky130_fd_sc_hd__a221o_1
X_11498_ _11495_/A _11495_/B _11532_/A vssd1 vssd1 vccd1 vccd1 _11499_/C sky130_fd_sc_hd__o21ba_2
XFILLER_137_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16025_ _16025_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16026_/B sky130_fd_sc_hd__nor2_2
X_13237_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__or2_2
X_10449_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__nand2_4
XFILLER_152_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _13298_/A _13300_/D _13169_/D _17391_/A vssd1 vssd1 vccd1 vccd1 _13170_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12119_ _11905_/X _11909_/A _12309_/A _12118_/Y vssd1 vssd1 vccd1 vccd1 _12309_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_111_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13099_ _13099_/A _13099_/B vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16927_ _16582_/A _15537_/X _16926_/Y vssd1 vssd1 vccd1 vccd1 _16927_/X sky130_fd_sc_hd__o21a_1
XFILLER_133_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ _14383_/A _17134_/C _16859_/A vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15809_ _15805_/Y _15806_/Y _15808_/Y vssd1 vssd1 vccd1 vccd1 _15809_/Y sky130_fd_sc_hd__o21ai_2
X_16789_ _16789_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _16789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09330_ _09462_/A _09468_/A _09462_/C vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__o21ai_4
XFILLER_34_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__nand2_1
XFILLER_178_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09192_ _11953_/B _12174_/D _12129_/B _11953_/A vssd1 vssd1 vccd1 vccd1 _09194_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08976_ _12770_/A _11920_/B _10446_/B _09172_/B vssd1 vssd1 vccd1 vccd1 _09238_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_103_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09528_ _09391_/C _09399_/Y _09458_/X _09628_/A vssd1 vssd1 vccd1 vccd1 _09528_/Y
+ sky130_fd_sc_hd__a211oi_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09334_/A _09334_/B _09334_/C vssd1 vssd1 vccd1 vccd1 _09459_/Y sky130_fd_sc_hd__a21oi_4
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ _12303_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__nand2b_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11421_ _11396_/A _11396_/C _11396_/B vssd1 vssd1 vccd1 vccd1 _11421_/Y sky130_fd_sc_hd__a21oi_4
X_14140_ _14213_/B _14052_/B _14141_/D _14290_/A vssd1 vssd1 vccd1 vccd1 _14142_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11352_ _11352_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__xnor2_2
XFILLER_193_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10303_ _10305_/B _10305_/C _10305_/A vssd1 vssd1 vccd1 vccd1 _10303_/Y sky130_fd_sc_hd__a21oi_4
X_14071_ _14071_/A _14071_/B vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__xor2_1
X_11283_ _11283_/A _11283_/B _11333_/A vssd1 vssd1 vccd1 vccd1 _11284_/B sky130_fd_sc_hd__or3_1
XFILLER_3_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13022_ _17401_/A _13564_/C _12872_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _13024_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_180_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10234_ _10234_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__nor2_4
XFILLER_140_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10165_ _10971_/A _10647_/D _10745_/D _10525_/A vssd1 vssd1 vccd1 vccd1 _10165_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10096_ _09968_/B _09970_/A _09968_/A vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__o21ai_4
X_14973_ _14886_/X _14972_/X _15056_/A vssd1 vssd1 vccd1 vccd1 _15749_/A sky130_fd_sc_hd__a21oi_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16712_ _16786_/A _16712_/B vssd1 vssd1 vccd1 vccd1 _16714_/B sky130_fd_sc_hd__and2_1
X_13924_ _13925_/A _13925_/B _13925_/C vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__a21o_2
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16643_ _16643_/A vssd1 vssd1 vccd1 vccd1 _16643_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13855_ _13856_/A _13856_/B vssd1 vssd1 vccd1 vccd1 _13961_/A sky130_fd_sc_hd__and2b_1
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12806_ _17415_/A _13434_/D vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__nand2_4
X_16574_ _16917_/A _16574_/B vssd1 vssd1 vccd1 vccd1 _16574_/Y sky130_fd_sc_hd__nand2_1
X_13786_ _13787_/A _13787_/B vssd1 vssd1 vccd1 vccd1 _13915_/A sky130_fd_sc_hd__and2b_1
X_10998_ _11159_/A _10998_/B vssd1 vssd1 vccd1 vccd1 _10999_/C sky130_fd_sc_hd__and2_2
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _15525_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15525_/X sky130_fd_sc_hd__and2_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12737_ _12737_/A _12737_/B vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__xnor2_2
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15456_ _15456_/A _16304_/A _15455_/X vssd1 vssd1 vccd1 vccd1 _15467_/B sky130_fd_sc_hd__or3b_2
X_12668_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _14340_/B _14342_/A _14424_/B _14406_/Y vssd1 vssd1 vccd1 vccd1 _14473_/A
+ sky130_fd_sc_hd__a211o_4
X_11619_ _11584_/A _11584_/B _11583_/Y vssd1 vssd1 vccd1 vccd1 _11620_/C sky130_fd_sc_hd__o21ba_1
X_15387_ _16115_/A _15463_/B _15381_/Y _15383_/X _15386_/Y vssd1 vssd1 vccd1 vccd1
+ _15387_/X sky130_fd_sc_hd__o311a_1
XFILLER_190_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ _12599_/A _12599_/B vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__and2_2
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17126_ _17127_/A _17127_/B vssd1 vssd1 vccd1 vccd1 _17128_/A sky130_fd_sc_hd__or2_1
XFILLER_184_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14338_ _14222_/A _14265_/B _14336_/X _14337_/Y vssd1 vssd1 vccd1 vccd1 _14340_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17057_ _17056_/B _17057_/B vssd1 vssd1 vccd1 vccd1 _17058_/B sky130_fd_sc_hd__and2b_1
XFILLER_132_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14269_ _14270_/A _14270_/B _14270_/C vssd1 vssd1 vccd1 vccd1 _14350_/A sky130_fd_sc_hd__a21oi_2
XFILLER_132_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ _16005_/B _14928_/Y _16008_/B1 _16014_/A _16008_/C1 vssd1 vssd1 vccd1 vccd1
+ _16008_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08830_ _08830_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08832_/B sky130_fd_sc_hd__nand2_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _11867_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _16302_/A sky130_fd_sc_hd__nand2_8
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09313_ _09338_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09391_/B sky130_fd_sc_hd__or2_2
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _11990_/B sky130_fd_sc_hd__a21o_4
XFILLER_167_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _09357_/A _09174_/Y _09502_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _09364_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__xnor2_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11970_ _11970_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__nand2_1
XTAP_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10921_ _14786_/A _15463_/A vssd1 vssd1 vccd1 vccd1 _14805_/A sky130_fd_sc_hd__nand2_1
XTAP_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13640_ _13745_/B _13745_/D _14175_/B _13641_/A vssd1 vssd1 vccd1 vccd1 _13642_/A
+ sky130_fd_sc_hd__a22oi_2
X_10852_ _11122_/B _11335_/B _11391_/B _11266_/A vssd1 vssd1 vccd1 vccd1 _10852_/Y
+ sky130_fd_sc_hd__a22oi_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13571_/A _13702_/A vssd1 vssd1 vccd1 vccd1 _13572_/C sky130_fd_sc_hd__and2_1
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10783_ _10784_/A _10784_/B _11768_/B vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__o21ba_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _14801_/A _14801_/B _14801_/C vssd1 vssd1 vccd1 vccd1 _15311_/B sky130_fd_sc_hd__o21a_1
X_12522_ _12522_/A _12522_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12524_/A sky130_fd_sc_hd__or3_1
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16290_ _16290_/A _16290_/B _16290_/C vssd1 vssd1 vccd1 vccd1 _16562_/C sky130_fd_sc_hd__or3_4
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _15241_/A _15241_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15242_/C sky130_fd_sc_hd__nand3_1
X_12453_ _12454_/A _12454_/B _12454_/C vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__a21o_2
XFILLER_166_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _11406_/A _11406_/B vssd1 vssd1 vccd1 vccd1 _11405_/A sky130_fd_sc_hd__or2_1
X_12384_ _12382_/X _12383_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__mux2_1
X_15172_ _15106_/A _11683_/B _16207_/B vssd1 vssd1 vccd1 vccd1 _15173_/B sky130_fd_sc_hd__a21oi_1
XFILLER_181_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14123_ _13939_/Y _14281_/A _14121_/X vssd1 vssd1 vccd1 vccd1 _14125_/B sky130_fd_sc_hd__a21oi_1
X_11335_ _11630_/A _11335_/B vssd1 vssd1 vccd1 vccd1 _11386_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14054_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14055_/B sky130_fd_sc_hd__and2_1
XFILLER_140_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11266_ _11266_/A _11377_/B _14899_/A _14906_/B vssd1 vssd1 vccd1 vccd1 _11268_/C
+ sky130_fd_sc_hd__nand4_2
X_10217_ _10209_/A _10210_/A _10209_/B _10211_/Y vssd1 vssd1 vccd1 vccd1 _10219_/B
+ sky130_fd_sc_hd__o31a_2
X_13005_ _13005_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__and2_1
X_11197_ _11198_/B _11198_/A vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__and2b_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10148_ _10148_/A _10148_/B _10148_/C vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__nor3_1
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10079_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__nand2_2
X_14956_ _14956_/A _14956_/B vssd1 vssd1 vccd1 vccd1 _14956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_48_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13907_ _14027_/A _13907_/B vssd1 vssd1 vccd1 vccd1 _13908_/C sky130_fd_sc_hd__nor2_1
XFILLER_63_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14887_ _14888_/A _14887_/B vssd1 vssd1 vccd1 vccd1 _14887_/Y sky130_fd_sc_hd__nor2_2
XFILLER_63_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16626_ _16624_/X _16626_/B vssd1 vssd1 vccd1 vccd1 _16627_/B sky130_fd_sc_hd__and2b_2
XFILLER_23_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13838_ _12857_/X _12861_/X _13838_/S vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__mux2_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16557_ _16557_/A _16557_/B _16557_/C vssd1 vssd1 vccd1 vccd1 _16558_/C sky130_fd_sc_hd__or3_4
X_13769_ _13770_/A _13770_/B _13770_/C vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__o21ai_4
XFILLER_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15508_ _15687_/A _16041_/A vssd1 vssd1 vccd1 vccd1 _15510_/B sky130_fd_sc_hd__or2_4
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16488_ _16480_/A _16400_/B _16487_/Y vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__o21ai_1
X_15439_ _15439_/A _15439_/B vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__xor2_4
XFILLER_117_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17109_ _17140_/A _17139_/B _17109_/C vssd1 vssd1 vccd1 vccd1 _17113_/A sky130_fd_sc_hd__or3_1
XFILLER_171_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__or2_1
XFILLER_113_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout805 _15617_/A vssd1 vssd1 vccd1 vccd1 _15624_/A sky130_fd_sc_hd__buf_4
Xfanout816 _12502_/B1 vssd1 vssd1 vccd1 vccd1 _11335_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_113_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09862_/A _09862_/B vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__xnor2_2
Xfanout827 _17486_/Q vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__clkbuf_16
Xfanout838 _12463_/D vssd1 vssd1 vccd1 vccd1 _09937_/B sky130_fd_sc_hd__buf_6
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout849 _17483_/Q vssd1 vssd1 vccd1 vccd1 _12295_/D sky130_fd_sc_hd__clkbuf_8
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08813_ _12245_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _08814_/B sky130_fd_sc_hd__nand2_4
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__nor2_2
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08744_ _15071_/A _14836_/A _08743_/Y vssd1 vssd1 vccd1 vccd1 _17611_/D sky130_fd_sc_hd__a21o_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09227_ _09227_/A _09227_/B _09227_/C vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__and3_1
XFILLER_107_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09158_ _09165_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__nor2_2
XFILLER_108_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09089_ _09317_/A _09323_/A _09317_/C vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__o21ai_2
X_11120_ _11121_/A _11121_/C vssd1 vssd1 vccd1 vccd1 _11126_/B sky130_fd_sc_hd__nor2_2
XFILLER_190_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11051_ _11051_/A _11051_/B _11051_/C vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__nand3_2
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10002_ _10003_/B _10003_/A vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__nand2b_1
XFILLER_88_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1004 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14810_ _15801_/B _15802_/A _16809_/B vssd1 vssd1 vccd1 vccd1 _15895_/C sky130_fd_sc_hd__a21o_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15790_ _15610_/Y _15611_/X _15700_/A _15789_/X vssd1 vssd1 vccd1 vccd1 _15790_/X
+ sky130_fd_sc_hd__a31o_2
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _14742_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__or2_1
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11953_ _11953_/A _11953_/B _12340_/B _12338_/C vssd1 vssd1 vccd1 vccd1 _12163_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ fanout942/X _17460_/D vssd1 vssd1 vccd1 vccd1 _17460_/Q sky130_fd_sc_hd__dfxtp_4
X_10904_ _10905_/B _10904_/B _11423_/C _11605_/B vssd1 vssd1 vccd1 vccd1 _11107_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_72_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _14633_/A _14631_/A _14669_/B _14671_/X vssd1 vssd1 vccd1 vccd1 _14701_/A
+ sky130_fd_sc_hd__a31oi_4
X_11884_ _11884_/A _11884_/B vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__xnor2_4
XFILLER_189_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16411_ _16411_/A _16505_/B vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__and2_2
XFILLER_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13623_ _12705_/X _12709_/B _13627_/S vssd1 vssd1 vccd1 vccd1 _13624_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10835_ _10836_/A _10834_/Y _11124_/C _11135_/B vssd1 vssd1 vccd1 vccd1 _10850_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17391_ _17391_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17391_/X sky130_fd_sc_hd__or2_1
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16342_ _16342_/A _16342_/B vssd1 vssd1 vccd1 vccd1 _16344_/B sky130_fd_sc_hd__xnor2_1
X_13554_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _13680_/B sky130_fd_sc_hd__nor2_2
XFILLER_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10766_ _10764_/X _10766_/B _10766_/C vssd1 vssd1 vccd1 vccd1 _11725_/A sky130_fd_sc_hd__nand3b_4
XFILLER_160_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _12659_/A _13194_/D vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__nand2_2
X_16273_ _16273_/A _16273_/B vssd1 vssd1 vccd1 vccd1 _16276_/A sky130_fd_sc_hd__xnor2_1
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13485_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13486_/C sky130_fd_sc_hd__nand2_2
X_10697_ _10694_/X _10697_/B vssd1 vssd1 vccd1 vccd1 _11036_/B sky130_fd_sc_hd__and2b_2
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15224_ _15222_/A _15222_/B _15225_/B vssd1 vssd1 vccd1 vccd1 _15296_/A sky130_fd_sc_hd__a21o_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12436_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__a21o_4
XFILLER_172_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15157_/B sky130_fd_sc_hd__xor2_4
X_12367_ _12198_/A _12367_/B vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__and2b_4
XFILLER_181_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14106_ _13974_/A _13974_/B _14015_/X vssd1 vssd1 vccd1 vccd1 _14108_/B sky130_fd_sc_hd__o21ai_2
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ _11423_/B _11561_/D _11317_/B _11314_/X vssd1 vssd1 vccd1 vccd1 _11320_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_180_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12298_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__nor2_2
XFILLER_99_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15086_ _15726_/A _16226_/C _15085_/B vssd1 vssd1 vccd1 vccd1 _15087_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11249_ _11249_/A _11249_/B _11249_/C vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__or3_1
XFILLER_80_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14037_ _12038_/X _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _14037_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15988_ _15989_/A _15989_/B _15987_/X vssd1 vssd1 vccd1 vccd1 _16096_/B sky130_fd_sc_hd__o21ba_2
XFILLER_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14939_ _17607_/Q _17477_/D _17476_/D _17608_/Q vssd1 vssd1 vccd1 vccd1 _14939_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16609_ _16609_/A _16609_/B _16609_/C vssd1 vssd1 vccd1 vccd1 _16610_/B sky130_fd_sc_hd__and3_1
X_17589_ fanout939/X _17589_/D vssd1 vssd1 vccd1 vccd1 _17589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _09012_/A _09012_/B _09012_/C vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__and3_1
XFILLER_136_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _09914_/A _09914_/B _10029_/A vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__nor3_1
Xfanout602 _15062_/S0 vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__buf_6
Xfanout613 _17153_/A vssd1 vssd1 vccd1 vccd1 _14554_/B sky130_fd_sc_hd__buf_6
Xfanout624 _12597_/B vssd1 vssd1 vccd1 vccd1 _12270_/C sky130_fd_sc_hd__buf_6
Xfanout635 _17506_/Q vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__buf_8
XFILLER_86_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout646 _14593_/D vssd1 vssd1 vccd1 vccd1 _13908_/B sky130_fd_sc_hd__buf_8
X_09845_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__nor2_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout657 _14428_/B vssd1 vssd1 vccd1 vccd1 _16974_/A sky130_fd_sc_hd__buf_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout668 _12576_/D vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__buf_8
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout679 _10180_/B vssd1 vssd1 vccd1 vccd1 _09928_/D sky130_fd_sc_hd__buf_4
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09776_/A _09776_/B _09776_/C vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__and3_1
XFILLER_6_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08727_ _14794_/B vssd1 vssd1 vccd1 vccd1 _08727_/Y sky130_fd_sc_hd__inv_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ _10963_/B _10920_/B _10962_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _10621_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ _10538_/Y _10550_/X _10566_/A _10523_/Y vssd1 vssd1 vccd1 vccd1 _10566_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_139_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10482_ _10709_/A _10370_/B _10481_/X vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__o21a_2
X_13270_ _13271_/A _13271_/B vssd1 vssd1 vccd1 vccd1 _13270_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12221_ _11831_/Y _11835_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _12316_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__a21o_2
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11103_ _11104_/B _11104_/C _11104_/A vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__a21o_4
X_16960_ _17012_/B _16960_/B vssd1 vssd1 vccd1 vccd1 _16960_/X sky130_fd_sc_hd__xor2_1
X_12083_ _12252_/B _12083_/B vssd1 vssd1 vccd1 vccd1 _12085_/C sky130_fd_sc_hd__or2_2
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15911_ _16317_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16813_/B sky130_fd_sc_hd__nand2_8
X_11034_ _11035_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__and2b_2
X_16891_ _16758_/A _16935_/B _16808_/X _16809_/X vssd1 vssd1 vccd1 vccd1 _16893_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _15760_/A _15760_/B _15758_/X vssd1 vssd1 vccd1 vccd1 _15863_/A sky130_fd_sc_hd__o21ai_4
XFILLER_65_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/A _15773_/B vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__nor2_1
XFILLER_18_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ _12985_/A _12985_/B _12985_/C vssd1 vssd1 vccd1 vccd1 _13125_/B sky130_fd_sc_hd__or3_4
XTAP_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ fanout925/X _17512_/D vssd1 vssd1 vccd1 vccd1 _17512_/Q sky130_fd_sc_hd__dfxtp_2
X_14724_ _14750_/A _14726_/C vssd1 vssd1 vccd1 vccd1 _14727_/B sky130_fd_sc_hd__and2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__nor2_4
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17443_ fanout934/X _17443_/D vssd1 vssd1 vccd1 vccd1 _17443_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _14655_/A _14655_/B vssd1 vssd1 vccd1 vccd1 _14656_/B sky130_fd_sc_hd__or2_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11867_/A _11867_/B _11867_/C _11867_/D vssd1 vssd1 vccd1 vccd1 _12093_/A
+ sky130_fd_sc_hd__and4_2
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13606_ _13607_/A _13607_/B _13607_/C vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__o21ai_4
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ _10823_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _10829_/A sky130_fd_sc_hd__nor2_2
X_17374_ input63/X _17396_/A2 _17373_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17515_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14586_ _14629_/C _14587_/B vssd1 vssd1 vccd1 vccd1 _14586_/X sky130_fd_sc_hd__or2_1
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ _14888_/B _11798_/B _11798_/C _11798_/D vssd1 vssd1 vccd1 vccd1 _11800_/C
+ sky130_fd_sc_hd__or4_4
X_16325_ _16667_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16326_/B sky130_fd_sc_hd__nor2_1
X_13537_ _13538_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13537_/Y sky130_fd_sc_hd__nor2_1
XFILLER_158_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10749_ _10750_/B _10750_/C _10750_/A vssd1 vssd1 vccd1 vccd1 _10760_/A sky130_fd_sc_hd__a21o_4
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16256_ _16257_/A _16257_/B vssd1 vssd1 vccd1 vccd1 _16256_/X sky130_fd_sc_hd__and2_1
XFILLER_174_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13468_ _17419_/A _17417_/A _13764_/C _13764_/D vssd1 vssd1 vccd1 vccd1 _13469_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _15262_/C _15208_/C _15208_/D vssd1 vssd1 vccd1 vccd1 _15207_/X sky130_fd_sc_hd__or3_4
XFILLER_127_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12419_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12421_/C sky130_fd_sc_hd__xnor2_4
X_16187_ _16188_/A _16188_/B _16188_/C vssd1 vssd1 vccd1 vccd1 _16187_/Y sky130_fd_sc_hd__o21ai_1
X_13399_ _13398_/C _13526_/A _13397_/Y vssd1 vssd1 vccd1 vccd1 _13401_/B sky130_fd_sc_hd__a21bo_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15138_ _16025_/A _16315_/B vssd1 vssd1 vccd1 vccd1 _15159_/A sky130_fd_sc_hd__nor2_2
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15069_ _15069_/A _15147_/C vssd1 vssd1 vccd1 vccd1 _15069_/X sky130_fd_sc_hd__and2_1
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _09574_/B _09574_/C _09574_/A vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__o21ai_2
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _09779_/A _09654_/D vssd1 vssd1 vccd1 vccd1 _14949_/A sky130_fd_sc_hd__and2_2
XFILLER_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout410 _14775_/A vssd1 vssd1 vccd1 vccd1 _17401_/A sky130_fd_sc_hd__buf_12
Xfanout421 _09030_/A vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__buf_8
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout432 _10241_/B vssd1 vssd1 vccd1 vccd1 _10694_/B sky130_fd_sc_hd__buf_6
XFILLER_150_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout443 _12079_/A vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__buf_6
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout454 _11791_/B vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__buf_12
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout465 _17523_/Q vssd1 vssd1 vccd1 vccd1 _11791_/C sky130_fd_sc_hd__buf_12
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout476 _12595_/A vssd1 vssd1 vccd1 vccd1 _17385_/A sky130_fd_sc_hd__buf_6
X_09828_ _09828_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__xor2_2
Xfanout487 _11240_/A vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__buf_8
XFILLER_98_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout498 _09748_/A vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__buf_2
XFILLER_87_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09759_ _09890_/A _09898_/A _09890_/C vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__o21ai_4
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12770_/A _12770_/B _12923_/D _12770_/D vssd1 vssd1 vccd1 vccd1 _12771_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _10774_/A _10774_/C _10774_/B vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__o21a_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/A _14440_/B _14440_/C vssd1 vssd1 vccd1 vccd1 _14441_/B sky130_fd_sc_hd__nor3_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _14796_/A _11675_/C vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__nor2_2
XFILLER_35_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__xor2_4
X_14371_ _14372_/A _14372_/B _14372_/C vssd1 vssd1 vccd1 vccd1 _14445_/A sky130_fd_sc_hd__o21ai_2
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11583_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16110_ _16107_/Y _16108_/X _16001_/A _16003_/X vssd1 vssd1 vccd1 vccd1 _16111_/C
+ sky130_fd_sc_hd__o211a_1
X_13322_ _13322_/A _13322_/B vssd1 vssd1 vccd1 vccd1 _13324_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ _17090_/A _17093_/B vssd1 vssd1 vccd1 vccd1 _17118_/B sky130_fd_sc_hd__nor2_1
X_10534_ _10535_/A _10533_/Y _10647_/C _10534_/D vssd1 vssd1 vccd1 vccd1 _10644_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_167_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16041_ _16041_/A _16041_/B _16041_/C vssd1 vssd1 vccd1 vccd1 _16043_/A sky130_fd_sc_hd__or3_1
X_10465_ _10465_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10469_/C sky130_fd_sc_hd__xnor2_1
X_13253_ _13249_/Y _13250_/X _13121_/A _13123_/A vssd1 vssd1 vccd1 vccd1 _13253_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ _12371_/A _12202_/Y _11967_/A _11971_/A vssd1 vssd1 vccd1 vccd1 _12206_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_182_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13186_/B sky130_fd_sc_hd__xnor2_1
X_10396_ _10397_/B _10397_/A vssd1 vssd1 vccd1 vccd1 _10396_/X sky130_fd_sc_hd__and2b_1
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ _12135_/A _12135_/B _12442_/B _17139_/A vssd1 vssd1 vccd1 vccd1 _12136_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16943_ _16943_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16944_/B sky130_fd_sc_hd__or2_2
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _17070_/B _12018_/Y _12065_/X vssd1 vssd1 vccd1 vccd1 _17577_/D sky130_fd_sc_hd__o21ai_1
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11017_ _11260_/C _10738_/D _10739_/A _10737_/Y vssd1 vssd1 vccd1 vccd1 _11018_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16874_ _16485_/A _16865_/Y _16873_/X vssd1 vssd1 vccd1 vccd1 _16874_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15825_ _15825_/A _15825_/B vssd1 vssd1 vccd1 vccd1 _15827_/B sky130_fd_sc_hd__xnor2_4
XTAP_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15756_ _15756_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _15759_/A sky130_fd_sc_hd__xnor2_4
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12968_ _12968_/A _12968_/B vssd1 vssd1 vccd1 vccd1 _12971_/A sky130_fd_sc_hd__xnor2_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _14708_/B _14708_/C _14708_/D _14738_/A vssd1 vssd1 vccd1 vccd1 _14713_/A
+ sky130_fd_sc_hd__a22o_1
X_11919_ _11920_/B _12127_/D _11920_/D _12770_/A vssd1 vssd1 vccd1 vccd1 _11921_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15687_ _15687_/A _15687_/B _15686_/Y vssd1 vssd1 vccd1 vccd1 _15782_/B sky130_fd_sc_hd__or3b_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _13049_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _13049_/B sky130_fd_sc_hd__nand3_2
XFILLER_166_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17426_ input60/X _17426_/A2 _17425_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17541_/D
+ sky130_fd_sc_hd__o211a_1
X_14638_ _14638_/A _14638_/B vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ input59/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17357_/X sky130_fd_sc_hd__or3_1
X_14569_ _14569_/A _14569_/B _14569_/C vssd1 vssd1 vccd1 vccd1 _14570_/C sky130_fd_sc_hd__nand3_2
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _16302_/A _17163_/A2 _16307_/X vssd1 vssd1 vccd1 vccd1 _16310_/C sky130_fd_sc_hd__o21ba_1
XFILLER_158_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17288_ _17605_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17288_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16239_ _16239_/A _16239_/B vssd1 vssd1 vccd1 vccd1 _16239_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_146_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08992_ _08994_/A vssd1 vssd1 vccd1 vccd1 _08992_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09613_ _09746_/A _09612_/Y _15537_/A _09928_/D vssd1 vssd1 vccd1 vccd1 _09754_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _09436_/A _09435_/C _09435_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__a21o_1
XFILLER_37_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _09602_/A _09610_/A _09602_/C vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__o21ai_4
XFILLER_180_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10250_ _10243_/B _10245_/B _10243_/A vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__o21ba_4
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _10431_/A _10311_/D _14952_/A vssd1 vssd1 vccd1 vccd1 _10181_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_191_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout240 _14871_/Y vssd1 vssd1 vccd1 vccd1 _16218_/C1 sky130_fd_sc_hd__clkbuf_8
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout251 _15794_/A vssd1 vssd1 vccd1 vccd1 _16207_/B sky130_fd_sc_hd__buf_8
Xfanout262 _15147_/Y vssd1 vssd1 vccd1 vccd1 _15551_/A sky130_fd_sc_hd__buf_6
X_13940_ _14122_/A _13941_/B vssd1 vssd1 vccd1 vccd1 _13940_/X sky130_fd_sc_hd__and2_1
Xfanout273 _15523_/A vssd1 vssd1 vccd1 vccd1 _17063_/A sky130_fd_sc_hd__buf_6
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout284 _15038_/A vssd1 vssd1 vccd1 vccd1 _12390_/S sky130_fd_sc_hd__buf_6
Xfanout295 _17369_/A vssd1 vssd1 vccd1 vccd1 _13838_/S sky130_fd_sc_hd__buf_6
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13871_ _13768_/A _13768_/B _13762_/A vssd1 vssd1 vccd1 vccd1 _13873_/B sky130_fd_sc_hd__a21o_1
XFILLER_189_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15610_ _15610_/A _15610_/B vssd1 vssd1 vccd1 vccd1 _15610_/Y sky130_fd_sc_hd__nor2_4
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12822_ _12823_/B _12822_/B vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__nand2b_4
X_16590_ _16590_/A _16686_/A vssd1 vssd1 vccd1 vccd1 _16591_/C sky130_fd_sc_hd__nor2_1
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15541_ _15541_/A _15541_/B vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__nor2_1
X_12753_ _12907_/A _13300_/C _12754_/A vssd1 vssd1 vccd1 vccd1 _12910_/B sky130_fd_sc_hd__and3_2
XFILLER_188_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11705_/A _11704_/B vssd1 vssd1 vccd1 vccd1 _15889_/A sky130_fd_sc_hd__xnor2_4
X_15472_ _15472_/A _15472_/B vssd1 vssd1 vccd1 vccd1 _15472_/Y sky130_fd_sc_hd__nand2_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12684_ _12685_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__or2_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17547_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17211_/X sky130_fd_sc_hd__and2_1
X_14423_ _14734_/A _14421_/X _14422_/X vssd1 vssd1 vccd1 vccd1 _14423_/Y sky130_fd_sc_hd__a21oi_4
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__xnor2_4
XFILLER_168_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _17167_/A _17163_/A2 _17141_/X vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__o21ba_1
X_14354_ _14416_/B _14354_/B vssd1 vssd1 vccd1 vccd1 _14354_/X sky130_fd_sc_hd__or2_1
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _11566_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__xnor2_1
X_13305_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _13305_/Y sky130_fd_sc_hd__nand2b_1
X_10517_ _10517_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10519_/B sky130_fd_sc_hd__nand2_2
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17073_ _17065_/A _17029_/B _17072_/Y vssd1 vssd1 vccd1 vccd1 _17077_/B sky130_fd_sc_hd__o21a_1
X_14285_ _17070_/B _14283_/X _14352_/B _14211_/X vssd1 vssd1 vccd1 vccd1 _17595_/D
+ sky130_fd_sc_hd__o31ai_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ _11502_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__nand2_2
XFILLER_115_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16024_ _15913_/A _16023_/Y _16022_/X vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__o21ai_4
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13236_ _13236_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _13238_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10448_ _10685_/A _10448_/B vssd1 vssd1 vccd1 vccd1 _10563_/B sky130_fd_sc_hd__nor2_2
XFILLER_170_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13027_/A _13029_/B _13027_/B vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__o21ba_4
X_10379_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__nor2_2
XFILLER_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ _12118_/A _12118_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__nand3_2
XFILLER_123_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13098_ _17419_/A _17417_/A _13551_/D _13434_/D vssd1 vssd1 vccd1 vccd1 _13099_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ _12700_/D _12049_/B vssd1 vssd1 vccd1 vccd1 _12049_/Y sky130_fd_sc_hd__nand2_1
X_16926_ _14080_/C _17075_/A2 _16925_/X vssd1 vssd1 vccd1 vccd1 _16926_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16857_ _16931_/A _16931_/B _16856_/Y vssd1 vssd1 vccd1 vccd1 _16857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15808_ _15808_/A _15808_/B vssd1 vssd1 vccd1 vccd1 _15808_/Y sky130_fd_sc_hd__nor2_1
X_16788_ _14168_/A _16644_/B _16789_/A vssd1 vssd1 vccd1 vccd1 _16788_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ _15740_/A _15740_/B vssd1 vssd1 vccd1 vccd1 _15861_/A sky130_fd_sc_hd__and2b_4
XFILLER_178_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09260_ _09050_/A _09049_/C _09049_/B vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__a21o_1
X_09191_ _11953_/A _11953_/B _12174_/D _12129_/B vssd1 vssd1 vccd1 vccd1 _09196_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17409_ _17409_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17409_/X sky130_fd_sc_hd__or2_1
XFILLER_193_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08975_ _11920_/B _10446_/B _09172_/B _12770_/A vssd1 vssd1 vccd1 vccd1 _08977_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_25_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09527_ _09487_/X _09488_/Y _09507_/Y _09525_/X vssd1 vssd1 vccd1 vccd1 _09530_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09483_/B _09483_/A vssd1 vssd1 vccd1 vccd1 _09458_/X sky130_fd_sc_hd__and2b_1
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _09387_/A _09388_/Y _09343_/X _09344_/Y vssd1 vssd1 vccd1 vccd1 _09393_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _11408_/A _11408_/C _11408_/B vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__o21ai_4
XFILLER_177_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11351_ _11351_/A _11402_/A _11351_/C vssd1 vssd1 vccd1 vccd1 _11354_/A sky130_fd_sc_hd__and3_1
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10302_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10305_/C sky130_fd_sc_hd__nand2_2
X_14070_ _14071_/B _14071_/A vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__and2b_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _11283_/B _11333_/A _11283_/A vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__o21ai_4
XFILLER_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13021_ _13021_/A _13021_/B vssd1 vssd1 vccd1 vccd1 _13024_/A sky130_fd_sc_hd__xnor2_4
X_10233_ _09981_/C _17468_/D _10112_/A _10110_/Y vssd1 vssd1 vccd1 vccd1 _10234_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_3_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10164_ _14786_/A _10971_/A _10647_/D _10745_/D vssd1 vssd1 vccd1 vccd1 _10167_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14972_ _14875_/X _14971_/X _15071_/A vssd1 vssd1 vccd1 vccd1 _14972_/X sky130_fd_sc_hd__a21o_1
X_10095_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__or2_4
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ _16711_/A _16711_/B _16711_/C vssd1 vssd1 vccd1 vccd1 _16712_/B sky130_fd_sc_hd__or3_1
X_13923_ _13923_/A _13923_/B vssd1 vssd1 vccd1 vccd1 _13925_/C sky130_fd_sc_hd__xor2_2
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16642_ _16644_/C _16644_/B _16651_/A vssd1 vssd1 vccd1 vccd1 _16643_/A sky130_fd_sc_hd__a21boi_4
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _13748_/A _13748_/B _13742_/A vssd1 vssd1 vccd1 vccd1 _13856_/B sky130_fd_sc_hd__a21o_1
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12805_ _12805_/A _12805_/B vssd1 vssd1 vccd1 vccd1 _12807_/A sky130_fd_sc_hd__nor2_2
X_16573_ _16481_/A _16482_/Y _16572_/Y vssd1 vssd1 vccd1 vccd1 _16574_/B sky130_fd_sc_hd__a21o_1
X_13785_ _13891_/A _13785_/B vssd1 vssd1 vccd1 vccd1 _13787_/B sky130_fd_sc_hd__nor2_1
XFILLER_62_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ _11164_/B _10996_/B _10996_/C vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__o21ai_1
XFILLER_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15524_ _11624_/Y _15524_/B _15524_/C vssd1 vssd1 vccd1 vccd1 _15525_/B sky130_fd_sc_hd__nand3b_1
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _17387_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _12737_/B sky130_fd_sc_hd__nand2_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15455_ _14805_/A _14805_/B _14805_/C vssd1 vssd1 vccd1 vccd1 _15455_/X sky130_fd_sc_hd__a21o_1
XFILLER_188_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__or2_4
XFILLER_175_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14406_ _14405_/B _14405_/C _14405_/A vssd1 vssd1 vccd1 vccd1 _14406_/Y sky130_fd_sc_hd__a21oi_4
X_11618_ _11617_/B _11616_/Y _11583_/B _11587_/X vssd1 vssd1 vccd1 vccd1 _11624_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_191_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15386_ _15386_/A _15386_/B vssd1 vssd1 vccd1 vccd1 _15386_/Y sky130_fd_sc_hd__nand2_1
X_12598_ _12599_/A _12599_/B vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__nor2_1
XFILLER_184_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17125_ _17125_/A _17125_/B vssd1 vssd1 vccd1 vccd1 _17127_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14337_ _14337_/A _14405_/A _14337_/C vssd1 vssd1 vccd1 vccd1 _14337_/Y sky130_fd_sc_hd__nor3_4
X_11549_ _15888_/A _11549_/B vssd1 vssd1 vccd1 vccd1 _15793_/A sky130_fd_sc_hd__and2_1
XFILLER_183_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17056_ _17057_/B _17056_/B vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__and2b_1
X_14268_ _14268_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14270_/C sky130_fd_sc_hd__xnor2_2
XFILLER_143_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16007_ _16007_/A _16007_/B _16007_/C vssd1 vssd1 vccd1 vccd1 _16007_/X sky130_fd_sc_hd__or3_1
X_13219_ _13220_/A _13220_/B _13220_/C vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__a21o_2
X_14199_ _14200_/A _14200_/B _14198_/X vssd1 vssd1 vccd1 vccd1 _14276_/B sky130_fd_sc_hd__o21ba_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _11027_/A _09892_/D vssd1 vssd1 vccd1 vccd1 _08760_/Y sky130_fd_sc_hd__nand2_8
XFILLER_97_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16909_ _16909_/A _16909_/B vssd1 vssd1 vccd1 vccd1 _16910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09312_ _09261_/A _09261_/B _09310_/B _09401_/A vssd1 vssd1 vccd1 vccd1 _09338_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09243_ _11990_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__nand2_1
XFILLER_193_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _09172_/A _09944_/D _09172_/B _09360_/A vssd1 vssd1 vccd1 vccd1 _09174_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08958_ _08958_/A _09084_/A vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__or2_1
XFILLER_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08889_ _08889_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _09020_/B sky130_fd_sc_hd__xnor2_4
XFILLER_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10920_ _14786_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__and2_4
XTAP_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10851_ _10933_/A _10933_/B _11335_/B _11391_/B vssd1 vssd1 vccd1 vccd1 _10854_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13570_ _13569_/A _13569_/B _13569_/C vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__o21ai_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10782_ _10685_/B _10688_/A _10579_/B _10584_/X vssd1 vssd1 vccd1 vccd1 _11768_/B
+ sky130_fd_sc_hd__a211oi_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ _12521_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12522_/C sky130_fd_sc_hd__xor2_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15241_/A _15241_/B _15241_/C vssd1 vssd1 vccd1 vccd1 _15242_/B sky130_fd_sc_hd__a21o_1
X_12452_ _12452_/A _12452_/B vssd1 vssd1 vccd1 vccd1 _12454_/C sky130_fd_sc_hd__xnor2_2
XFILLER_138_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _11403_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11406_/B sky130_fd_sc_hd__and2_2
XFILLER_172_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15171_ _15171_/A _15171_/B vssd1 vssd1 vccd1 vccd1 _15171_/Y sky130_fd_sc_hd__xnor2_1
X_12383_ _12046_/Y _12049_/Y _12383_/S vssd1 vssd1 vccd1 vccd1 _12383_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _14122_/A _14122_/B vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__nor2_1
XFILLER_181_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11334_ _11480_/A _11437_/B _11334_/C _14897_/A vssd1 vssd1 vccd1 vccd1 _11337_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ _14054_/A _14054_/B vssd1 vssd1 vccd1 vccd1 _14158_/B sky130_fd_sc_hd__nor2_2
X_11265_ _11266_/A _11561_/C vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__and2_4
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13004_ _13004_/A _13004_/B vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__nor2_1
XFILLER_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10216_ _10216_/A _10216_/B _10216_/C vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__and3_2
X_11196_ _11088_/A _11087_/B _11087_/A vssd1 vssd1 vccd1 vccd1 _11198_/B sky130_fd_sc_hd__o21ba_2
XFILLER_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _10148_/B _10148_/C _10148_/A vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__o21a_2
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14955_ _14958_/A _14952_/Y _14954_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14955_/X
+ sky130_fd_sc_hd__a211o_1
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__xor2_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _13906_/A _13906_/B _13906_/C vssd1 vssd1 vccd1 vccd1 _13907_/B sky130_fd_sc_hd__and3_1
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14886_ _15373_/C _15305_/C _14924_/A _14886_/D vssd1 vssd1 vccd1 vccd1 _14886_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16625_ _16625_/A _16625_/B _16623_/X vssd1 vssd1 vccd1 vccd1 _16626_/B sky130_fd_sc_hd__or3b_4
XFILLER_63_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13837_ _13837_/A _17164_/B _13837_/C vssd1 vssd1 vccd1 vccd1 _14841_/B sky130_fd_sc_hd__or3_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16556_ _16638_/A vssd1 vssd1 vccd1 vccd1 _16558_/B sky130_fd_sc_hd__inv_2
X_13768_ _13768_/A _13768_/B vssd1 vssd1 vccd1 vccd1 _13770_/C sky130_fd_sc_hd__xor2_4
X_15507_ _15507_/A _15507_/B vssd1 vssd1 vccd1 vccd1 _15510_/A sky130_fd_sc_hd__xnor2_4
X_12719_ _12720_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__and2_2
X_16487_ _16480_/A _16400_/B _16652_/A vssd1 vssd1 vccd1 vccd1 _16487_/Y sky130_fd_sc_hd__a21oi_1
X_13699_ _14248_/A _16859_/A _13698_/C vssd1 vssd1 vccd1 vccd1 _13700_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15438_ _15439_/A _15439_/B vssd1 vssd1 vccd1 vccd1 _15520_/B sky130_fd_sc_hd__and2b_1
XFILLER_129_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _15369_/A _15369_/B vssd1 vssd1 vccd1 vccd1 _15369_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17108_ _17065_/A _17029_/B _14867_/A vssd1 vssd1 vccd1 vccd1 _17109_/C sky130_fd_sc_hd__a21oi_1
XFILLER_171_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17039_ _17038_/C _17040_/B _17040_/A vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__o21a_1
X_09930_ _09930_/A _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__or3_4
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout806 _15617_/A vssd1 vssd1 vccd1 vccd1 _11334_/C sky130_fd_sc_hd__buf_6
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _09862_/B _09862_/A vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__nand2b_1
Xfanout817 _17487_/Q vssd1 vssd1 vccd1 vccd1 _12502_/B1 sky130_fd_sc_hd__buf_12
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout828 _12618_/D vssd1 vssd1 vccd1 vccd1 _12174_/D sky130_fd_sc_hd__buf_8
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_975 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout839 _17484_/Q vssd1 vssd1 vccd1 vccd1 _12463_/D sky130_fd_sc_hd__clkbuf_16
X_08812_ _08812_/A _08812_/B vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__nor2_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _10067_/A _12129_/B _09643_/C vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__a21oi_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _14836_/A _14872_/A vssd1 vssd1 vccd1 vccd1 _08743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09226_ _09227_/A _09227_/B _09227_/C vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__a21oi_4
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09157_ _12546_/B _12597_/B _09101_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _09165_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_148_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09088_ _09088_/A _09088_/B vssd1 vssd1 vccd1 vccd1 _09317_/C sky130_fd_sc_hd__xnor2_1
XFILLER_123_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11050_ _11051_/A _11051_/B _11051_/C vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__and3_2
XFILLER_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10001_ _10123_/A _10000_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__o21ba_2
XFILLER_190_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _17151_/A _14739_/Y _14737_/X vssd1 vssd1 vccd1 vccd1 _14742_/B sky130_fd_sc_hd__o21a_1
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _11953_/B _12340_/B _12338_/C _11953_/A vssd1 vssd1 vccd1 vccd1 _11956_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _11005_/A _11370_/D vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__nand2_1
XFILLER_189_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _14660_/B _14662_/A _14670_/X vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__a21o_1
XFILLER_45_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _12258_/A _12565_/C vssd1 vssd1 vccd1 vccd1 _11884_/B sky130_fd_sc_hd__nand2_4
X_16410_ _16410_/A _16938_/D _16504_/B vssd1 vssd1 vccd1 vccd1 _16505_/B sky130_fd_sc_hd__or3_1
XFILLER_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13622_ _14756_/A1 _13620_/Y _13621_/X _13517_/Y _13520_/X vssd1 vssd1 vccd1 vccd1
+ _17588_/D sky130_fd_sc_hd__a32o_1
XFILLER_189_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10834_ _10933_/B _10970_/B _11335_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _10834_/Y
+ sky130_fd_sc_hd__a22oi_2
X_17390_ input40/X _17396_/A2 _17389_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17523_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16341_ _16342_/A _16342_/B vssd1 vssd1 vccd1 vccd1 _16444_/B sky130_fd_sc_hd__and2b_1
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _14215_/A _13764_/D vssd1 vssd1 vccd1 vccd1 _13555_/B sky130_fd_sc_hd__nand2_1
XFILLER_160_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10765_ _10631_/X _10693_/Y _10712_/X _10730_/Y vssd1 vssd1 vccd1 vccd1 _10766_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12504_ _12504_/A _12504_/B vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__nor2_1
X_16272_ _16272_/A _16272_/B vssd1 vssd1 vccd1 vccd1 _16273_/B sky130_fd_sc_hd__xnor2_2
XFILLER_157_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13484_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13603_/B sky130_fd_sc_hd__or2_4
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10696_ _10694_/B _11027_/C _11027_/D _10694_/A vssd1 vssd1 vccd1 vccd1 _10697_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15223_ _15774_/A _15647_/A vssd1 vssd1 vccd1 vccd1 _15225_/B sky130_fd_sc_hd__nand2_4
XFILLER_172_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _12435_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _12437_/C sky130_fd_sc_hd__nand2_2
XFILLER_185_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15154_ _15155_/A _15155_/B vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__or2_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12366_ _12366_/A _12366_/B vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__or2_4
X_14105_ _14192_/B _14105_/B vssd1 vssd1 vccd1 vccd1 _14108_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _11314_/X _11317_/B vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__and2b_2
X_15085_ _15913_/A _15085_/B vssd1 vssd1 vccd1 vccd1 _15161_/A sky130_fd_sc_hd__nand2b_1
XFILLER_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12297_ _12620_/A _12618_/D vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__nand2_1
XFILLER_141_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14036_ _12057_/X _12063_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _14036_/X sky130_fd_sc_hd__mux2_4
XFILLER_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11248_ _11249_/B _11249_/C _11249_/A vssd1 vssd1 vccd1 vccd1 _11255_/B sky130_fd_sc_hd__o21ai_4
XFILLER_171_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11179_ _11175_/Y _11176_/X _11015_/X _11019_/X vssd1 vssd1 vccd1 vccd1 _11182_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15987_ _15987_/A _15987_/B vssd1 vssd1 vccd1 vccd1 _15987_/X sky130_fd_sc_hd__xor2_1
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14938_ _17607_/Q _14938_/B vssd1 vssd1 vccd1 vccd1 _14938_/X sky130_fd_sc_hd__or2_2
XFILLER_180_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14869_ _12442_/B _15248_/C _17140_/B _14838_/X _14842_/X vssd1 vssd1 vccd1 vccd1
+ _14869_/X sky130_fd_sc_hd__a311o_1
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _16609_/A _16609_/B _16609_/C vssd1 vssd1 vccd1 vccd1 _16697_/A sky130_fd_sc_hd__a21oi_2
X_17588_ fanout939/X _17588_/D vssd1 vssd1 vccd1 vccd1 _17588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16539_ _16541_/A _16541_/B vssd1 vssd1 vccd1 vccd1 _16627_/A sky130_fd_sc_hd__nand2_4
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09011_ _09012_/A _09012_/B _09012_/C vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__a21oi_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09913_ _09913_/A _09913_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__nand2_2
Xfanout603 _17510_/Q vssd1 vssd1 vccd1 vccd1 _15062_/S0 sky130_fd_sc_hd__buf_6
Xfanout614 _08969_/B vssd1 vssd1 vccd1 vccd1 _17153_/A sky130_fd_sc_hd__buf_6
Xfanout625 _08968_/B vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__buf_8
Xfanout636 _14089_/B vssd1 vssd1 vccd1 vccd1 _13844_/D sky130_fd_sc_hd__buf_6
XFILLER_99_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout647 _17028_/A vssd1 vssd1 vccd1 vccd1 _14545_/C sky130_fd_sc_hd__buf_8
X_09844_ _10241_/B _10377_/B _10491_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _09845_/B
+ sky130_fd_sc_hd__a22oi_4
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout658 _17504_/Q vssd1 vssd1 vccd1 vccd1 _14428_/B sky130_fd_sc_hd__buf_12
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout669 fanout676/X vssd1 vssd1 vccd1 vccd1 _12576_/D sky130_fd_sc_hd__buf_8
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09775_ _09776_/A _09776_/B _09776_/C vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__a21oi_4
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08726_ _15401_/A vssd1 vssd1 vccd1 vccd1 _15274_/A sky130_fd_sc_hd__clkinv_4
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10550_ _10550_/A _10550_/B _10550_/C vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__and3_4
XFILLER_168_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _12166_/A _09509_/B _09209_/C vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__and3_2
X_10481_ _10235_/A _17467_/D _11027_/D _10366_/A vssd1 vssd1 vccd1 vccd1 _10481_/X
+ sky130_fd_sc_hd__a22o_1
X_12220_ _11826_/Y _11829_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ _12316_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__nand3_4
XFILLER_29_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11102_ _11238_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11104_/C sky130_fd_sc_hd__nand2_1
XFILLER_190_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12082_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ _16317_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16129_/B sky130_fd_sc_hd__and2_2
X_11033_ _11005_/A _11005_/B _11007_/X _11006_/X _10957_/D vssd1 vssd1 vccd1 vccd1
+ _11035_/B sky130_fd_sc_hd__a32o_4
X_16890_ _16890_/A _16952_/A vssd1 vssd1 vccd1 vccd1 _16895_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ _15841_/A _15841_/B vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__xnor2_1
XTAP_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ _15772_/A _15772_/B _15772_/C vssd1 vssd1 vccd1 vccd1 _15773_/B sky130_fd_sc_hd__and3_1
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12984_ _12984_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _12985_/C sky130_fd_sc_hd__nand2_2
XTAP_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ fanout925/X _17511_/D vssd1 vssd1 vccd1 vccd1 _17511_/Q sky130_fd_sc_hd__dfxtp_1
X_14723_ _14723_/A _14723_/B _14723_/C vssd1 vssd1 vccd1 vccd1 _14726_/C sky130_fd_sc_hd__or3_1
X_11935_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__nor2_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14655_/A _14655_/B vssd1 vssd1 vccd1 vccd1 _14691_/A sky130_fd_sc_hd__nand2_1
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17442_ fanout934/X _17442_/D vssd1 vssd1 vccd1 vccd1 _17442_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11866_ _11867_/B _11867_/C _11867_/D _12243_/A vssd1 vssd1 vccd1 vccd1 _11868_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13605_/A _13605_/B vssd1 vssd1 vccd1 vccd1 _13607_/C sky130_fd_sc_hd__xor2_4
X_10817_ _10962_/A _11005_/B _10812_/A _10810_/Y vssd1 vssd1 vccd1 vccd1 _10823_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14585_ _14585_/A _14585_/B vssd1 vssd1 vccd1 vccd1 _14587_/B sky130_fd_sc_hd__nand2_1
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17373_ _17373_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17373_/X sky130_fd_sc_hd__or2_1
X_11797_ _14832_/A _17134_/A _17421_/A _14765_/A vssd1 vssd1 vccd1 vccd1 _11798_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13536_ _13403_/B _13409_/B _13403_/A vssd1 vssd1 vccd1 vccd1 _13538_/B sky130_fd_sc_hd__a21boi_4
X_16324_ _16324_/A _16324_/B vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__nand2_1
X_10748_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _10750_/C sky130_fd_sc_hd__nand2_1
XFILLER_174_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16255_ _16158_/A _16158_/B _16145_/Y vssd1 vssd1 vccd1 vccd1 _16257_/B sky130_fd_sc_hd__a21bo_1
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ _14766_/A _13764_/C _13764_/D _14765_/A vssd1 vssd1 vccd1 vccd1 _13469_/A
+ sky130_fd_sc_hd__a22oi_2
X_10679_ _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__and2_2
XFILLER_185_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15206_ _15206_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15206_/X sky130_fd_sc_hd__and2_1
XFILLER_173_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12418_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__and2_1
X_16186_ _16188_/A _16188_/B _16188_/C vssd1 vssd1 vccd1 vccd1 _16189_/A sky130_fd_sc_hd__o21a_1
X_13398_ _13397_/Y _13526_/A _13398_/C vssd1 vssd1 vccd1 vccd1 _13526_/B sky130_fd_sc_hd__nand3b_2
XFILLER_12_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15137_ _11629_/C _14944_/A _15133_/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17546_/D
+ sky130_fd_sc_hd__a22oi_1
XFILLER_126_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _12349_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ _15274_/A _16977_/A _15065_/Y _15067_/X vssd1 vssd1 vccd1 vccd1 _17545_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14019_ _14113_/A _14019_/B vssd1 vssd1 vccd1 vccd1 _14021_/B sky130_fd_sc_hd__and2_1
XFILLER_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09560_ _09689_/A _09689_/B vssd1 vssd1 vccd1 vccd1 _09574_/C sky130_fd_sc_hd__and2_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09491_ _09491_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout400 _13948_/A vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__buf_6
XFILLER_28_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout411 _17529_/Q vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__buf_12
Xfanout422 _11867_/A vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__buf_12
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout433 _11027_/A vssd1 vssd1 vccd1 vccd1 _10241_/B sky130_fd_sc_hd__buf_6
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout444 _12079_/A vssd1 vssd1 vccd1 vccd1 _16108_/C sky130_fd_sc_hd__buf_6
Xfanout455 _11791_/B vssd1 vssd1 vccd1 vccd1 _16317_/A sky130_fd_sc_hd__buf_8
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout466 _17387_/A vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__buf_12
XFILLER_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__xnor2_4
Xfanout477 _17521_/Q vssd1 vssd1 vccd1 vccd1 _12595_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout488 _15262_/B vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__buf_6
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout499 _12592_/A vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__buf_8
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09758_ _09758_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09890_/C sky130_fd_sc_hd__xnor2_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _09689_/A _09689_/B vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__xnor2_2
XFILLER_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__or2_4
XFILLER_27_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ _11651_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _11675_/C sky130_fd_sc_hd__nand2_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10602_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14370_ _14370_/A _14370_/B vssd1 vssd1 vccd1 vccd1 _14372_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11582_ _11582_/A _11583_/A _11582_/C vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__nand3_4
XFILLER_156_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13321_ _17425_/A _17423_/A _13434_/D _13321_/D vssd1 vssd1 vccd1 vccd1 _13322_/B
+ sky130_fd_sc_hd__and4_1
X_10533_ _10171_/B _10647_/D _10645_/C _14789_/A vssd1 vssd1 vccd1 vccd1 _10533_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _16040_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _16041_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13252_ _13252_/A vssd1 vssd1 vccd1 vccd1 _13252_/Y sky130_fd_sc_hd__inv_2
X_10464_ _10465_/B _10465_/A vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__and2b_1
XFILLER_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12203_ _11967_/A _11971_/A _12371_/A _12202_/Y vssd1 vssd1 vccd1 vccd1 _12371_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13183_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13326_/A sky130_fd_sc_hd__and2_1
X_10395_ _10395_/A _10505_/A vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__nor2_4
XFILLER_135_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12134_ _14421_/S _12442_/B _17134_/B _11849_/A vssd1 vssd1 vccd1 vccd1 _12136_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16942_ _16943_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16994_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12065_ _11849_/A _12058_/X _12064_/X _13625_/B vssd1 vssd1 vccd1 vccd1 _12065_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_42_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11016_ _11016_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__xnor2_4
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16873_ _11766_/X _16389_/A _16866_/Y _16872_/X vssd1 vssd1 vccd1 vccd1 _16873_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15824_ _15825_/A _15825_/B vssd1 vssd1 vccd1 vccd1 _15926_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15755_ _16262_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15756_/B sky130_fd_sc_hd__nor2_4
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12967_ _12968_/A _12968_/B vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__and2b_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11918_ _11914_/X _11916_/A _08874_/A _08873_/X vssd1 vssd1 vccd1 vccd1 _11918_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14706_ _13516_/S _12548_/B _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14706_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15686_ _15686_/A _15686_/B vssd1 vssd1 vccd1 vccd1 _15686_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _13049_/A _12899_/B _12899_/C vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__a21o_1
XFILLER_178_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17425_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17425_/X sky130_fd_sc_hd__or2_1
XFILLER_21_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11849_ _11849_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _11849_/Y sky130_fd_sc_hd__nand2_2
X_14637_ _14637_/A1 _12218_/A _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14637_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14569_/A _14569_/B _14569_/C vssd1 vssd1 vccd1 vccd1 _14621_/A sky130_fd_sc_hd__a21o_2
X_17356_ _13300_/D _17360_/A2 _17355_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17507_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16307_ _16302_/B _16580_/A2 _16733_/B1 _16298_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16307_/X sky130_fd_sc_hd__a221o_1
X_13519_ _14666_/S _13519_/B vssd1 vssd1 vccd1 vccd1 _13519_/Y sky130_fd_sc_hd__nor2_1
X_14499_ _17023_/A _14492_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14500_/B sky130_fd_sc_hd__o21ba_1
X_17287_ _17463_/Q _17293_/A2 _17285_/X _17286_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17463_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16238_ _16238_/A _16238_/B vssd1 vssd1 vccd1 vccd1 _16239_/B sky130_fd_sc_hd__xor2_2
XFILLER_174_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _16695_/A _16589_/B _16814_/B _16352_/A vssd1 vssd1 vccd1 vccd1 _16170_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08991_ _08991_/A _08991_/B vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__xnor2_4
XFILLER_125_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09612_ _12135_/B _14863_/B _10431_/B _12135_/A vssd1 vssd1 vccd1 vccd1 _09612_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09543_ _09543_/A _09543_/B vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09474_ _09478_/B _09474_/B vssd1 vssd1 vccd1 vccd1 _09602_/C sky130_fd_sc_hd__and2_2
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10180_ _10431_/A _10180_/B _10180_/C vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__and3_1
XFILLER_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout230 _14931_/X vssd1 vssd1 vccd1 vccd1 _17163_/A2 sky130_fd_sc_hd__buf_6
Xfanout241 _16806_/A2 vssd1 vssd1 vccd1 vccd1 _17170_/B1 sky130_fd_sc_hd__buf_6
Xfanout252 _11784_/X vssd1 vssd1 vccd1 vccd1 _15794_/A sky130_fd_sc_hd__buf_8
XFILLER_120_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout274 _08733_/Y vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__buf_6
Xfanout285 _12383_/S vssd1 vssd1 vccd1 vccd1 _15038_/A sky130_fd_sc_hd__buf_6
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout296 _15458_/A vssd1 vssd1 vccd1 vccd1 _17369_/A sky130_fd_sc_hd__buf_6
XFILLER_115_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _13870_/A _13870_/B vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__xnor2_2
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _12821_/A _12821_/B vssd1 vssd1 vccd1 vccd1 _12823_/B sky130_fd_sc_hd__or2_1
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15540_ _14356_/S _15537_/X _15539_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15540_/X
+ sky130_fd_sc_hd__a211o_1
X_12752_ _12907_/A _12752_/B vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__nand2_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11703_ _11703_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11704_/B sky130_fd_sc_hd__xor2_4
XFILLER_187_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15471_ _15472_/A _15472_/B vssd1 vssd1 vccd1 vccd1 _16604_/B sky130_fd_sc_hd__and2_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12519_/A _12519_/B _12520_/Y vssd1 vssd1 vccd1 vccd1 _12685_/B sky130_fd_sc_hd__o21a_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _17579_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__a21o_1
X_14422_ _12849_/X _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _14422_/X sky130_fd_sc_hd__o21a_1
X_11634_ _11635_/B _11635_/A vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__nand2b_1
XFILLER_30_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14416_/B _14354_/B vssd1 vssd1 vccd1 vccd1 _14353_/Y sky130_fd_sc_hd__nand2_1
X_17141_ _14829_/X _17162_/A2 _16974_/B _14829_/B _17170_/B1 vssd1 vssd1 vccd1 vccd1
+ _17141_/X sky130_fd_sc_hd__a221o_1
X_11565_ _11565_/A _11565_/B _11566_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__or3_1
XFILLER_155_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ _13304_/A _13304_/B vssd1 vssd1 vccd1 vccd1 _13306_/B sky130_fd_sc_hd__xor2_4
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10516_ _10502_/X _10503_/Y _10510_/X _10514_/X vssd1 vssd1 vccd1 vccd1 _10517_/B
+ sky130_fd_sc_hd__a211o_1
X_17072_ _17065_/A _17029_/B _17140_/A vssd1 vssd1 vccd1 vccd1 _17072_/Y sky130_fd_sc_hd__a21oi_1
X_14284_ _14283_/B _14284_/B vssd1 vssd1 vccd1 vccd1 _14352_/B sky130_fd_sc_hd__and2b_1
XFILLER_144_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11496_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16023_ _16938_/A _17119_/C vssd1 vssd1 vccd1 vccd1 _16023_/Y sky130_fd_sc_hd__nand2_2
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13235_ _13235_/A _13235_/B vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__xor2_1
X_10447_ _10559_/A _17302_/A1 _10446_/C vssd1 vssd1 vccd1 vccd1 _10448_/B sky130_fd_sc_hd__a21oi_1
X_13166_ _13036_/A _13038_/B _13036_/B vssd1 vssd1 vccd1 vccd1 _13176_/A sky130_fd_sc_hd__o21ba_4
X_10378_ _11006_/B _10491_/B _10911_/B _11006_/A vssd1 vssd1 vccd1 vccd1 _10379_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_151_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12117_ _12118_/A _12118_/B _12118_/C vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__a21o_4
X_13097_ _17417_/A _13551_/D _13434_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _13099_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _15811_/A _15709_/A _12060_/S vssd1 vssd1 vccd1 vccd1 _12049_/B sky130_fd_sc_hd__mux2_1
X_16925_ _16918_/B _17162_/A2 _16974_/B _14865_/B _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16925_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16856_ _16931_/A _16931_/B _17131_/A vssd1 vssd1 vccd1 vccd1 _16856_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15807_ _13627_/S _15180_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _15808_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16787_ _16787_/A _16853_/C vssd1 vssd1 vccd1 vccd1 _16787_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13999_ _17409_/A _13897_/B _13898_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _14001_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15738_ _15647_/A _16246_/A _15644_/X _15645_/Y vssd1 vssd1 vccd1 vccd1 _15740_/B
+ sky130_fd_sc_hd__a31o_4
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15669_ _15568_/A _15570_/B _15568_/B vssd1 vssd1 vccd1 vccd1 _15671_/B sky130_fd_sc_hd__a21bo_4
XFILLER_34_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17408_ input50/X _17422_/A2 _17407_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17532_/D
+ sky130_fd_sc_hd__o211a_1
X_09190_ _09190_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09196_/A sky130_fd_sc_hd__nor2_2
XFILLER_92_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17339_ input49/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17339_/X sky130_fd_sc_hd__or3_1
XFILLER_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _09242_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__and2_2
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _09507_/Y _09525_/X _09487_/X _09488_/Y vssd1 vssd1 vccd1 vccd1 _09530_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09455_/A _09455_/B _09543_/B _09437_/X vssd1 vssd1 vccd1 vccd1 _09483_/B
+ sky130_fd_sc_hd__a31oi_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ _09388_/A vssd1 vssd1 vccd1 vccd1 _09388_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11350_ _11291_/B _11288_/C _11288_/A vssd1 vssd1 vccd1 vccd1 _11351_/C sky130_fd_sc_hd__a21o_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10411_/B sky130_fd_sc_hd__xnor2_4
XFILLER_152_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11281_ _11520_/C _11334_/C _11281_/C vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__and3_4
XFILLER_180_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _17401_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13021_/B sky130_fd_sc_hd__nand2_4
XFILLER_193_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10232_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__xnor2_4
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10163_ _10163_/A _10163_/B vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__nand2_2
XFILLER_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14971_ _15147_/C _11789_/X _14877_/Y vssd1 vssd1 vccd1 vccd1 _14971_/X sky130_fd_sc_hd__a21o_1
X_10094_ _10094_/A _10348_/A vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16710_ _16711_/A _16711_/B _16711_/C vssd1 vssd1 vccd1 vccd1 _16786_/A sky130_fd_sc_hd__o21ai_4
X_13922_ _13922_/A _13922_/B vssd1 vssd1 vccd1 vccd1 _13923_/B sky130_fd_sc_hd__nand2_2
XFILLER_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _16641_/A _16641_/B vssd1 vssd1 vccd1 vccd1 _16641_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13853_ _13853_/A _13853_/B vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__xor2_2
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12804_ _17419_/A _17417_/A _13321_/D _13194_/D vssd1 vssd1 vccd1 vccd1 _12805_/B
+ sky130_fd_sc_hd__and4_1
X_16572_ _16572_/A _16572_/B vssd1 vssd1 vccd1 vccd1 _16572_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13784_ _13784_/A _13784_/B vssd1 vssd1 vccd1 vccd1 _13785_/B sky130_fd_sc_hd__and2_1
XFILLER_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10996_ _11164_/B _10996_/B _10996_/C vssd1 vssd1 vccd1 vccd1 _11159_/A sky130_fd_sc_hd__or3_4
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _15523_/A _15523_/B vssd1 vssd1 vccd1 vccd1 _15523_/X sky130_fd_sc_hd__or2_2
XFILLER_187_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12735_ _12735_/A _12735_/B vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__nor2_1
XFILLER_188_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12509_/B _12511_/B _12509_/A vssd1 vssd1 vccd1 vccd1 _12668_/B sky130_fd_sc_hd__o21ba_1
X_15454_ _15454_/A _15454_/B _15532_/B vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__and3_1
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14405_ _14405_/A _14405_/B _14405_/C vssd1 vssd1 vccd1 vccd1 _14424_/B sky130_fd_sc_hd__and3_2
X_11617_ _11617_/A _11617_/B _11617_/C vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__or3_2
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15385_ _12858_/Y _17164_/D _15384_/X _15711_/A vssd1 vssd1 vccd1 vccd1 _15386_/B
+ sky130_fd_sc_hd__o22ai_4
X_12597_ _12907_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _12599_/B sky130_fd_sc_hd__and2_1
X_17124_ _17124_/A _17124_/B vssd1 vssd1 vccd1 vccd1 _17125_/B sky130_fd_sc_hd__or2_1
XFILLER_190_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14336_ _14405_/A _14337_/C _14337_/A vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__o21a_2
X_11548_ _11705_/A _11547_/C _11586_/A vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__a21bo_1
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14267_ _14268_/A _14268_/B vssd1 vssd1 vccd1 vccd1 _14344_/B sky130_fd_sc_hd__and2_1
X_17055_ _17093_/B _17055_/B vssd1 vssd1 vccd1 vccd1 _17057_/B sky130_fd_sc_hd__xor2_1
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11479_ _11479_/A _11479_/B vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__nor2_1
XFILLER_109_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16006_ _17119_/B _16005_/B _16005_/C vssd1 vssd1 vccd1 vccd1 _16007_/C sky130_fd_sc_hd__a21oi_1
X_13218_ _13346_/B _13218_/B vssd1 vssd1 vccd1 vccd1 _13220_/C sky130_fd_sc_hd__nand2_1
XFILLER_174_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14198_ _14276_/A _14198_/B vssd1 vssd1 vccd1 vccd1 _14198_/X sky130_fd_sc_hd__or2_1
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13149_ _13149_/A _13149_/B vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__nor2_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16908_ _16908_/A _16908_/B vssd1 vssd1 vccd1 vccd1 _16909_/B sky130_fd_sc_hd__xnor2_2
XFILLER_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16839_ _16775_/A _16775_/B _16771_/A vssd1 vssd1 vccd1 vccd1 _16841_/B sky130_fd_sc_hd__a21bo_1
XFILLER_93_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09311_ _09311_/A _09316_/B _09311_/C vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__and3_2
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09242_ _09242_/A _09242_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09173_ _09360_/A _09944_/D _09502_/C vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__and3_1
XFILLER_193_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08957_ _11932_/A _17505_/Q _08957_/C _08957_/D vssd1 vssd1 vccd1 vccd1 _09084_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08888_ _16315_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__xnor2_4
XFILLER_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10850_ _10850_/A _10855_/A _10850_/C vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__or3_4
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _10560_/B _09509_/B vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__nand2_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _10682_/Y _10689_/X _10779_/B _10780_/Y vssd1 vssd1 vccd1 vccd1 _10784_/B
+ sky130_fd_sc_hd__o31a_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12521_/B _12521_/A vssd1 vssd1 vccd1 vccd1 _12520_/Y sky130_fd_sc_hd__nand2b_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__xnor2_4
XFILLER_138_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ _11402_/A _11402_/B _11451_/A vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__nor3b_4
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15170_ _15170_/A _15170_/B _15170_/C vssd1 vssd1 vccd1 vccd1 _15171_/B sky130_fd_sc_hd__and3_1
X_12382_ _12042_/Y _12044_/Y _12383_/S vssd1 vssd1 vccd1 vccd1 _12382_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_90 _09654_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14121_ _14032_/A _14029_/Y _14031_/B vssd1 vssd1 vccd1 vccd1 _14121_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ _11333_/A _11333_/B vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__nor2_4
XFILLER_193_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _14215_/A _14052_/B vssd1 vssd1 vccd1 vccd1 _14054_/B sky130_fd_sc_hd__nand2_1
XFILLER_193_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11264_ _11264_/A _11270_/A _11264_/C vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__or3_4
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13003_ _13003_/A _13003_/B vssd1 vssd1 vccd1 vccd1 _13004_/B sky130_fd_sc_hd__or2_1
X_10215_ _10214_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10216_/C sky130_fd_sc_hd__nand2b_1
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11195_ _11195_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11198_/A sky130_fd_sc_hd__xnor2_4
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _10508_/C _10743_/C _10268_/B vssd1 vssd1 vccd1 vccd1 _10148_/C sky130_fd_sc_hd__and3_1
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10077_ _10033_/B _10055_/B _10033_/A vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__o21bai_2
X_14954_ _14958_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _14954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13905_ _13906_/A _13906_/B _13906_/C vssd1 vssd1 vccd1 vccd1 _14027_/A sky130_fd_sc_hd__a21oi_2
XFILLER_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14885_ _15396_/A _14888_/B _14888_/C _14888_/D vssd1 vssd1 vccd1 vccd1 _14886_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16624_ _16625_/A _16625_/B _16623_/X vssd1 vssd1 vccd1 vccd1 _16624_/X sky130_fd_sc_hd__o21ba_2
X_13836_ _14756_/A1 _13829_/Y _13830_/X _13835_/X vssd1 vssd1 vccd1 vccd1 _17590_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16555_ _16557_/A _16557_/B _16557_/C vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__o21a_4
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13767_ _13767_/A _13767_/B vssd1 vssd1 vccd1 vccd1 _13768_/B sky130_fd_sc_hd__xnor2_4
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10979_ _11049_/A _11049_/B _11049_/C vssd1 vssd1 vccd1 vccd1 _11051_/A sky130_fd_sc_hd__o21ai_4
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15506_ _15660_/A _16812_/A _15414_/A _15416_/Y vssd1 vssd1 vccd1 vccd1 _15507_/B
+ sky130_fd_sc_hd__a31o_4
X_12718_ _17401_/A _13450_/D _12557_/X _12869_/C _12235_/C vssd1 vssd1 vccd1 vccd1
+ _12720_/B sky130_fd_sc_hd__a32o_2
XFILLER_188_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16486_ _12560_/A _14775_/X _14816_/X _16485_/Y vssd1 vssd1 vccd1 vccd1 _16493_/B
+ sky130_fd_sc_hd__a31o_1
X_13698_ _14248_/A _16859_/A _13698_/C vssd1 vssd1 vccd1 vccd1 _13800_/B sky130_fd_sc_hd__nand3_2
XFILLER_148_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15437_ _15358_/A _15358_/B _15356_/A vssd1 vssd1 vccd1 vccd1 _15439_/B sky130_fd_sc_hd__o21ai_4
XFILLER_30_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ _12650_/B _12649_/B vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__nand2b_4
XFILLER_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15368_ _15233_/X _15299_/Y _15298_/Y vssd1 vssd1 vccd1 vccd1 _15369_/B sky130_fd_sc_hd__o21bai_2
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17107_ _11775_/Y _17105_/Y _17106_/Y vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__a21o_2
XFILLER_190_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14319_ _14319_/A _14389_/A vssd1 vssd1 vccd1 vccd1 _14321_/C sky130_fd_sc_hd__nor2_1
XFILLER_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15299_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15299_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_171_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17038_ _17081_/A _17038_/B _17038_/C vssd1 vssd1 vccd1 vccd1 _17040_/B sky130_fd_sc_hd__nor3_2
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09860_ _09994_/A _15801_/A _09855_/X vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__o21ba_2
Xfanout807 _10839_/D vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__buf_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout818 _09647_/B vssd1 vssd1 vccd1 vccd1 _12338_/D sky130_fd_sc_hd__buf_8
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout829 _12618_/D vssd1 vssd1 vccd1 vccd1 _09791_/B sky130_fd_sc_hd__buf_4
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _09030_/A _11867_/B _12638_/B _12171_/B vssd1 vssd1 vccd1 vccd1 _08812_/B
+ sky130_fd_sc_hd__and4_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_987 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09791_ _10560_/B _09791_/B vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__nand2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08742_ _17607_/Q _17608_/Q vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__or2_4
XFILLER_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09225_ _09225_/A _09225_/B vssd1 vssd1 vccd1 vccd1 _09227_/C sky130_fd_sc_hd__xor2_4
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09152_/A _09153_/X _09131_/X _09138_/X vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_175_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _09317_/A _09086_/Y _15538_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09323_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__nor2_2
XFILLER_66_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _10106_/B sky130_fd_sc_hd__xnor2_4
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11951_ _09014_/A _09013_/B _09013_/A vssd1 vssd1 vccd1 vccd1 _11993_/A sky130_fd_sc_hd__o21ba_2
XFILLER_83_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10902_ _10995_/B _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10953_/A sky130_fd_sc_hd__or3_4
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _14633_/A _14631_/B _14669_/B _14669_/X vssd1 vssd1 vccd1 vccd1 _14670_/X
+ sky130_fd_sc_hd__a31o_1
X_11882_ _11882_/A _11882_/B vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__nor2_2
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10833_ _11266_/A _11122_/B _10970_/B _10971_/B vssd1 vssd1 vccd1 vccd1 _10836_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _13729_/B _13621_/B vssd1 vssd1 vccd1 vccd1 _13621_/X sky130_fd_sc_hd__or2_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _16444_/A _16340_/B vssd1 vssd1 vccd1 vccd1 _16342_/B sky130_fd_sc_hd__nor2_1
X_13552_ _13552_/A _13680_/A vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__or2_1
XFILLER_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10764_ _10771_/B _10764_/B vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__or2_1
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12503_ _12657_/A _12657_/B _13067_/D _12923_/D vssd1 vssd1 vccd1 vccd1 _12504_/B
+ sky130_fd_sc_hd__and4_1
X_16271_ _16271_/A _16271_/B vssd1 vssd1 vccd1 vccd1 _16272_/B sky130_fd_sc_hd__nor2_1
X_13483_ _13603_/A _13483_/B vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10695_ _11027_/B _10809_/D vssd1 vssd1 vccd1 vccd1 _11036_/A sky130_fd_sc_hd__nand2_2
XFILLER_186_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12434_ _12588_/A _12434_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__nand3_4
X_15222_ _15222_/A _15222_/B vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__nand2_2
XFILLER_185_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15153_ _14881_/X _14889_/X _15932_/A _11841_/A vssd1 vssd1 vccd1 vccd1 _15155_/B
+ sky130_fd_sc_hd__a211o_4
X_12365_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12366_/B sky130_fd_sc_hd__a21oi_4
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ _14104_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14105_/B sky130_fd_sc_hd__or2_1
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11316_ _11423_/A _15402_/A _11370_/C _11314_/A vssd1 vssd1 vccd1 vccd1 _11317_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15084_ _15081_/A _15734_/A _15157_/A _15083_/X vssd1 vssd1 vccd1 vccd1 _15085_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12296_ _12296_/A _12508_/A vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__or2_1
XFILLER_10_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14035_ _14763_/S _14033_/X _14034_/Y _13945_/Y vssd1 vssd1 vccd1 vccd1 _17592_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11247_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11249_/C sky130_fd_sc_hd__and2b_1
XFILLER_113_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11178_ _11015_/X _11019_/X _11175_/Y _11176_/X vssd1 vssd1 vccd1 vccd1 _11178_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10129_ _10255_/A _10736_/C vssd1 vssd1 vccd1 vccd1 _10251_/B sky130_fd_sc_hd__nand2_4
X_15986_ _15987_/A _15987_/B vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__and2b_2
X_14937_ _17607_/Q _14938_/B vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__nor2_2
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14868_ _17139_/A _17139_/B vssd1 vssd1 vccd1 vccd1 _17140_/B sky130_fd_sc_hd__and2_1
X_16607_ _16607_/A _16607_/B vssd1 vssd1 vccd1 vccd1 _16609_/C sky130_fd_sc_hd__xor2_2
XFILLER_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _13820_/A _13820_/B vssd1 vssd1 vccd1 vccd1 _13930_/A sky130_fd_sc_hd__and2b_1
XFILLER_91_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17587_ fanout935/X _17587_/D vssd1 vssd1 vccd1 vccd1 _17587_/Q sky130_fd_sc_hd__dfxtp_1
X_14799_ _14790_/Y _14798_/Y _11321_/X vssd1 vssd1 vccd1 vccd1 _15244_/C sky130_fd_sc_hd__o21ba_1
X_16538_ _16447_/Y _16450_/B _16446_/X vssd1 vssd1 vccd1 vccd1 _16541_/B sky130_fd_sc_hd__o21ai_4
XFILLER_149_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16469_ _16469_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16470_/C sky130_fd_sc_hd__xor2_2
XFILLER_192_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09010_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _09012_/C sky130_fd_sc_hd__nand2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09912_ _09912_/A _09912_/B _09912_/C vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__or3_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout604 _11437_/B vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__buf_6
Xfanout615 _17509_/Q vssd1 vssd1 vccd1 vccd1 _08969_/B sky130_fd_sc_hd__buf_12
Xfanout626 _14175_/B vssd1 vssd1 vccd1 vccd1 _13948_/D sky130_fd_sc_hd__buf_6
Xfanout637 _13169_/D vssd1 vssd1 vccd1 vccd1 _14089_/B sky130_fd_sc_hd__buf_6
X_09843_ _10115_/A _10241_/B _10377_/B _10491_/B vssd1 vssd1 vccd1 vccd1 _09845_/A
+ sky130_fd_sc_hd__and4_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout648 _14593_/D vssd1 vssd1 vccd1 vccd1 _17028_/A sky130_fd_sc_hd__clkbuf_16
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout659 _09654_/D vssd1 vssd1 vccd1 vccd1 _12734_/D sky130_fd_sc_hd__buf_8
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09776_/C sky130_fd_sc_hd__xnor2_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08725_ _15703_/A vssd1 vssd1 vccd1 vccd1 _15206_/A sky130_fd_sc_hd__clkinv_4
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1056 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _09208_/A _09208_/B vssd1 vssd1 vccd1 vccd1 _09209_/C sky130_fd_sc_hd__xnor2_1
XFILLER_6_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10480_ _10480_/A _10480_/B vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__xnor2_4
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09150_/A sky130_fd_sc_hd__nor2_2
XFILLER_135_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12150_ _12150_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _12151_/C sky130_fd_sc_hd__xnor2_4
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _11101_/A _11101_/B vssd1 vssd1 vccd1 vccd1 _11238_/B sky130_fd_sc_hd__xnor2_4
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12081_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12252_/B sky130_fd_sc_hd__and2_2
XFILLER_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11035_/A sky130_fd_sc_hd__xnor2_4
XFILLER_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ _15841_/A _15841_/B vssd1 vssd1 vccd1 vccd1 _15840_/Y sky130_fd_sc_hd__nand2_1
XTAP_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15772_/A _15772_/B _15772_/C vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__a21oi_1
XFILLER_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12983_ _12982_/B _12983_/B vssd1 vssd1 vccd1 vccd1 _12984_/B sky130_fd_sc_hd__nand2b_1
XTAP_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ fanout925/X _17510_/D vssd1 vssd1 vccd1 vccd1 _17510_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _14723_/A _14723_/B _14723_/C vssd1 vssd1 vccd1 vccd1 _14750_/A sky130_fd_sc_hd__o21ai_2
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11934_ _11935_/A _11935_/B vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__and2_2
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ fanout934/X _17441_/D vssd1 vssd1 vccd1 vccd1 _17441_/Q sky130_fd_sc_hd__dfxtp_4
X_14653_ _14693_/B _14653_/B vssd1 vssd1 vccd1 vccd1 _14655_/B sky130_fd_sc_hd__xnor2_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__xor2_2
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13604_/A _13604_/B vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__nor2_4
X_10816_ _10816_/A _10816_/B vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__xnor2_1
X_17372_ input62/X _17377_/B _17371_/Y _17372_/C1 vssd1 vssd1 vccd1 vccd1 _17514_/D
+ sky130_fd_sc_hd__o211a_1
X_14584_ _14584_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14629_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11796_ _14766_/A _17415_/A _14769_/A _14770_/A vssd1 vssd1 vccd1 vccd1 _11798_/C
+ sky130_fd_sc_hd__or4_1
X_16323_ _16410_/A _16595_/A _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16324_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13535_ _13535_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__xnor2_4
X_10747_ _10747_/A _10747_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__xnor2_4
XFILLER_159_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16254_ _16254_/A _16254_/B vssd1 vssd1 vccd1 vccd1 _16257_/A sky130_fd_sc_hd__xor2_4
XFILLER_159_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13466_ _13322_/A _13324_/B _13322_/B vssd1 vssd1 vccd1 vccd1 _13473_/A sky130_fd_sc_hd__o21ba_1
X_10678_ _10678_/A _10678_/B vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__nand2_4
X_15205_ _15205_/A _15205_/B vssd1 vssd1 vccd1 vccd1 _15206_/B sky130_fd_sc_hd__nor2_2
X_12417_ _12417_/A _12417_/B vssd1 vssd1 vccd1 vccd1 _12419_/B sky130_fd_sc_hd__xnor2_4
X_16185_ _16165_/A _16533_/B _16060_/A _16058_/A vssd1 vssd1 vccd1 vccd1 _16188_/C
+ sky130_fd_sc_hd__a31o_1
X_13397_ _13950_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _13397_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15136_ _16012_/S _15104_/X _15135_/Y _15808_/A vssd1 vssd1 vccd1 vccd1 _15136_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_182_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12348_ _12349_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__or2_4
XFILLER_154_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12279_ _12108_/A _12110_/B _12108_/B vssd1 vssd1 vccd1 vccd1 _12281_/B sky130_fd_sc_hd__o21ba_1
X_15067_ _17131_/A _15093_/B _15031_/X _15066_/Y vssd1 vssd1 vccd1 vccd1 _15067_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14018_ _14018_/A _14018_/B _14018_/C vssd1 vssd1 vccd1 vccd1 _14019_/B sky130_fd_sc_hd__nand3_1
XFILLER_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15969_ _15969_/A _15969_/B vssd1 vssd1 vccd1 vccd1 _15970_/B sky130_fd_sc_hd__nor2_1
X_09490_ _09928_/C _11813_/B _09353_/A _09351_/Y vssd1 vssd1 vccd1 vccd1 _09491_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout401 _14774_/A vssd1 vssd1 vccd1 vccd1 _13948_/A sky130_fd_sc_hd__buf_6
Xfanout412 _17528_/Q vssd1 vssd1 vccd1 vccd1 _09023_/B sky130_fd_sc_hd__buf_6
XFILLER_120_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout423 _10115_/A vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__buf_6
XFILLER_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout434 _17526_/Q vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__buf_12
XFILLER_87_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout445 _12079_/A vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__buf_2
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout456 _17524_/Q vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__buf_12
X_09826_ _09826_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _12016_/B sky130_fd_sc_hd__nor2_2
XFILLER_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout467 _12578_/A vssd1 vssd1 vccd1 vccd1 _17387_/A sky130_fd_sc_hd__buf_12
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout478 _11095_/A vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__buf_8
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout489 _17520_/Q vssd1 vssd1 vccd1 vccd1 _15262_/B sky130_fd_sc_hd__buf_8
XFILLER_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09757_ _09890_/A _09756_/Y _15537_/A _14863_/B vssd1 vssd1 vccd1 vccd1 _09898_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09688_ _09721_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11651_/A _14792_/B _15008_/B _14792_/A vssd1 vssd1 vccd1 vccd1 _11650_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10601_ _10601_/A _10601_/B vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__xnor2_4
XFILLER_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _11538_/B _11551_/X _11579_/A _11614_/A vssd1 vssd1 vccd1 vccd1 _11582_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13320_ _17423_/A _13434_/D _13321_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _13322_/A
+ sky130_fd_sc_hd__a22oi_2
X_10532_ _14789_/A _10532_/B _10647_/D _10645_/C vssd1 vssd1 vccd1 vccd1 _10535_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _10463_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__nor2_1
X_13251_ _13121_/A _13123_/A _13249_/Y _13250_/X vssd1 vssd1 vccd1 vccd1 _13252_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12202_ _12367_/B _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13182_ _17385_/A _13947_/B _13182_/C vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__and3_1
X_10394_ _10395_/A _10393_/Y _10508_/C _10933_/D vssd1 vssd1 vccd1 vccd1 _10505_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_124_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12133_ _11932_/A _12592_/C _11933_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _12141_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16941_ _16813_/Y _16986_/A _16940_/X _16994_/A vssd1 vssd1 vccd1 vccd1 _16943_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12064_ _14356_/S _12063_/X _15457_/A vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _11016_/B _11016_/A vssd1 vssd1 vccd1 vccd1 _11015_/X sky130_fd_sc_hd__and2b_4
XFILLER_42_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16872_ _16872_/A _16872_/B _16871_/X vssd1 vssd1 vccd1 vccd1 _16872_/X sky130_fd_sc_hd__or3b_4
XFILLER_77_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15823_ _15821_/X _15823_/B vssd1 vssd1 vccd1 vccd1 _15825_/B sky130_fd_sc_hd__and2b_4
XTAP_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15666_/B _15853_/A _15753_/X vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__a21oi_4
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12966_ _12966_/A _12966_/B vssd1 vssd1 vccd1 vccd1 _12968_/B sky130_fd_sc_hd__xnor2_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14705_ _14734_/A _14705_/B vssd1 vssd1 vccd1 vccd1 _14705_/Y sky130_fd_sc_hd__nand2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ _08874_/A _08873_/X _11914_/X _11916_/A vssd1 vssd1 vccd1 vccd1 _11917_/X
+ sky130_fd_sc_hd__o211a_4
X_15685_ _15686_/B _15685_/B _15587_/B vssd1 vssd1 vccd1 vccd1 _15782_/A sky130_fd_sc_hd__or3b_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12897_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _12899_/C sky130_fd_sc_hd__xnor2_2
X_17424_ input59/X _17426_/A2 _17423_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17540_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14734_/A _14636_/B vssd1 vssd1 vccd1 vccd1 _14636_/Y sky130_fd_sc_hd__nand2_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ _14734_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _11848_/Y sky130_fd_sc_hd__nor2_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17355_ input57/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17355_/X sky130_fd_sc_hd__or3_1
X_14567_ _14567_/A _14567_/B vssd1 vssd1 vccd1 vccd1 _14569_/C sky130_fd_sc_hd__xnor2_2
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11779_ _11778_/A _17138_/A _17138_/B _11777_/Y vssd1 vssd1 vccd1 vccd1 _11781_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16306_ _16652_/A _16399_/B _16306_/C vssd1 vssd1 vccd1 vccd1 _16310_/B sky130_fd_sc_hd__or3_1
XFILLER_158_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13518_ _12544_/X _12547_/X _13838_/S vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__mux2_2
X_17286_ _17572_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17286_/X sky130_fd_sc_hd__and2_1
X_14498_ _14562_/A _14498_/B vssd1 vssd1 vccd1 vccd1 _14501_/B sky130_fd_sc_hd__and2_1
XFILLER_174_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16237_ _16238_/A _16238_/B vssd1 vssd1 vccd1 vccd1 _16339_/B sky130_fd_sc_hd__nand2_1
X_13449_ _14383_/A _13564_/D _13450_/D _16913_/C vssd1 vssd1 vccd1 vccd1 _13451_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_173_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16168_ _16619_/A _16168_/B _16168_/C vssd1 vssd1 vccd1 vccd1 _16170_/A sky130_fd_sc_hd__or3_4
XFILLER_127_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _15119_/A _15119_/B vssd1 vssd1 vccd1 vccd1 _15119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16099_ _15994_/A _15994_/B _16100_/B _15991_/X vssd1 vssd1 vccd1 vccd1 _16099_/X
+ sky130_fd_sc_hd__a211o_1
X_08990_ _12772_/A _12127_/D vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__nand2_4
XFILLER_115_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09611_ _12135_/A _12135_/B _14863_/B _10431_/B vssd1 vssd1 vccd1 vccd1 _09746_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09542_ _09484_/A _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__a21oi_4
XFILLER_37_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09473_ _09473_/A _09591_/A _09473_/C vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__or3_1
XFILLER_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout220 _16020_/B vssd1 vssd1 vccd1 vccd1 _16054_/B sky130_fd_sc_hd__buf_12
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout231 _15804_/A2 vssd1 vssd1 vccd1 vccd1 _17075_/A2 sky130_fd_sc_hd__buf_4
Xfanout242 _14871_/Y vssd1 vssd1 vccd1 vccd1 _16806_/A2 sky130_fd_sc_hd__buf_6
Xfanout253 _16389_/A vssd1 vssd1 vccd1 vccd1 _16922_/A sky130_fd_sc_hd__buf_6
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout264 _15891_/B vssd1 vssd1 vccd1 vccd1 _15796_/B sky130_fd_sc_hd__buf_4
XFILLER_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout275 _16911_/A vssd1 vssd1 vccd1 vccd1 _17131_/A sky130_fd_sc_hd__buf_6
XFILLER_189_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout286 _15056_/A vssd1 vssd1 vccd1 vccd1 _12383_/S sky130_fd_sc_hd__buf_4
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09809_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__nand2_1
Xfanout297 _15458_/A vssd1 vssd1 vccd1 vccd1 _15901_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12820_ _12820_/A _12820_/B _12820_/C vssd1 vssd1 vccd1 vccd1 _12821_/B sky130_fd_sc_hd__and3_1
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ _12751_/A _12910_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__nor2_2
XFILLER_188_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _15793_/A _15793_/B vssd1 vssd1 vccd1 vccd1 _15888_/B sky130_fd_sc_hd__nand2_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15442_/Y _15443_/X _15441_/X vssd1 vssd1 vccd1 vccd1 _15522_/A sky130_fd_sc_hd__a21o_2
XFILLER_188_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12685_/A sky130_fd_sc_hd__xnor2_2
XFILLER_91_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _12847_/B _12852_/X _14421_/S vssd1 vssd1 vccd1 vccd1 _14421_/X sky130_fd_sc_hd__mux2_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11649_/A _11632_/B _11632_/A vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__o21ba_2
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _17140_/A _17140_/B _17140_/C vssd1 vssd1 vccd1 vccd1 _17140_/X sky130_fd_sc_hd__or3_1
X_14352_ _14352_/A _14352_/B vssd1 vssd1 vccd1 vccd1 _14354_/B sky130_fd_sc_hd__or2_1
XFILLER_156_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11564_ _11564_/A _11590_/A vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__nor2_1
XFILLER_183_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13303_ _13303_/A _13303_/B vssd1 vssd1 vccd1 vccd1 _13304_/B sky130_fd_sc_hd__xnor2_4
X_10515_ _10510_/X _10514_/X _10502_/X _10503_/Y vssd1 vssd1 vccd1 vccd1 _10517_/A
+ sky130_fd_sc_hd__o211ai_4
X_17071_ _11773_/A _11773_/B _17070_/Y vssd1 vssd1 vccd1 vccd1 _17077_/A sky130_fd_sc_hd__o21a_2
X_14283_ _14284_/B _14283_/B vssd1 vssd1 vccd1 vccd1 _14283_/X sky130_fd_sc_hd__and2b_1
X_11495_ _11495_/A _11495_/B _11532_/A vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__nor3b_4
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16022_ _16226_/C _16165_/B _17119_/C _15726_/A vssd1 vssd1 vccd1 vccd1 _16022_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10446_ _10559_/A _10446_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10685_/A sky130_fd_sc_hd__and3_2
XFILLER_108_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13234_ _13235_/B _13235_/A vssd1 vssd1 vccd1 vccd1 _13361_/B sky130_fd_sc_hd__and2b_1
XFILLER_164_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ _13165_/A _13165_/B _13165_/C vssd1 vssd1 vccd1 vccd1 _13178_/B sky130_fd_sc_hd__nand3_4
X_10377_ _11005_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__nand2_4
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12116_ _12116_/A _12116_/B vssd1 vssd1 vccd1 vccd1 _12118_/C sky130_fd_sc_hd__or2_2
XFILLER_111_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13096_ _12924_/A _12926_/B _12924_/B vssd1 vssd1 vccd1 vccd1 _13103_/A sky130_fd_sc_hd__o21ba_1
XFILLER_123_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12047_ _12040_/Y _12042_/Y _12044_/Y _12046_/Y _12383_/S _15312_/S vssd1 vssd1 vccd1
+ vccd1 _12047_/X sky130_fd_sc_hd__mux4_2
X_16924_ _14865_/B _16868_/A _16923_/Y vssd1 vssd1 vccd1 vccd1 _16924_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16855_ _16716_/Y _16854_/D _16854_/X _16852_/Y vssd1 vssd1 vccd1 vccd1 _16931_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_66_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15806_ _15458_/A _15179_/X _15806_/B1 vssd1 vssd1 vccd1 vccd1 _15806_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16786_ _16786_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16853_/C sky130_fd_sc_hd__xor2_4
XFILLER_168_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13998_ _13998_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _14001_/A sky130_fd_sc_hd__nor2_2
XFILLER_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15737_ _15737_/A _15737_/B vssd1 vssd1 vccd1 vccd1 _15740_/A sky130_fd_sc_hd__xnor2_4
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12949_ _12949_/A _13092_/A vssd1 vssd1 vccd1 vccd1 _12950_/C sky130_fd_sc_hd__and2_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15668_ _15668_/A _15668_/B vssd1 vssd1 vccd1 vccd1 _15671_/A sky130_fd_sc_hd__xor2_4
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17407_ _17407_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17407_/X sky130_fd_sc_hd__or2_1
X_14619_ _14658_/B _14619_/B vssd1 vssd1 vccd1 vccd1 _14621_/C sky130_fd_sc_hd__or2_1
XFILLER_21_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15599_ _15599_/A _15599_/B vssd1 vssd1 vccd1 vccd1 _15601_/B sky130_fd_sc_hd__nand2_4
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17338_ _13094_/B _17360_/A2 _17337_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17498_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17269_ _17457_/Q _17293_/A2 _17267_/X _17268_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17457_/D sky130_fd_sc_hd__o221a_1
XFILLER_140_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ _08973_/A _08973_/B _09095_/A vssd1 vssd1 vccd1 vccd1 _08974_/B sky130_fd_sc_hd__or3_1
XFILLER_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09525_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__and2_2
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09456_ _09456_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__xnor2_4
XFILLER_40_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09387_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__and3_4
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10300_ _10300_/A _10418_/A vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__or2_4
XFILLER_180_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11280_ _11283_/B _11280_/B vssd1 vssd1 vccd1 vccd1 _11281_/C sky130_fd_sc_hd__nor2_1
XFILLER_119_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10231_ _10134_/A _10134_/C _10134_/B vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10162_ _10162_/A _10170_/A _10162_/C vssd1 vssd1 vccd1 vccd1 _10163_/B sky130_fd_sc_hd__or3_1
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14970_ _14899_/X _14968_/X _08727_/Y vssd1 vssd1 vccd1 vccd1 _16025_/A sky130_fd_sc_hd__a21o_4
X_10093_ _09806_/A _09807_/Y _10094_/A _10092_/X vssd1 vssd1 vccd1 vccd1 _10348_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_94_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13921_ _13921_/A _13921_/B _13921_/C vssd1 vssd1 vccd1 vccd1 _13922_/B sky130_fd_sc_hd__nand3_1
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16640_ _11756_/A _11756_/B _16568_/B _16568_/A vssd1 vssd1 vccd1 vccd1 _16641_/B
+ sky130_fd_sc_hd__a22o_2
X_13852_ _13852_/A _13947_/B _13853_/B vssd1 vssd1 vccd1 vccd1 _13958_/B sky130_fd_sc_hd__and3_1
XFILLER_63_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _17417_/A _13321_/D _13194_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _12805_/A
+ sky130_fd_sc_hd__a22oi_4
X_16571_ _16571_/A _17153_/B _14774_/A vssd1 vssd1 vccd1 vccd1 _16572_/B sky130_fd_sc_hd__or3b_1
XFILLER_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _13784_/A _13784_/B vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__nor2_1
X_10995_ _10995_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _10996_/C sky130_fd_sc_hd__nor2_1
XFILLER_76_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _15522_/A _15522_/B vssd1 vssd1 vccd1 vccd1 _15523_/B sky130_fd_sc_hd__xor2_1
X_12734_ _17391_/A _17389_/A _12734_/C _12734_/D vssd1 vssd1 vccd1 vccd1 _12735_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15532_/A _15453_/B _15453_/C vssd1 vssd1 vccd1 vccd1 _15532_/B sky130_fd_sc_hd__nand3_1
XFILLER_176_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__xor2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ _14399_/X _14466_/B _14296_/X _14337_/Y vssd1 vssd1 vccd1 vccd1 _14405_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_169_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11616_ _11617_/A _11617_/B _11617_/C vssd1 vssd1 vccd1 vccd1 _11616_/Y sky130_fd_sc_hd__nor3_2
X_15384_ _15097_/X _15100_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _15384_/X sky130_fd_sc_hd__mux2_2
X_12596_ _12596_/A _12755_/A vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__nor2_1
X_17123_ _17124_/A _17124_/B vssd1 vssd1 vccd1 vccd1 _17125_/A sky130_fd_sc_hd__nand2_1
X_14335_ _14332_/X _14333_/Y _14239_/A _14256_/X vssd1 vssd1 vccd1 vccd1 _14337_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_129_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11547_ _11586_/A _11705_/A _11547_/C vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__nand3b_2
XFILLER_51_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17054_ _17090_/A _17093_/A vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14266_ _14266_/A _14266_/B vssd1 vssd1 vccd1 vccd1 _14268_/B sky130_fd_sc_hd__xnor2_2
X_11478_ _11520_/C _11480_/C _11440_/A _11438_/Y vssd1 vssd1 vccd1 vccd1 _11479_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16005_ _17119_/B _16005_/B _16005_/C vssd1 vssd1 vccd1 vccd1 _16007_/B sky130_fd_sc_hd__and3_1
XFILLER_171_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13217_ _17407_/A _13564_/D _13216_/C vssd1 vssd1 vccd1 vccd1 _13218_/B sky130_fd_sc_hd__a21o_1
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__nor2_4
X_14197_ _14197_/A _14197_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__and3_1
XFILLER_124_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13148_ _13948_/A _13948_/B _14153_/C _13566_/B vssd1 vssd1 vccd1 vccd1 _13149_/B
+ sky130_fd_sc_hd__and4_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _17411_/A _13866_/D _13229_/B _14769_/A vssd1 vssd1 vccd1 vccd1 _13083_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16907_ _16906_/A _16906_/B _16908_/A vssd1 vssd1 vccd1 vccd1 _17012_/A sky130_fd_sc_hd__a21o_1
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16838_ _16838_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _16841_/A sky130_fd_sc_hd__xnor2_2
XFILLER_93_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16769_ _16770_/A _16770_/B _16770_/C vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__o21ai_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _09310_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _09311_/C sky130_fd_sc_hd__xnor2_1
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _09242_/A _09242_/B _09242_/C vssd1 vssd1 vccd1 vccd1 _11990_/A sky130_fd_sc_hd__a21o_2
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09172_ _09172_/A _09172_/B vssd1 vssd1 vccd1 vccd1 _09502_/C sky130_fd_sc_hd__and2_1
XFILLER_193_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08956_ _11930_/B _09652_/B _11808_/B _12135_/A vssd1 vssd1 vccd1 vccd1 _08957_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08887_ _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08888_/B sky130_fd_sc_hd__nor2_2
XFILLER_57_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__xor2_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _10780_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09439_ _09439_/A _09439_/B vssd1 vssd1 vccd1 vccd1 _09441_/C sky130_fd_sc_hd__or2_2
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12450_ _12451_/B _12451_/A vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__and2b_1
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ _11349_/A _11349_/B _11349_/C vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__a21oi_4
XFILLER_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ _12696_/A _12379_/B _12380_/Y vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__a21o_1
XANTENNA_80 _17459_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_91 _09654_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _14279_/A _14120_/B vssd1 vssd1 vccd1 vccd1 _14278_/A sky130_fd_sc_hd__nand2b_2
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11332_ _11520_/C _11334_/C _11281_/C vssd1 vssd1 vccd1 vccd1 _11333_/B sky130_fd_sc_hd__a21oi_2
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14051_ _14051_/A _14158_/A vssd1 vssd1 vccd1 vccd1 _14054_/A sky130_fd_sc_hd__or2_1
XFILLER_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11263_ _11264_/A _11264_/C vssd1 vssd1 vccd1 vccd1 _11270_/B sky130_fd_sc_hd__nor2_2
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__or2_1
XFILLER_97_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10214_ _10214_/A _10214_/B _10214_/C vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__or3_4
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__nor2_2
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10076_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__nor2_2
X_14953_ _12054_/A _15101_/A1 _10180_/C vssd1 vssd1 vccd1 vccd1 _15038_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13904_ _13904_/A _13904_/B vssd1 vssd1 vccd1 vccd1 _13906_/C sky130_fd_sc_hd__xnor2_2
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14884_ _14888_/B _14888_/C _14888_/D vssd1 vssd1 vccd1 vccd1 _14887_/B sky130_fd_sc_hd__or3_4
XFILLER_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16623_ _16699_/A _16623_/B vssd1 vssd1 vccd1 vccd1 _16623_/X sky130_fd_sc_hd__or2_1
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13835_ _14839_/A _11848_/Y _13834_/Y _13832_/Y _12853_/X vssd1 vssd1 vccd1 vccd1
+ _13835_/X sky130_fd_sc_hd__a32o_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16554_ _16554_/A _16554_/B vssd1 vssd1 vccd1 vccd1 _16557_/C sky130_fd_sc_hd__xnor2_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _14215_/A _13866_/C vssd1 vssd1 vccd1 vccd1 _13767_/B sky130_fd_sc_hd__nand2_4
XFILLER_188_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _11049_/C sky130_fd_sc_hd__xor2_4
X_15505_ _15505_/A _15505_/B vssd1 vssd1 vccd1 vccd1 _15512_/A sky130_fd_sc_hd__xnor2_2
XFILLER_189_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12717_ _12717_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _12720_/A sky130_fd_sc_hd__xnor2_2
X_16485_ _16485_/A _16485_/B vssd1 vssd1 vccd1 vccd1 _16485_/Y sky130_fd_sc_hd__nand2_1
X_13697_ _13697_/A _13800_/A vssd1 vssd1 vccd1 vccd1 _13698_/C sky130_fd_sc_hd__and2_1
X_15436_ _15436_/A _15436_/B vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__xnor2_4
X_12648_ _12795_/A _12638_/B _12496_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12649_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15367_ _15365_/X _15367_/B vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__nand2b_1
X_12579_ _12579_/A _12579_/B vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__xnor2_2
XFILLER_157_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17106_ _11775_/Y _17105_/Y _16922_/A vssd1 vssd1 vccd1 vccd1 _17106_/Y sky130_fd_sc_hd__o21ai_1
X_14318_ _14450_/A _14318_/B _14318_/C _14641_/D vssd1 vssd1 vccd1 vccd1 _14389_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_102_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15298_ _15299_/A _15299_/B vssd1 vssd1 vccd1 vccd1 _15298_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17037_ _17037_/A _17037_/B vssd1 vssd1 vccd1 vccd1 _17056_/B sky130_fd_sc_hd__nor2_1
X_14249_ _14248_/A _14599_/D _14248_/C vssd1 vssd1 vccd1 vccd1 _14250_/B sky130_fd_sc_hd__a21o_1
XFILLER_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout808 _17488_/Q vssd1 vssd1 vccd1 vccd1 _10839_/D sky130_fd_sc_hd__buf_12
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout819 _12770_/D vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_140_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ _11867_/B _12638_/B _12171_/B _09030_/A vssd1 vssd1 vccd1 vccd1 _08812_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09933_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__xnor2_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08741_ _15147_/C _14836_/A _08740_/Y vssd1 vssd1 vccd1 vccd1 _17612_/D sky130_fd_sc_hd__a21o_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _12166_/A _12158_/C vssd1 vssd1 vccd1 vccd1 _09225_/B sky130_fd_sc_hd__nand2_2
XFILLER_179_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09155_ _09155_/A vssd1 vssd1 vccd1 vccd1 _09155_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09086_ _12135_/B _11808_/B _09926_/B _12135_/A vssd1 vssd1 vccd1 vccd1 _09086_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09988_ _09988_/A _09988_/B vssd1 vssd1 vccd1 vccd1 _10106_/A sky130_fd_sc_hd__xnor2_4
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08939_ _11930_/B _12270_/D _12102_/D _17373_/A vssd1 vssd1 vccd1 vccd1 _08941_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_130_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11950_ _11947_/X _11948_/Y _09016_/A _09016_/Y vssd1 vssd1 vccd1 vccd1 _11998_/B
+ sky130_fd_sc_hd__o211a_4
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _10901_/A _10901_/B vssd1 vssd1 vccd1 vccd1 _10902_/C sky130_fd_sc_hd__nor2_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11881_ _12256_/A _12256_/B _12088_/D _11881_/D vssd1 vssd1 vccd1 vccd1 _11882_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13620_ _13729_/B _13621_/B vssd1 vssd1 vccd1 vccd1 _13620_/Y sky130_fd_sc_hd__nand2_1
X_10832_ _10863_/A vssd1 vssd1 vccd1 vccd1 _11075_/A sky130_fd_sc_hd__inv_2
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13551_ _14050_/A _14050_/B _13664_/D _13551_/D vssd1 vssd1 vccd1 vccd1 _13680_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ _10771_/A _10734_/X _10760_/A _10761_/Y vssd1 vssd1 vccd1 vccd1 _10764_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_186_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12502_ _12657_/B _13067_/D _12502_/B1 _12657_/A vssd1 vssd1 vccd1 vccd1 _12504_/A
+ sky130_fd_sc_hd__a22oi_2
X_16270_ _16270_/A _16270_/B _16270_/C vssd1 vssd1 vccd1 vccd1 _16271_/B sky130_fd_sc_hd__nor3_1
XFILLER_185_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13482_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__or2_1
XFILLER_185_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10694_ _10694_/A _10694_/B _11027_/C _11027_/D vssd1 vssd1 vccd1 vccd1 _10694_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15221_ _15221_/A _15221_/B vssd1 vssd1 vccd1 vccd1 _15226_/A sky130_fd_sc_hd__xnor2_4
XFILLER_157_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ _12588_/A _12434_/B _12434_/C vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__a21o_1
XFILLER_185_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ _15551_/A _15152_/B _15175_/B vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__or3b_4
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12364_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__and3_2
XFILLER_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _14104_/A _14104_/B vssd1 vssd1 vccd1 vccd1 _14192_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11315_ _11423_/B _11561_/D vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__nand2_2
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15083_ _15278_/A _15821_/A _15647_/A _15660_/A vssd1 vssd1 vccd1 vccd1 _15083_/X
+ sky130_fd_sc_hd__a22o_1
X_12295_ _12618_/A _12770_/B _12463_/D _12295_/D vssd1 vssd1 vccd1 vccd1 _12508_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ _14122_/B _14034_/B vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11246_ _11246_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__nor2_4
XFILLER_106_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11177_ _11015_/X _11019_/X _11175_/Y _11176_/X vssd1 vssd1 vccd1 vccd1 _11182_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10128_ _10128_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__nor2_2
X_15985_ _15867_/B _15875_/B _15867_/A vssd1 vssd1 vccd1 vccd1 _15987_/B sky130_fd_sc_hd__a21bo_1
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10059_ _10059_/A _10059_/B _10059_/C vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__nor3_4
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14936_ _14942_/A _10560_/D _15248_/C _15899_/A2 _14935_/X vssd1 vssd1 vccd1 vccd1
+ _14944_/B sky130_fd_sc_hd__o32a_1
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ _14867_/A _17065_/A _17029_/B vssd1 vssd1 vccd1 vccd1 _17139_/B sky130_fd_sc_hd__and3_1
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16606_ _16807_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16607_/B sky130_fd_sc_hd__nand2_1
X_13818_ _13818_/A _13818_/B vssd1 vssd1 vccd1 vccd1 _13820_/B sky130_fd_sc_hd__nand2_2
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17586_ fanout936/X _17586_/D vssd1 vssd1 vccd1 vccd1 _17586_/Q sky130_fd_sc_hd__dfxtp_1
X_14798_ _14791_/X _14797_/X _11469_/X vssd1 vssd1 vccd1 vccd1 _14798_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_189_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16537_ _16537_/A _16537_/B vssd1 vssd1 vccd1 vccd1 _16541_/A sky130_fd_sc_hd__xnor2_4
X_13749_ _13749_/A _13749_/B vssd1 vssd1 vccd1 vccd1 _13751_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16468_ _16469_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16558_/A sky130_fd_sc_hd__and2b_2
XFILLER_176_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15419_ _15419_/A _15419_/B vssd1 vssd1 vccd1 vccd1 _15422_/A sky130_fd_sc_hd__xor2_4
XFILLER_191_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16399_ _16399_/A _16399_/B vssd1 vssd1 vccd1 vccd1 _16400_/C sky130_fd_sc_hd__nor2_1
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09911_ _09912_/A _09912_/B _09912_/C vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout605 _11437_/B vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__buf_6
Xfanout616 _17139_/A vssd1 vssd1 vccd1 vccd1 _12752_/B sky130_fd_sc_hd__clkbuf_16
Xfanout627 _13300_/D vssd1 vssd1 vccd1 vccd1 _14175_/B sky130_fd_sc_hd__clkbuf_8
X_09842_ _09842_/A _09842_/B _09848_/B vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__or3_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout638 _17506_/Q vssd1 vssd1 vccd1 vccd1 _13169_/D sky130_fd_sc_hd__buf_6
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout649 _17505_/Q vssd1 vssd1 vccd1 vccd1 _14593_/D sky130_fd_sc_hd__clkbuf_16
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B _09773_/C vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__or3_2
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _17139_/A vssd1 vssd1 vccd1 vccd1 _17134_/B sky130_fd_sc_hd__inv_2
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09207_ _09208_/B _09208_/A vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__and2b_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09138_ _09170_/B _09170_/A vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__and2b_1
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09069_ _09069_/A _09076_/B vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__nand2_2
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11238_/A sky130_fd_sc_hd__xnor2_4
X_12080_ _12080_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__xnor2_1
XFILLER_104_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _11032_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11176_/A sky130_fd_sc_hd__and2_2
XFILLER_104_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15770_ _15662_/A _15774_/B _15663_/A _15660_/X vssd1 vssd1 vccd1 vccd1 _15772_/C
+ sky130_fd_sc_hd__a31oi_4
XTAP_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12983_/B _12982_/B vssd1 vssd1 vccd1 vccd1 _12984_/A sky130_fd_sc_hd__nand2b_4
XTAP_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14747_/B _14721_/B vssd1 vssd1 vccd1 vccd1 _14723_/C sky130_fd_sc_hd__and2_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _11933_/A _11933_/B vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ fanout934/X _17440_/D vssd1 vssd1 vccd1 vccd1 _17440_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14683_/A _14693_/A vssd1 vssd1 vccd1 vccd1 _14653_/B sky130_fd_sc_hd__nor2_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13603_/A _13603_/B _13603_/C vssd1 vssd1 vccd1 vccd1 _13604_/B sky130_fd_sc_hd__and3_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10816_/A _10816_/B vssd1 vssd1 vccd1 vccd1 _11057_/B sky130_fd_sc_hd__nand2_2
X_17371_ _17371_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17371_/Y sky130_fd_sc_hd__nand2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _14583_/A _14583_/B _14583_/C vssd1 vssd1 vccd1 vccd1 _14584_/B sky130_fd_sc_hd__and3_1
X_11795_ _14775_/A _14776_/A _14777_/A _16209_/C vssd1 vssd1 vccd1 vccd1 _11799_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_158_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16322_ _16505_/A _16743_/C _17043_/B _15209_/Y vssd1 vssd1 vccd1 vccd1 _16324_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13534_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__xnor2_4
XFILLER_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ _10746_/A _10984_/A vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__or2_2
XFILLER_186_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16253_ _16254_/A _16254_/B vssd1 vssd1 vccd1 vccd1 _16347_/B sky130_fd_sc_hd__nor2_1
XFILLER_185_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13465_ _13465_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__xor2_2
X_10677_ _10678_/A _10677_/B _10677_/C vssd1 vssd1 vccd1 vccd1 _10678_/B sky130_fd_sc_hd__nand3_4
XFILLER_185_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15204_ _15204_/A _16880_/A _15270_/A vssd1 vssd1 vccd1 vccd1 _15205_/B sky130_fd_sc_hd__or3b_4
X_12416_ _17393_/A _12565_/C vssd1 vssd1 vccd1 vccd1 _12417_/B sky130_fd_sc_hd__nand2_4
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16184_ _16184_/A _16184_/B vssd1 vssd1 vccd1 vccd1 _16192_/A sky130_fd_sc_hd__nor2_2
X_13396_ _13844_/A _13844_/B _13523_/B _13895_/C vssd1 vssd1 vccd1 vccd1 _13526_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15135_ _15711_/A _15711_/B _15134_/X vssd1 vssd1 vccd1 vccd1 _15135_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_153_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12347_ _12180_/B _12182_/B _12180_/A vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__o21ba_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15066_ _17164_/C _15064_/X _15055_/X vssd1 vssd1 vccd1 vccd1 _15066_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_114_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12278_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12281_/A sky130_fd_sc_hd__xnor2_2
X_14017_ _14018_/A _14018_/B _14018_/C vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _11229_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11229_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15968_ _15969_/A _15969_/B vssd1 vssd1 vccd1 vccd1 _16084_/B sky130_fd_sc_hd__and2_1
XFILLER_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14919_ _14916_/X _14918_/Y _15130_/S vssd1 vssd1 vccd1 vccd1 _14919_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15899_ _15895_/B _15899_/A2 _16008_/B1 _15898_/A _16008_/C1 vssd1 vssd1 vccd1 vccd1
+ _15899_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17569_ fanout945/X _17569_/D vssd1 vssd1 vccd1 vccd1 _17569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 _14774_/A vssd1 vssd1 vccd1 vccd1 _17403_/A sky130_fd_sc_hd__buf_8
XFILLER_63_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout413 _17528_/Q vssd1 vssd1 vccd1 vccd1 _12068_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout424 _11867_/A vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__buf_6
XFILLER_98_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout435 _13405_/B vssd1 vssd1 vccd1 vccd1 _17395_/A sky130_fd_sc_hd__buf_8
XFILLER_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout446 _17525_/Q vssd1 vssd1 vccd1 vccd1 _12079_/A sky130_fd_sc_hd__buf_12
X_09825_ _09825_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__and2_1
Xfanout457 _12256_/B vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__buf_8
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout468 _10904_/B vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__buf_12
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout479 _10392_/A vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__buf_6
XFILLER_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ _10171_/B _10431_/B _10543_/B _14789_/A vssd1 vssd1 vccd1 vccd1 _09756_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09576_/A _09575_/C _09575_/B vssd1 vssd1 vccd1 vccd1 _09721_/B sky130_fd_sc_hd__a21o_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10600_ _11027_/B _17469_/D _10593_/A _10592_/A vssd1 vssd1 vccd1 vccd1 _10603_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_167_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11580_ _11579_/A _11614_/A _11538_/B _11551_/X vssd1 vssd1 vccd1 vccd1 _11583_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_167_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10531_ _10531_/A _10536_/A _10531_/C vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__or3_4
XFILLER_168_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13250_ _13249_/A _13249_/B _13249_/C _13249_/D vssd1 vssd1 vccd1 vccd1 _13250_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10462_ _10454_/A _10455_/X _10463_/A _10461_/X vssd1 vssd1 vccd1 vccd1 _10463_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12201_ _12367_/B _12201_/B _12201_/C vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__and3_4
XFILLER_108_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _13181_/A _13181_/B vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10393_ _14784_/A _10970_/B _10392_/D _10392_/A vssd1 vssd1 vccd1 vccd1 _10393_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ _12343_/B _12132_/B vssd1 vssd1 vccd1 vccd1 _12145_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16940_ _16317_/A _16165_/B _17119_/C _16809_/C vssd1 vssd1 vccd1 vccd1 _16940_/X
+ sky130_fd_sc_hd__a22o_1
X_12063_ _13837_/A _16011_/B _12063_/C vssd1 vssd1 vccd1 vccd1 _12063_/X sky130_fd_sc_hd__or3_4
XFILLER_81_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _10966_/A _10965_/B _10965_/A vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__o21ba_2
XFILLER_49_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16871_ _17165_/A1 _14481_/X _17164_/C _15460_/X vssd1 vssd1 vccd1 vccd1 _16871_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15822_ _16226_/B _16745_/B _15821_/C _15821_/D vssd1 vssd1 vccd1 vccd1 _15823_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15753_ _16446_/A _15752_/A _16619_/A _16410_/A vssd1 vssd1 vccd1 vccd1 _15753_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12965_ _17415_/A _13551_/D vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__nand2_2
XTAP_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _11916_/A vssd1 vssd1 vccd1 vccd1 _11916_/Y sky130_fd_sc_hd__inv_2
X_14704_ _13516_/X _13519_/B _14840_/A vssd1 vssd1 vccd1 vccd1 _14705_/B sky130_fd_sc_hd__mux2_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15684_ _15580_/B _15582_/B _15580_/A vssd1 vssd1 vccd1 vccd1 _15686_/B sky130_fd_sc_hd__o21ba_1
XFILLER_61_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12897_/A _12897_/B vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__and2b_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17423_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17423_/X sky130_fd_sc_hd__or2_1
X_14635_ _13273_/X _13276_/B _17371_/A vssd1 vssd1 vccd1 vccd1 _14636_/B sky130_fd_sc_hd__mux2_4
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _12442_/A _14933_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__or3_4
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14566_/A _14566_/B vssd1 vssd1 vccd1 vccd1 _14567_/B sky130_fd_sc_hd__nor2_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _13169_/D _17354_/A2 _17353_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17506_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11778_ _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11778_/Y sky130_fd_sc_hd__nand2_2
XFILLER_158_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16305_ _14859_/B _16115_/B _16298_/A vssd1 vssd1 vccd1 vccd1 _16306_/C sky130_fd_sc_hd__a21oi_1
X_13517_ _12401_/A _13516_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13517_/Y sky130_fd_sc_hd__o21ai_1
X_17285_ _17604_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__a21o_1
X_10729_ _10729_/A _10729_/B vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__xor2_4
X_14497_ _14497_/A _14497_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14498_/B sky130_fd_sc_hd__or3_1
XFILLER_146_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16236_ _16595_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16238_/B sky130_fd_sc_hd__nor2_2
XFILLER_146_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13448_ _16723_/A _16722_/A vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__and2_4
XFILLER_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _16619_/A _16168_/B vssd1 vssd1 vccd1 vccd1 _16259_/C sky130_fd_sc_hd__nor2_1
XFILLER_115_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ _13252_/Y _13256_/A _13500_/B _13378_/X vssd1 vssd1 vccd1 vccd1 _13504_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15118_ _15042_/X _15043_/X _15041_/X vssd1 vssd1 vccd1 vccd1 _15119_/B sky130_fd_sc_hd__a21boi_4
X_16098_ _16098_/A vssd1 vssd1 vccd1 vccd1 _16100_/B sky130_fd_sc_hd__clkinv_2
XFILLER_88_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15049_ _16115_/A _15110_/B _15046_/Y _15048_/Y vssd1 vssd1 vccd1 vccd1 _15049_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09610_ _09610_/A _09614_/A _09610_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__or3_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09541_ _09530_/B _09530_/C _09528_/Y _09485_/X vssd1 vssd1 vccd1 vccd1 _09541_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_3_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _09602_/A _09471_/Y _15537_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _09610_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout210 _14911_/B vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__buf_2
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout221 _16991_/A vssd1 vssd1 vccd1 vccd1 _16020_/B sky130_fd_sc_hd__buf_8
XFILLER_114_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout232 _14930_/Y vssd1 vssd1 vccd1 vccd1 _15804_/A2 sky130_fd_sc_hd__buf_6
Xfanout243 _16015_/A vssd1 vssd1 vccd1 vccd1 _17140_/A sky130_fd_sc_hd__buf_4
Xfanout254 _14756_/A1 vssd1 vssd1 vccd1 vccd1 _14763_/S sky130_fd_sc_hd__buf_4
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout265 _16391_/B vssd1 vssd1 vccd1 vccd1 _15891_/B sky130_fd_sc_hd__buf_2
Xfanout276 _08732_/X vssd1 vssd1 vccd1 vccd1 _16911_/A sky130_fd_sc_hd__buf_8
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__xnor2_1
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout287 _08722_/Y vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__buf_6
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout298 _15116_/A vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _09739_/A _09739_/B vssd1 vssd1 vccd1 vccd1 _09740_/C sky130_fd_sc_hd__xnor2_1
XFILLER_189_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ _17385_/A _17383_/A _13300_/D _13169_/D vssd1 vssd1 vccd1 vccd1 _12910_/A
+ sky130_fd_sc_hd__and4_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11701_ _11700_/B _11700_/C _11700_/A vssd1 vssd1 vccd1 vccd1 _15793_/B sky130_fd_sc_hd__a21bo_1
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12681_ _12682_/A _12682_/B vssd1 vssd1 vccd1 vccd1 _12681_/Y sky130_fd_sc_hd__nor2_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14763_/S _14418_/X _14419_/Y _14358_/Y vssd1 vssd1 vccd1 vccd1 _17597_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/A _11632_/B vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__or2_4
XFILLER_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14351_ _14349_/X _14351_/B vssd1 vssd1 vccd1 vccd1 _14416_/B sky130_fd_sc_hd__and2b_1
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ _11564_/A _11562_/Y _11630_/A _11563_/D vssd1 vssd1 vccd1 vccd1 _11590_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_156_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13302_ _17387_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _13303_/B sky130_fd_sc_hd__nand2_4
XFILLER_183_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10514_ _10613_/A _10613_/B vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__and2_2
X_17070_ _17105_/B _17070_/B vssd1 vssd1 vccd1 vccd1 _17070_/Y sky130_fd_sc_hd__nor2_1
X_14282_ _13939_/A _14281_/Y _14280_/X vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _11453_/B _11449_/B _11449_/C vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__a21oi_4
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16021_ _16108_/C _16054_/B vssd1 vssd1 vccd1 vccd1 _16409_/B sky130_fd_sc_hd__nand2_2
X_13233_ _13099_/A _13101_/B _13099_/B vssd1 vssd1 vccd1 vccd1 _13235_/B sky130_fd_sc_hd__o21ba_1
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/C sky130_fd_sc_hd__nor2_1
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13164_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13312_/A sky130_fd_sc_hd__inv_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _11006_/A _11006_/B _10491_/B _10911_/B vssd1 vssd1 vccd1 vccd1 _10379_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_152_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12115_ _12115_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12116_/B sky130_fd_sc_hd__nor2_1
X_13095_ _13095_/A _13095_/B vssd1 vssd1 vccd1 vccd1 _13114_/A sky130_fd_sc_hd__xnor2_1
XFILLER_111_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12046_ _12700_/D _12046_/B vssd1 vssd1 vccd1 vccd1 _12046_/Y sky130_fd_sc_hd__nand2_1
X_16923_ _14865_/B _16868_/A _17140_/A vssd1 vssd1 vccd1 vccd1 _16923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16854_ _16566_/A _16566_/B _16854_/C _16854_/D vssd1 vssd1 vccd1 vccd1 _16854_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _16011_/A _15805_/B vssd1 vssd1 vccd1 vccd1 _15805_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16785_ _16850_/A _16785_/B vssd1 vssd1 vccd1 vccd1 _16786_/B sky130_fd_sc_hd__or2_4
X_13997_ _13997_/A _13997_/B vssd1 vssd1 vccd1 vccd1 _13998_/B sky130_fd_sc_hd__and2_1
XFILLER_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15736_ _16136_/B _16246_/A vssd1 vssd1 vccd1 vccd1 _15737_/B sky130_fd_sc_hd__nand2_4
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _12947_/A _12947_/B _12947_/C vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__o21ai_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15667_ _16536_/A _15667_/B vssd1 vssd1 vccd1 vccd1 _15668_/B sky130_fd_sc_hd__nand2_2
X_12879_ _13643_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ input49/X _17422_/A2 _17405_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17531_/D
+ sky130_fd_sc_hd__o211a_1
X_14618_ _14618_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _14619_/B sky130_fd_sc_hd__nor2_1
X_15598_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15599_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14549_ _14549_/A _14601_/B vssd1 vssd1 vccd1 vccd1 _14570_/A sky130_fd_sc_hd__nor2_2
XFILLER_159_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17337_ input48/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17337_/X sky130_fd_sc_hd__or3_1
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17268_ _17566_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__and2_1
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16219_ _16735_/A _13839_/X _16582_/A _14961_/X vssd1 vssd1 vccd1 vccd1 _16219_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17199_ _17543_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__and2_1
XFILLER_143_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08972_ _08973_/B _09095_/A _08973_/A vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__o21ai_4
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__xnor2_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09455_/A _09455_/B vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__nand2_1
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09386_ _09386_/A _09386_/B vssd1 vssd1 vccd1 vccd1 _09387_/C sky130_fd_sc_hd__xnor2_4
XFILLER_40_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10230_ _10157_/C _10157_/B _10155_/Y vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__a21bo_2
XFILLER_180_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10161_ _10054_/B _10159_/Y _10155_/A _10137_/X vssd1 vssd1 vccd1 vccd1 _10161_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _10091_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13920_ _13921_/A _13921_/B _13921_/C vssd1 vssd1 vccd1 vccd1 _13922_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13851_ _13851_/A _13958_/A vssd1 vssd1 vccd1 vccd1 _13853_/B sky130_fd_sc_hd__nor2_2
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12802_ _12619_/A _12621_/B _12619_/B vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__o21ba_4
XFILLER_142_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13782_ _13681_/B _13683_/B _13681_/A vssd1 vssd1 vccd1 vccd1 _13784_/B sky130_fd_sc_hd__o21ba_1
X_16570_ _14774_/A _16644_/B _16571_/A vssd1 vssd1 vccd1 vccd1 _16572_/A sky130_fd_sc_hd__a21bo_1
XFILLER_76_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10994_ _14794_/A _10993_/D _11164_/A _10992_/Y vssd1 vssd1 vccd1 vccd1 _10996_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12733_ _17389_/A _12578_/B _12576_/C _17391_/A vssd1 vssd1 vccd1 vccd1 _12735_/A
+ sky130_fd_sc_hd__a22oi_2
X_15521_ _15519_/X _15521_/B vssd1 vssd1 vccd1 vccd1 _15522_/B sky130_fd_sc_hd__nand2b_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _15532_/A _15453_/B _15453_/C vssd1 vssd1 vccd1 vccd1 _15454_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12504_/A _12506_/B _12504_/B vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__o21ba_1
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14424_/A vssd1 vssd1 vccd1 vccd1 _14405_/B sky130_fd_sc_hd__inv_2
X_11615_ _11614_/A _11614_/B _11614_/C vssd1 vssd1 vccd1 vccd1 _11617_/C sky130_fd_sc_hd__a21oi_2
XFILLER_168_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15383_ _10799_/Y _14931_/X _15382_/X _16977_/A vssd1 vssd1 vccd1 vccd1 _15383_/X
+ sky130_fd_sc_hd__o211a_1
X_12595_ _12595_/A _12595_/B _12595_/C _12736_/B vssd1 vssd1 vccd1 vccd1 _12755_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14334_ _14239_/A _14256_/X _14332_/X _14333_/Y vssd1 vssd1 vccd1 vccd1 _14405_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_168_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17122_ _17091_/A _17118_/A _17089_/A vssd1 vssd1 vccd1 vccd1 _17124_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11546_ _11461_/B _11544_/Y _11543_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11547_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _17091_/A _17053_/B vssd1 vssd1 vccd1 vccd1 _17093_/B sky130_fd_sc_hd__nand2b_2
X_14265_ _14265_/A _14265_/B _14266_/B vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__and3_1
XFILLER_100_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11477_ _11477_/A _11514_/A _11477_/C vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__and3_4
XFILLER_109_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16004_ _16004_/A _16004_/B vssd1 vssd1 vccd1 vccd1 _16004_/Y sky130_fd_sc_hd__xnor2_1
X_13216_ _17407_/A _13564_/D _13216_/C vssd1 vssd1 vccd1 vccd1 _13346_/B sky130_fd_sc_hd__nand3_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _12398_/S _10431_/B _10312_/A _10310_/Y vssd1 vssd1 vccd1 vccd1 _10429_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14196_ _14197_/A _14197_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _14276_/A sky130_fd_sc_hd__a21oi_2
XFILLER_112_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ _13948_/B _14153_/C _13566_/B _13948_/A vssd1 vssd1 vccd1 vccd1 _13149_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _11027_/B _10912_/C vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__nand2_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _12979_/A _12978_/B _12978_/A vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__a21bo_2
XFILLER_140_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16906_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16908_/B sky130_fd_sc_hd__nand2_1
X_12029_ _12700_/C _12700_/D vssd1 vssd1 vccd1 vccd1 _12035_/C sky130_fd_sc_hd__nand2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16837_ _16762_/A _16762_/B _16765_/A vssd1 vssd1 vccd1 vccd1 _16838_/B sky130_fd_sc_hd__a21o_1
XFILLER_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16768_ _16768_/A _16835_/B vssd1 vssd1 vccd1 vccd1 _16770_/C sky130_fd_sc_hd__nor2_1
XFILLER_81_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15719_ _16917_/A _15705_/Y _15706_/X _15718_/X vssd1 vssd1 vccd1 vccd1 _15719_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_22_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16699_ _16699_/A _16699_/B vssd1 vssd1 vccd1 vccd1 _16701_/B sky130_fd_sc_hd__xnor2_1
X_09240_ _09240_/A _09240_/B vssd1 vssd1 vccd1 vccd1 _09242_/C sky130_fd_sc_hd__xnor2_1
XFILLER_178_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ _09178_/A _09178_/B _09178_/C vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__a21oi_4
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08955_ _08958_/A vssd1 vssd1 vccd1 vccd1 _08957_/C sky130_fd_sc_hd__inv_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _09030_/A _11867_/B _12171_/B _12166_/B vssd1 vssd1 vccd1 vccd1 _08887_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09507_/Y sky130_fd_sc_hd__nor2_2
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09439_/B sky130_fd_sc_hd__nor2_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09369_ _09370_/B _09370_/C _09370_/A vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__a21o_4
XFILLER_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _11403_/B _11400_/B _11400_/C vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__and3_4
XFILLER_184_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _16922_/A _12380_/B vssd1 vssd1 vccd1 vccd1 _12380_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_70 _17529_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_81 _17461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_92 _12088_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11331_/A _11331_/B _11331_/C vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__nand3_2
XFILLER_158_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14050_ _14050_/A _14050_/B _14141_/D _14050_/D vssd1 vssd1 vccd1 vccd1 _14158_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_158_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11262_ _11553_/B _11391_/B _11125_/A _11123_/Y vssd1 vssd1 vccd1 vccd1 _11264_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _13001_/A _13001_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__and3_1
X_10213_ _10194_/A _10194_/B _10194_/C vssd1 vssd1 vccd1 vccd1 _10214_/C sky130_fd_sc_hd__o21a_1
XFILLER_122_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11193_ _11222_/B _11191_/X _11067_/Y _11069_/X vssd1 vssd1 vccd1 vccd1 _11194_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_97_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10144_ _10508_/C _10743_/C vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__nand2_1
X_14952_ _14952_/A _14952_/B vssd1 vssd1 vccd1 vccd1 _14952_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13903_ _14326_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _13904_/B sky130_fd_sc_hd__nand2_2
XFILLER_130_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ _15262_/B _15472_/A _15071_/A vssd1 vssd1 vccd1 vccd1 _14888_/D sky130_fd_sc_hd__or3b_1
XFILLER_78_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16622_ _16622_/A _16622_/B _16622_/C vssd1 vssd1 vccd1 vccd1 _16623_/B sky130_fd_sc_hd__nor3_1
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16553_ _16554_/A _16554_/B vssd1 vssd1 vccd1 vccd1 _16636_/B sky130_fd_sc_hd__nand2b_1
X_13765_ _13765_/A _13765_/B vssd1 vssd1 vccd1 vccd1 _13767_/A sky130_fd_sc_hd__nor2_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10977_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10977_/X sky130_fd_sc_hd__or2_2
XFILLER_189_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15504_ _15504_/A _15504_/B vssd1 vssd1 vccd1 vccd1 _15505_/B sky130_fd_sc_hd__xor2_4
X_12716_ _17401_/A _13564_/D vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__nand2_2
X_13696_ _13695_/A _13695_/B _13695_/C vssd1 vssd1 vccd1 vccd1 _13800_/A sky130_fd_sc_hd__o21ai_2
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16484_ _12560_/A _14775_/X _14816_/X vssd1 vssd1 vccd1 vccd1 _16485_/B sky130_fd_sc_hd__a21o_1
XFILLER_189_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12647_ _12798_/B _12647_/B vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__nand2_1
X_15435_ _15436_/A _15436_/B vssd1 vssd1 vccd1 vccd1 _15520_/A sky130_fd_sc_hd__and2_1
XFILLER_30_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15366_ _15365_/B _15366_/B vssd1 vssd1 vccd1 vccd1 _15367_/B sky130_fd_sc_hd__nand2b_1
XFILLER_191_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12578_ _12578_/A _12578_/B vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17105_ _17105_/A _17105_/B vssd1 vssd1 vccd1 vccd1 _17105_/Y sky130_fd_sc_hd__nor2_1
X_14317_ _14318_/B _14318_/C _14641_/D _14450_/A vssd1 vssd1 vccd1 vccd1 _14319_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_157_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11530_/C sky130_fd_sc_hd__xnor2_4
X_15297_ _15228_/A _15228_/B _15231_/A vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__o21a_1
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14248_ _14248_/A _14599_/D _14248_/C vssd1 vssd1 vccd1 vccd1 _14330_/B sky130_fd_sc_hd__nand3_4
X_17036_ _17028_/A _17170_/B1 _17035_/X vssd1 vssd1 vccd1 vccd1 _17570_/D sky130_fd_sc_hd__a21oi_1
XFILLER_98_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14179_ _14180_/A _14180_/B vssd1 vssd1 vccd1 vccd1 _14273_/A sky130_fd_sc_hd__nand2b_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout809 _12338_/C vssd1 vssd1 vccd1 vccd1 _09509_/B sky130_fd_sc_hd__buf_8
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _14836_/A _14933_/A vssd1 vssd1 vccd1 vccd1 _08740_/Y sky130_fd_sc_hd__nor2_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09223_ _09223_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__nor2_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _09131_/X _09138_/X _09152_/A _09153_/X vssd1 vssd1 vccd1 vccd1 _09155_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_175_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09085_ _12135_/A _12135_/B _11808_/B _09926_/B vssd1 vssd1 vccd1 vccd1 _09317_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_147_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ _11026_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _09988_/B sky130_fd_sc_hd__nand2_4
XFILLER_89_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08938_ _08923_/A _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__o21ba_1
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08869_ _08869_/A _08869_/B _08869_/C vssd1 vssd1 vccd1 vccd1 _08869_/Y sky130_fd_sc_hd__nand3_2
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _10899_/C _10899_/D _10995_/A _10898_/Y vssd1 vssd1 vccd1 vccd1 _10902_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_123_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11880_ _12256_/B _12565_/D _11881_/D _12256_/A vssd1 vssd1 vccd1 vccd1 _11882_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ _11072_/B _11072_/C _11072_/A vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__a21o_2
XFILLER_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _14050_/B _13664_/D _13551_/D _14050_/A vssd1 vssd1 vccd1 vccd1 _13552_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ _10760_/A _10761_/Y _10771_/A _10734_/X vssd1 vssd1 vccd1 vccd1 _10771_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_38_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12501_ _12501_/A _12501_/B vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__xnor2_4
XFILLER_186_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13481_ _13482_/A _13482_/B vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__nand2_2
X_10693_ _10632_/B _10632_/C _10632_/D _10632_/A vssd1 vssd1 vccd1 vccd1 _10693_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15220_ _15220_/A _15220_/B vssd1 vssd1 vccd1 vccd1 _15221_/B sky130_fd_sc_hd__xnor2_4
XFILLER_185_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12432_ _12432_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12434_/C sky130_fd_sc_hd__xnor2_4
XFILLER_173_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _15152_/B _15175_/B _16991_/A vssd1 vssd1 vccd1 vccd1 _15151_/X sky130_fd_sc_hd__and3b_2
X_12363_ _12190_/A _12189_/A _12189_/B _12191_/X vssd1 vssd1 vccd1 vccd1 _12364_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_126_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14194_/A _14102_/B vssd1 vssd1 vccd1 vccd1 _14104_/B sky130_fd_sc_hd__xnor2_1
X_11314_ _11314_/A _11423_/A _15402_/A _11370_/C vssd1 vssd1 vccd1 vccd1 _11314_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_181_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15082_ _15278_/A _15821_/A _15342_/A vssd1 vssd1 vccd1 vccd1 _15164_/B sky130_fd_sc_hd__and3_1
XFILLER_180_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ _12770_/B _12463_/D _12295_/D _12618_/A vssd1 vssd1 vccd1 vccd1 _12296_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _14122_/B _14034_/B vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__or2_1
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11245_ _11260_/C _14906_/B _11118_/A _11116_/Y vssd1 vssd1 vccd1 vccd1 _11246_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _11176_/A _11176_/B _11176_/C vssd1 vssd1 vccd1 vccd1 _11176_/X sky130_fd_sc_hd__or3_4
XFILLER_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10127_ _10254_/B _10392_/D _10377_/B _10254_/A vssd1 vssd1 vccd1 vccd1 _10128_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15984_ _15984_/A _15984_/B vssd1 vssd1 vccd1 vccd1 _15987_/A sky130_fd_sc_hd__xnor2_2
X_10058_ _10057_/B _10057_/C _10057_/A vssd1 vssd1 vccd1 vccd1 _10059_/C sky130_fd_sc_hd__a21boi_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14935_ _10560_/D _15108_/A _15248_/C _14934_/X vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14866_ _17028_/A _17028_/B vssd1 vssd1 vccd1 vccd1 _17029_/B sky130_fd_sc_hd__and2_2
XFILLER_35_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16605_ _16827_/B _16681_/C _16514_/C _16603_/X vssd1 vssd1 vccd1 vccd1 _16607_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13817_ _13817_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _13820_/A sky130_fd_sc_hd__xnor2_4
XFILLER_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17585_ fanout935/X _17585_/D vssd1 vssd1 vccd1 vccd1 _17585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14797_ _14796_/B _14796_/C _14796_/D _11595_/B vssd1 vssd1 vccd1 vccd1 _14797_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_189_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16536_ _16536_/A _16695_/B _16537_/A vssd1 vssd1 vccd1 vccd1 _16622_/B sky130_fd_sc_hd__and3_1
X_13748_ _13748_/A _13748_/B vssd1 vssd1 vccd1 vccd1 _13751_/A sky130_fd_sc_hd__xnor2_4
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16467_ _16369_/A _16369_/B _16371_/Y vssd1 vssd1 vccd1 vccd1 _16469_/B sky130_fd_sc_hd__a21bo_1
XFILLER_176_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ _13680_/A _13680_/B _13680_/C vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__o21a_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15418_ _15501_/A _15418_/B _15419_/B vssd1 vssd1 vccd1 vccd1 _15501_/B sky130_fd_sc_hd__and3b_1
XFILLER_164_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16398_ _16398_/A _16398_/B vssd1 vssd1 vccd1 vccd1 _16398_/X sky130_fd_sc_hd__xor2_1
XFILLER_191_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15349_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__nor2_4
XFILLER_144_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17019_ _17028_/A _17153_/B _14766_/A vssd1 vssd1 vccd1 vccd1 _17066_/A sky130_fd_sc_hd__or3b_2
X_09910_ _09910_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09912_/C sky130_fd_sc_hd__nor2_2
XFILLER_125_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout606 _11437_/B vssd1 vssd1 vccd1 vccd1 _11561_/B sky130_fd_sc_hd__buf_4
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _09841_/A _09983_/A vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__nor2_4
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout617 _17508_/Q vssd1 vssd1 vccd1 vccd1 _17139_/A sky130_fd_sc_hd__clkbuf_16
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout628 _08968_/B vssd1 vssd1 vccd1 vccd1 _13300_/D sky130_fd_sc_hd__buf_6
Xfanout639 _14593_/C vssd1 vssd1 vccd1 vccd1 _14641_/D sky130_fd_sc_hd__clkbuf_8
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09773_/C _09812_/A vssd1 vssd1 vccd1 vccd1 _09772_/X sky130_fd_sc_hd__and2b_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _11629_/B vssd1 vssd1 vccd1 vccd1 _08723_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ _09206_/A _09375_/A vssd1 vssd1 vccd1 vccd1 _09208_/B sky130_fd_sc_hd__nor2_1
XFILLER_176_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09137_ _09167_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09170_/B sky130_fd_sc_hd__xnor2_4
XFILLER_108_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _09062_/X _09294_/A _09076_/A _09055_/Y vssd1 vssd1 vccd1 vccd1 _09076_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11030_ _11030_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _11032_/B sky130_fd_sc_hd__xnor2_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12981_ _12981_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _12983_/B sky130_fd_sc_hd__xnor2_1
XTAP_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14719_/A _14719_/B _14719_/C vssd1 vssd1 vccd1 vccd1 _14721_/B sky130_fd_sc_hd__o21ai_1
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11932_ _11932_/A _12592_/C vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__nand2_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14710_/C _14651_/B vssd1 vssd1 vccd1 vccd1 _14693_/B sky130_fd_sc_hd__xnor2_4
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _12237_/A _12171_/B _08748_/A _08747_/A vssd1 vssd1 vccd1 vccd1 _11865_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13603_/A _13603_/B _13603_/C vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__a21oi_4
X_10814_ _10814_/A _10814_/B vssd1 vssd1 vccd1 vccd1 _10816_/B sky130_fd_sc_hd__xnor2_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ input61/X _17377_/B _17369_/Y _17372_/C1 vssd1 vssd1 vccd1 vccd1 _17513_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _14582_/A vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__inv_2
X_11794_ _14771_/A _16723_/A _16644_/C _14774_/A vssd1 vssd1 vccd1 vccd1 _11798_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16321_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__xor2_1
XFILLER_185_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13533_ _13643_/A _13745_/D vssd1 vssd1 vccd1 vccd1 _13534_/B sky130_fd_sc_hd__nand2_2
X_10745_ _10746_/A _10744_/Y _11124_/C _10745_/D vssd1 vssd1 vccd1 vccd1 _10984_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_159_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16252_ _16252_/A _16252_/B vssd1 vssd1 vccd1 vccd1 _16254_/B sky130_fd_sc_hd__xnor2_4
X_13464_ _17405_/A _16789_/A vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ _10556_/B _10587_/Y wire120/X _10667_/Y vssd1 vssd1 vccd1 vccd1 _10677_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_159_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15203_ _14877_/Y _14967_/D _15143_/A vssd1 vssd1 vccd1 vccd1 _15203_/X sky130_fd_sc_hd__a21o_2
X_12415_ _12415_/A _12415_/B vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__nor2_2
X_16183_ _16183_/A _16183_/B _16183_/C vssd1 vssd1 vccd1 vccd1 _16184_/B sky130_fd_sc_hd__nor3_1
X_13395_ _13844_/B _13523_/B _13895_/C _13844_/A vssd1 vssd1 vccd1 vccd1 _13398_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12346_ _12346_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__xor2_1
X_15134_ _15116_/A _15131_/A _15130_/X _10171_/B vssd1 vssd1 vccd1 vccd1 _15134_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_182_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ _14963_/X _15040_/X _15044_/Y _15045_/X vssd1 vssd1 vccd1 vccd1 _15065_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_142_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12277_ _17381_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__nand2_2
XFILLER_142_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14016_ _14016_/A _14016_/B vssd1 vssd1 vccd1 vccd1 _14018_/C sky130_fd_sc_hd__xor2_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__xor2_4
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11159_ _11159_/A _11159_/B vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__xnor2_4
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15967_ _16084_/A _15967_/B vssd1 vssd1 vccd1 vccd1 _15969_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14918_ _15131_/A _14918_/B vssd1 vssd1 vccd1 vccd1 _14918_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15898_ _15898_/A _15898_/B vssd1 vssd1 vccd1 vccd1 _15898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14849_ _14906_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15381_/B sky130_fd_sc_hd__and2_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17568_ fanout942/X _17568_/D vssd1 vssd1 vccd1 vccd1 _17568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16519_ _16519_/A _16519_/B _16519_/C vssd1 vssd1 vccd1 vccd1 _16520_/B sky130_fd_sc_hd__and3_1
XFILLER_149_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17499_ fanout932/X _17499_/D vssd1 vssd1 vccd1 vccd1 _17499_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout403 _17530_/Q vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__buf_6
XFILLER_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout414 _10236_/B vssd1 vssd1 vccd1 vccd1 _10235_/A sky130_fd_sc_hd__buf_6
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout425 _17527_/Q vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__buf_8
XFILLER_101_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout436 _13405_/B vssd1 vssd1 vccd1 vccd1 _13745_/B sky130_fd_sc_hd__buf_6
XFILLER_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _09825_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__nor2_4
Xfanout447 _12256_/A vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__buf_8
Xfanout458 _17523_/Q vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__buf_12
XFILLER_150_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout469 _10904_/B vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__buf_12
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09755_ _12135_/A _12135_/B _10431_/B _10543_/B vssd1 vssd1 vccd1 vccd1 _09890_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09686_ _09686_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09768_/A sky130_fd_sc_hd__xnor2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10530_ _10531_/A _10531_/C vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__nor2_2
XFILLER_122_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10461_ _10336_/Y _10353_/X _10459_/A _10459_/Y vssd1 vssd1 vccd1 vccd1 _10461_/X
+ sky130_fd_sc_hd__o211a_2
X_12200_ _12200_/A _12200_/B vssd1 vssd1 vccd1 vccd1 _12201_/C sky130_fd_sc_hd__or2_2
XFILLER_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13180_ _13177_/Y _13312_/B _13046_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13189_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_124_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10392_ _10392_/A _14784_/A _10970_/B _10392_/D vssd1 vssd1 vccd1 vccd1 _10395_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12132_/B sky130_fd_sc_hd__and2_1
XFILLER_124_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ _12397_/B _12061_/Y _12383_/S vssd1 vssd1 vccd1 vccd1 _12063_/C sky130_fd_sc_hd__mux2_1
XFILLER_150_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11013_ _11013_/A _11013_/B vssd1 vssd1 vccd1 vccd1 _11016_/A sky130_fd_sc_hd__nor2_4
XFILLER_89_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16870_ _14770_/A _14864_/A _17075_/A2 _16869_/X vssd1 vssd1 vccd1 vccd1 _16872_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15821_ _15821_/A _16745_/B _15821_/C _15821_/D vssd1 vssd1 vccd1 vccd1 _15821_/X
+ sky130_fd_sc_hd__and4_1
XTAP_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15752_/A _15752_/B vssd1 vssd1 vccd1 vccd1 _15853_/A sky130_fd_sc_hd__nor2_8
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _12964_/A _12964_/B vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__nor2_1
XFILLER_161_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14756_/A1 _14700_/Y _14702_/Y _14667_/Y _14668_/X vssd1 vssd1 vccd1 vccd1
+ _17603_/D sky130_fd_sc_hd__a32o_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _11915_/A _11915_/B _12148_/B _11913_/X vssd1 vssd1 vccd1 vccd1 _11916_/A
+ sky130_fd_sc_hd__or4bb_4
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15769_/B _15682_/B _15682_/C vssd1 vssd1 vccd1 vccd1 _15690_/B sky130_fd_sc_hd__o21a_2
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A _12895_/B vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__xnor2_2
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ input57/X _17422_/A2 _17421_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17539_/D
+ sky130_fd_sc_hd__o211a_1
X_14634_ _14756_/A1 _14632_/X _14638_/B _14590_/Y _14591_/X vssd1 vssd1 vccd1 vccd1
+ _17601_/D sky130_fd_sc_hd__a32o_1
XFILLER_127_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _12442_/A _14933_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _13626_/B sky130_fd_sc_hd__nor3_4
XFILLER_54_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ input56/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__or3_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14565_/A _14565_/B vssd1 vssd1 vccd1 vccd1 _14566_/B sky130_fd_sc_hd__nor2_1
X_11777_ _10098_/A _11778_/B _11778_/A vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_186_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16304_ _16304_/A _16304_/B _16304_/C vssd1 vssd1 vccd1 vccd1 _16310_/A sky130_fd_sc_hd__or3_1
XFILLER_158_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10728_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__nand2_4
X_13516_ _12543_/X _12552_/B _13516_/S vssd1 vssd1 vccd1 vccd1 _13516_/X sky130_fd_sc_hd__mux2_4
X_17284_ _17462_/Q _17293_/A2 _17282_/X _17283_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17462_/D sky130_fd_sc_hd__o221a_1
X_14496_ _14497_/A _14497_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__o21ai_2
XFILLER_146_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16235_ _16235_/A _16339_/A vssd1 vssd1 vccd1 vccd1 _16238_/A sky130_fd_sc_hd__and2_2
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13447_ _13444_/A _13445_/Y _13329_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13490_/B
+ sky130_fd_sc_hd__o211a_2
X_10659_ _10660_/A _10658_/Y _10993_/C _10659_/D vssd1 vssd1 vccd1 vccd1 _10757_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_139_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16166_ _15746_/X _16164_/Y _16279_/A vssd1 vssd1 vccd1 vccd1 _16175_/A sky130_fd_sc_hd__a21oi_4
XFILLER_154_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13378_ _13500_/A _13376_/X _13246_/A _13249_/C vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15117_ _15117_/A _15117_/B vssd1 vssd1 vccd1 vccd1 _15119_/A sky130_fd_sc_hd__nand2_1
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _12795_/A _12637_/C _12328_/C vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16097_ _16096_/A _16096_/B _16096_/C vssd1 vssd1 vccd1 vccd1 _16098_/A sky130_fd_sc_hd__o21ai_4
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15048_ _14796_/B _15899_/A2 _15047_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15048_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16999_ _17000_/A _17000_/B vssd1 vssd1 vccd1 vccd1 _17052_/B sky130_fd_sc_hd__and2_1
XFILLER_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09540_ _09540_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09471_ _12135_/B _09928_/D _10309_/B _12135_/A vssd1 vssd1 vccd1 vccd1 _09471_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout200 _13841_/A vssd1 vssd1 vccd1 vccd1 _14210_/B sky130_fd_sc_hd__buf_4
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout211 _14911_/B vssd1 vssd1 vccd1 vccd1 _12700_/D sky130_fd_sc_hd__buf_4
Xfanout222 _17083_/A vssd1 vssd1 vccd1 vccd1 _16991_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout233 _16580_/A2 vssd1 vssd1 vccd1 vccd1 _17162_/A2 sky130_fd_sc_hd__buf_4
Xfanout244 _16015_/A vssd1 vssd1 vccd1 vccd1 _16652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout255 _16389_/A vssd1 vssd1 vccd1 vccd1 _14756_/A1 sky130_fd_sc_hd__buf_4
XFILLER_189_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout266 _16391_/B vssd1 vssd1 vccd1 vccd1 _17153_/B sky130_fd_sc_hd__buf_4
X_09807_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09807_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout277 _08727_/Y vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__buf_8
Xfanout288 _15384_/S vssd1 vssd1 vccd1 vccd1 _17367_/A sky130_fd_sc_hd__buf_6
Xfanout299 _08720_/Y vssd1 vssd1 vccd1 vccd1 _15116_/A sky130_fd_sc_hd__buf_6
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09738_ _09732_/X _09868_/A _09724_/X _09725_/Y vssd1 vssd1 vccd1 vccd1 _09740_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_189_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ _09668_/A _09668_/Y _09530_/X _09541_/X vssd1 vssd1 vccd1 vccd1 _09674_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11700_/A _11700_/B _11700_/C vssd1 vssd1 vccd1 vccd1 _11700_/Y sky130_fd_sc_hd__nand3_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ _12522_/B _12522_/C _12522_/A vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__o21ba_2
XFILLER_131_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11629_/B _15116_/B _14794_/B _11629_/A vssd1 vssd1 vccd1 vccd1 _11632_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14350_ _14350_/A _14350_/B _14350_/C vssd1 vssd1 vccd1 vccd1 _14351_/B sky130_fd_sc_hd__or3_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _11561_/B _11561_/C _11561_/D _11561_/A vssd1 vssd1 vccd1 vccd1 _11562_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13301_ _13301_/A _13301_/B vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__nor2_2
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10513_ _10513_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10613_/B sky130_fd_sc_hd__nor2_2
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14281_ _14281_/A _14281_/B vssd1 vssd1 vccd1 vccd1 _14281_/Y sky130_fd_sc_hd__nand2_2
X_11493_ _11496_/B _11493_/B _11493_/C vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__and3_2
XFILLER_183_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16020_ _16108_/C _16020_/B vssd1 vssd1 vccd1 vccd1 _17119_/C sky130_fd_sc_hd__and2_4
X_13232_ _13232_/A _13232_/B vssd1 vssd1 vccd1 vccd1 _13235_/A sky130_fd_sc_hd__xnor2_1
X_10444_ _10560_/A _10321_/C _10560_/D _10321_/A vssd1 vssd1 vccd1 vccd1 _10445_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13163_ _13165_/A _13165_/B _13165_/C vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__a21o_2
XFILLER_40_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10375_ _10390_/A _10375_/B vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__and2_2
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12114_ _12115_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12116_/A sky130_fd_sc_hd__and2_2
X_13094_ _17405_/A _13094_/B vssd1 vssd1 vccd1 vccd1 _13095_/B sky130_fd_sc_hd__nand2_1
XFILLER_152_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16922_ _16922_/A _16922_/B vssd1 vssd1 vccd1 vccd1 _16922_/Y sky130_fd_sc_hd__nand2_2
X_12045_ _11841_/A _11334_/C _11387_/C vssd1 vssd1 vccd1 vccd1 _12046_/B sky130_fd_sc_hd__a21o_1
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16853_ _16853_/A _16853_/B _16853_/C vssd1 vssd1 vccd1 vccd1 _16854_/D sky130_fd_sc_hd__and3_2
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15804_ _16809_/B _15804_/A2 _15803_/X vssd1 vssd1 vccd1 vccd1 _15804_/Y sky130_fd_sc_hd__a21oi_1
X_16784_ _16784_/A _16784_/B _16784_/C vssd1 vssd1 vccd1 vccd1 _16785_/B sky130_fd_sc_hd__and3_1
XFILLER_168_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13996_ _13997_/A _13997_/B vssd1 vssd1 vccd1 vccd1 _13998_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15735_ _15735_/A _15735_/B vssd1 vssd1 vccd1 vccd1 _15737_/A sky130_fd_sc_hd__nand2_4
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12947_/A _12947_/B _12947_/C vssd1 vssd1 vccd1 vccd1 _12949_/A sky130_fd_sc_hd__or3_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _15666_/A _15666_/B vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__xnor2_4
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12878_/A _13040_/A vssd1 vssd1 vccd1 vccd1 _12881_/A sky130_fd_sc_hd__or2_1
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17405_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17405_/X sky130_fd_sc_hd__or2_1
X_14617_ _14618_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _14658_/B sky130_fd_sc_hd__and2_1
X_11829_ _12031_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nand2_1
X_15597_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15599_/A sky130_fd_sc_hd__or2_4
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17336_ _13088_/B _17360_/A2 _17335_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17497_/D
+ sky130_fd_sc_hd__o211a_1
X_14548_ _14548_/A _14601_/A _14548_/C vssd1 vssd1 vccd1 vccd1 _14601_/B sky130_fd_sc_hd__nor3_2
XFILLER_187_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17267_ _17598_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17267_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14479_ _14479_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14479_/Y sky130_fd_sc_hd__nand2_1
X_16218_ _14778_/X _16580_/A2 _14933_/Y _14859_/B _16218_/C1 vssd1 vssd1 vccd1 vccd1
+ _16218_/X sky130_fd_sc_hd__a221o_1
XFILLER_146_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17198_ input25/X input28/X _17198_/C _17428_/C vssd1 vssd1 vccd1 vccd1 _17198_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16149_ _16041_/A _16039_/B _16150_/B _16595_/A vssd1 vssd1 vccd1 vccd1 _16149_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_143_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _08993_/C _08973_/B _08971_/C vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__nor3_4
XFILLER_170_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09523_ _09523_/A _09523_/B vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09454_ _09448_/X _09579_/A _09440_/X _09441_/Y vssd1 vssd1 vccd1 vccd1 _09455_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _09385_/A _09385_/B vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__xnor2_4
XFILLER_71_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _10137_/X _10155_/A _10159_/Y _10054_/B vssd1 vssd1 vccd1 vccd1 _10207_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ _10091_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__nor3_4
XFILLER_86_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13850_ _13849_/A _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13958_/A sky130_fd_sc_hd__o21a_2
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ _12801_/A _12801_/B vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__xnor2_4
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13781_ _13781_/A _13781_/B vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__xor2_1
XFILLER_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10993_ _11164_/A _10992_/Y _10993_/C _10993_/D vssd1 vssd1 vccd1 vccd1 _11164_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _15520_/A _15520_/B _15520_/C vssd1 vssd1 vccd1 vccd1 _15521_/B sky130_fd_sc_hd__or3_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12732_ _12566_/A _12568_/B _12566_/B vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__o21ba_1
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15451_ _15374_/B _15375_/X _15374_/A vssd1 vssd1 vccd1 vccd1 _15453_/C sky130_fd_sc_hd__o21bai_2
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12663_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__nor2_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14296_/X _14337_/Y _14399_/X _14466_/B vssd1 vssd1 vccd1 vccd1 _14424_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11614_ _11614_/A _11614_/B _11614_/C vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__and3_4
X_15382_ _15381_/A _15713_/B1 _14929_/X _14803_/A vssd1 vssd1 vccd1 vccd1 _15382_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12594_ _12595_/B _12595_/C _12736_/B _17385_/A vssd1 vssd1 vccd1 vccd1 _12596_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _17121_/A _17121_/B vssd1 vssd1 vccd1 vccd1 _17124_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14333_ _14333_/A _14333_/B vssd1 vssd1 vccd1 vccd1 _14333_/Y sky130_fd_sc_hd__nand2_2
X_11545_ _11502_/B _11543_/A _11544_/Y _11461_/B vssd1 vssd1 vccd1 vccd1 _11705_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17052_ _17052_/A _17052_/B _17050_/X vssd1 vssd1 vccd1 vccd1 _17053_/B sky130_fd_sc_hd__or3b_1
X_14264_ _14190_/A _14190_/B _14151_/A vssd1 vssd1 vccd1 vccd1 _14266_/B sky130_fd_sc_hd__a21o_2
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11476_ _11433_/A _11433_/C _11433_/B vssd1 vssd1 vccd1 vccd1 _11477_/C sky130_fd_sc_hd__a21o_2
XFILLER_100_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _16004_/A _16004_/B vssd1 vssd1 vccd1 vccd1 _16003_/X sky130_fd_sc_hd__or2_2
XFILLER_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10427_ _10427_/A _10427_/B _10427_/C vssd1 vssd1 vccd1 vccd1 _10437_/B sky130_fd_sc_hd__nand3_2
X_13215_ _13215_/A _13346_/A vssd1 vssd1 vccd1 vccd1 _13216_/C sky130_fd_sc_hd__and2_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14195_ _14195_/A _14195_/B vssd1 vssd1 vccd1 vccd1 _14197_/C sky130_fd_sc_hd__xor2_2
XFILLER_124_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ _10358_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__xnor2_4
X_13146_ _17371_/A _13516_/S _12037_/A _13145_/Y _15457_/A vssd1 vssd1 vccd1 vccd1
+ _13146_/X sky130_fd_sc_hd__a311o_1
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13074_/X _13075_/Y _12933_/B _12935_/A vssd1 vssd1 vccd1 vccd1 _13121_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_183_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__nand2_2
XFILLER_111_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16905_ _16905_/A _16905_/B vssd1 vssd1 vccd1 vccd1 _16908_/A sky130_fd_sc_hd__xnor2_4
X_12028_ _12020_/Y _12022_/Y _12024_/Y _12026_/Y _15038_/A _15312_/S vssd1 vssd1 vccd1
+ vccd1 _12028_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16836_ _16836_/A _16836_/B vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__nor2_2
XFILLER_65_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16767_ _16767_/A _16767_/B vssd1 vssd1 vccd1 vccd1 _16835_/B sky130_fd_sc_hd__nor2_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13979_ _14226_/A _14063_/C vssd1 vssd1 vccd1 vccd1 _13980_/B sky130_fd_sc_hd__nand2_4
XFILLER_80_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15718_ _16485_/A _15707_/Y _15708_/X _15717_/Y vssd1 vssd1 vccd1 vccd1 _15718_/X
+ sky130_fd_sc_hd__a31o_1
X_16698_ _16698_/A _16698_/B vssd1 vssd1 vccd1 vccd1 _16699_/B sky130_fd_sc_hd__and2_1
XFILLER_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15649_ _16226_/B _16246_/A _15557_/A _15554_/Y vssd1 vssd1 vccd1 vccd1 _15651_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09170_ _09170_/A _09170_/B vssd1 vssd1 vccd1 vccd1 _09178_/C sky130_fd_sc_hd__xor2_4
X_17319_ input38/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17319_/X sky130_fd_sc_hd__or3_1
XFILLER_174_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08954_ _17373_/A _11930_/B _09652_/B _11808_/B vssd1 vssd1 vccd1 vccd1 _08958_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_69_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08885_ _11867_/B _12171_/B _12166_/B _09030_/A vssd1 vssd1 vccd1 vccd1 _08887_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09506_ _09499_/Y _09658_/A _09500_/X vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__a21boi_4
XFILLER_53_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ _09437_/A _09437_/B _09456_/B vssd1 vssd1 vccd1 vccd1 _09437_/X sky130_fd_sc_hd__and3_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ _09498_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09370_/C sky130_fd_sc_hd__nand2_1
XFILLER_36_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09299_ _12107_/A _12595_/B _11867_/C _12795_/B vssd1 vssd1 vccd1 vccd1 _09302_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA_60 _17377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_71 i_wb_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_82 _17436_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11331_/B _11331_/C _11331_/A vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__a21o_1
XFILLER_193_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_93 _15101_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11261_ _11261_/A _11304_/A vssd1 vssd1 vccd1 vccd1 _11270_/A sky130_fd_sc_hd__nor2_4
XFILLER_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10214_/B sky130_fd_sc_hd__xnor2_2
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13000_ _13001_/A _13001_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__a21oi_2
XFILLER_97_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11192_ _11067_/Y _11069_/X _11222_/B _11191_/X vssd1 vssd1 vccd1 vccd1 _11194_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _10145_/A _15707_/A vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__nor2_2
XFILLER_97_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14951_ _15180_/B _14950_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15460_/B sky130_fd_sc_hd__mux2_1
XFILLER_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13902_ _13902_/A _13902_/B vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__nand2_4
XFILLER_43_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14882_ _15262_/A _15262_/C _15262_/D vssd1 vssd1 vccd1 vccd1 _14882_/X sky130_fd_sc_hd__or3_2
XFILLER_130_1058 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16621_ _16622_/A _16622_/B _16622_/C vssd1 vssd1 vccd1 vccd1 _16699_/A sky130_fd_sc_hd__o21a_1
XFILLER_78_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13833_ _12845_/X _12849_/B _13838_/S vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16552_ _16455_/A _16455_/B _16456_/Y vssd1 vssd1 vccd1 vccd1 _16554_/B sky130_fd_sc_hd__a21bo_2
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ _14050_/A _14050_/B _13764_/C _13764_/D vssd1 vssd1 vccd1 vccd1 _13765_/B
+ sky130_fd_sc_hd__and4_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__xnor2_4
X_15503_ _15504_/A _15504_/B vssd1 vssd1 vccd1 vccd1 _15590_/B sky130_fd_sc_hd__nand2_2
XFILLER_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12715_ _12715_/A _12715_/B vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__nor2_1
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16483_ _16390_/Y _16395_/Y _16481_/X _16482_/Y _16917_/A vssd1 vssd1 vccd1 vccd1
+ _16483_/X sky130_fd_sc_hd__o311a_1
X_13695_ _13695_/A _13695_/B _13695_/C vssd1 vssd1 vccd1 vccd1 _13697_/A sky130_fd_sc_hd__or3_1
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ _15359_/A _15359_/B _15351_/X vssd1 vssd1 vccd1 vccd1 _15436_/B sky130_fd_sc_hd__o21ai_4
XFILLER_188_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ _12795_/A _12645_/B _12645_/C vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__a21o_1
XFILLER_169_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15365_ _15366_/B _15365_/B vssd1 vssd1 vccd1 vccd1 _15365_/X sky130_fd_sc_hd__and2b_1
XFILLER_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ _12577_/A _12577_/B vssd1 vssd1 vccd1 vccd1 _12579_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17104_ _14597_/B _14827_/Y _14826_/X _14492_/A vssd1 vssd1 vccd1 vccd1 _17104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14316_ _14316_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11528_ _11527_/A _11527_/B _11526_/Y vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__o21bai_4
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15296_ _15296_/A _15296_/B vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__xnor2_4
XFILLER_171_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17035_ _17035_/A _17035_/B _17035_/C vssd1 vssd1 vccd1 vccd1 _17035_/X sky130_fd_sc_hd__and3_1
X_14247_ _14247_/A _14330_/A vssd1 vssd1 vccd1 vccd1 _14248_/C sky130_fd_sc_hd__and2_2
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _11458_/A _11458_/B _11458_/C vssd1 vssd1 vccd1 vccd1 _11460_/C sky130_fd_sc_hd__a21oi_4
XFILLER_131_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _14090_/A _14090_/B _14088_/B vssd1 vssd1 vccd1 vccd1 _14180_/B sky130_fd_sc_hd__o21ai_4
XFILLER_152_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _12987_/X _12993_/A _13127_/X _13128_/Y vssd1 vssd1 vccd1 vccd1 _13264_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ _16819_/A _16888_/B vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _09221_/A _09221_/B _09221_/C vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__o21a_2
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09153_/A _09153_/B _09153_/C vssd1 vssd1 vccd1 vccd1 _09153_/X sky130_fd_sc_hd__or3_1
XFILLER_148_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _09084_/A _09088_/A _09084_/C vssd1 vssd1 vccd1 vccd1 _09091_/B sky130_fd_sc_hd__or3_1
XFILLER_190_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09986_ _09986_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__nor2_2
XFILLER_118_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08937_ _08937_/A _08953_/A vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__or2_2
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08868_ _08869_/A _08869_/B _08869_/C vssd1 vssd1 vccd1 vccd1 _08868_/X sky130_fd_sc_hd__a21o_2
XFILLER_123_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08799_ _11911_/B _08799_/B vssd1 vssd1 vccd1 vccd1 _08801_/C sky130_fd_sc_hd__and2_2
X_10830_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11072_/C sky130_fd_sc_hd__nand2_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10761_ _10761_/A vssd1 vssd1 vccd1 vccd1 _10761_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ _12500_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__nand2_2
X_13480_ _13595_/A _13480_/B vssd1 vssd1 vccd1 vccd1 _13482_/B sky130_fd_sc_hd__and2_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10692_ wire120/X _10667_/C _10667_/B vssd1 vssd1 vccd1 vccd1 _10692_/X sky130_fd_sc_hd__o21a_2
XFILLER_186_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ _12432_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12607_/B sky130_fd_sc_hd__and2b_1
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15150_ _15208_/C _15208_/D _14905_/C _15149_/X _15143_/A vssd1 vssd1 vccd1 vccd1
+ _15152_/B sky130_fd_sc_hd__o32a_1
XFILLER_126_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _12526_/B _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__a21o_1
X_14101_ _14188_/B _14101_/B _14102_/B vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__and3_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__xnor2_4
X_15081_ _15081_/A _16315_/C vssd1 vssd1 vccd1 vccd1 _15342_/A sky130_fd_sc_hd__nor2_2
XFILLER_126_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12293_ _12143_/A _12143_/B _12146_/A vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__o21ai_4
XFILLER_181_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14032_ _14032_/A _14032_/B vssd1 vssd1 vccd1 vccd1 _14034_/B sky130_fd_sc_hd__nor2_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11244_ _11306_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__xnor2_4
XFILLER_106_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11175_ _11176_/A _11176_/B _11176_/C vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _10254_/A _10254_/B _10392_/D _10377_/B vssd1 vssd1 vccd1 vccd1 _10128_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15983_ _15983_/A _15983_/B vssd1 vssd1 vccd1 vccd1 _15984_/B sky130_fd_sc_hd__xnor2_4
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10057_ _10057_/A _10057_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__and3_1
X_14934_ _11841_/A _15108_/A _14932_/Y _15713_/B1 _15553_/A vssd1 vssd1 vccd1 vccd1
+ _14934_/X sky130_fd_sc_hd__a2111o_1
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14865_ _16974_/A _14865_/B _16868_/A vssd1 vssd1 vccd1 vccd1 _17028_/B sky130_fd_sc_hd__and3_1
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _16938_/A _16604_/B _16758_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16604_/X
+ sky130_fd_sc_hd__and4_1
X_13816_ _13817_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _13925_/B sky130_fd_sc_hd__nand2_1
X_17584_ fanout936/X _17584_/D vssd1 vssd1 vccd1 vccd1 _17584_/Q sky130_fd_sc_hd__dfxtp_1
X_14796_ _14796_/A _14796_/B _14796_/C _14796_/D vssd1 vssd1 vccd1 vccd1 _15051_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_189_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16535_ _16536_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16537_/B sky130_fd_sc_hd__nand2_2
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13747_ _13747_/A vssd1 vssd1 vccd1 vccd1 _13748_/B sky130_fd_sc_hd__clkinv_2
XFILLER_188_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10959_ _11010_/B _10961_/B vssd1 vssd1 vccd1 vccd1 _11043_/A sky130_fd_sc_hd__nor2_2
XFILLER_73_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16466_ _16466_/A _16466_/B vssd1 vssd1 vccd1 vccd1 _16469_/A sky130_fd_sc_hd__xnor2_4
XFILLER_176_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13678_ _13678_/A _13678_/B vssd1 vssd1 vccd1 vccd1 _13680_/C sky130_fd_sc_hd__xnor2_1
X_15417_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15419_/B sky130_fd_sc_hd__xor2_4
X_12629_ _12629_/A _12629_/B vssd1 vssd1 vccd1 vccd1 _12631_/C sky130_fd_sc_hd__xor2_4
X_16397_ _12235_/C _16397_/B vssd1 vssd1 vccd1 vccd1 _16398_/B sky130_fd_sc_hd__nand2b_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15348_ _15428_/A _15428_/B vssd1 vssd1 vccd1 vccd1 _15350_/B sky130_fd_sc_hd__xnor2_4
XFILLER_184_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15279_ _15279_/A _15279_/B vssd1 vssd1 vccd1 vccd1 _15281_/B sky130_fd_sc_hd__xor2_4
XFILLER_172_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17018_ _17018_/A vssd1 vssd1 vccd1 vccd1 _17018_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ _09841_/A _09839_/Y _10366_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _09983_/A
+ sky130_fd_sc_hd__and4bb_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout607 _17510_/Q vssd1 vssd1 vccd1 vccd1 _11437_/B sky130_fd_sc_hd__buf_4
Xfanout618 _14181_/B vssd1 vssd1 vccd1 vccd1 _13745_/D sky130_fd_sc_hd__clkbuf_8
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout629 _14318_/C vssd1 vssd1 vccd1 vccd1 _14641_/C sky130_fd_sc_hd__buf_6
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_916 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ _09812_/B _09812_/C vssd1 vssd1 vccd1 vccd1 _09773_/C sky130_fd_sc_hd__nor2_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _14794_/A vssd1 vssd1 vccd1 vccd1 _08722_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ _09206_/A _09204_/Y _10062_/A _09791_/B vssd1 vssd1 vccd1 vccd1 _09375_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09136_ _09502_/A _09947_/B _09176_/B _09135_/A vssd1 vssd1 vccd1 vccd1 _09170_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09067_ _09076_/A _09055_/Y _09062_/X _09294_/A vssd1 vssd1 vccd1 vccd1 _09069_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _09969_/A _09969_/B _09969_/C vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__nor3_1
XTAP_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ _12981_/A _12981_/B vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__or2_4
XTAP_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11931_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14651_/B vssd1 vssd1 vccd1 vccd1 _14710_/B sky130_fd_sc_hd__inv_2
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _11862_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__xnor2_4
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13601_/A _13601_/B vssd1 vssd1 vccd1 vccd1 _13603_/C sky130_fd_sc_hd__or2_2
X_10813_ _10814_/B _10814_/A vssd1 vssd1 vccd1 vccd1 _11057_/A sky130_fd_sc_hd__nand2b_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14583_/A _14583_/B _14583_/C vssd1 vssd1 vccd1 vccd1 _14582_/A sky130_fd_sc_hd__a21o_1
XFILLER_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _17520_/Q _15472_/A vssd1 vssd1 vccd1 vccd1 _14876_/C sky130_fd_sc_hd__or2_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16320_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16425_/A sky130_fd_sc_hd__and2b_1
XFILLER_186_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13532_ _13532_/A _13532_/B vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__nor2_4
X_10744_ _10933_/B _10743_/C _11132_/C _10933_/A vssd1 vssd1 vccd1 vccd1 _10744_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_185_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16251_ _16251_/A _16251_/B vssd1 vssd1 vccd1 vccd1 _16252_/B sky130_fd_sc_hd__nor2_4
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13463_ _13463_/A _13463_/B vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__nor2_2
XFILLER_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10675_ _10769_/A _10675_/B vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__xor2_4
X_15202_ _14899_/X _14968_/X _15948_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15214_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12414_ _17397_/A _17395_/A _12565_/D _13094_/B vssd1 vssd1 vccd1 vccd1 _12415_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_185_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16182_ _16183_/A _16183_/B _16183_/C vssd1 vssd1 vccd1 vccd1 _16184_/A sky130_fd_sc_hd__o21a_1
XFILLER_127_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13394_ _14840_/A _17164_/A _12394_/A _13393_/Y _14667_/A vssd1 vssd1 vccd1 vccd1
+ _13394_/X sky130_fd_sc_hd__a311o_1
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15133_ _14836_/A _15094_/X _15114_/X _15132_/X vssd1 vssd1 vccd1 vccd1 _15133_/X
+ sky130_fd_sc_hd__o211a_1
X_12345_ _12175_/A _12177_/B _12175_/B vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__o21ba_2
XFILLER_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15064_ _15057_/X _15059_/Y _15061_/Y _15063_/Y _15035_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15064_/X sky130_fd_sc_hd__mux4_2
X_12276_ _12276_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _14016_/A _14015_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14015_/X sky130_fd_sc_hd__or3_1
X_11227_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__and2_4
XFILLER_96_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11158_ _11159_/A _11159_/B vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__or2_4
XFILLER_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _10236_/A _10235_/A _17469_/D _17467_/D vssd1 vssd1 vccd1 vccd1 _10112_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_67_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15966_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _15967_/B sky130_fd_sc_hd__and3_1
X_11089_ _11084_/A _11084_/C _11084_/B vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__o21a_1
XFILLER_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14917_ _15463_/A _15541_/A _15624_/A _15709_/A _10430_/A _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14918_/B sky130_fd_sc_hd__mux4_1
X_15897_ _16304_/A _15897_/B _15897_/C vssd1 vssd1 vccd1 vccd1 _15897_/X sky130_fd_sc_hd__or3_1
XFILLER_64_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14848_ _14848_/A _14848_/B _14848_/C vssd1 vssd1 vccd1 vccd1 _15314_/B sky130_fd_sc_hd__and3_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ fanout945/X _17567_/D vssd1 vssd1 vccd1 vccd1 _17567_/Q sky130_fd_sc_hd__dfxtp_1
X_14779_ _16108_/C _17119_/A vssd1 vssd1 vccd1 vccd1 _16112_/B sky130_fd_sc_hd__or2_2
XFILLER_189_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16518_ _16519_/A _16519_/B _16519_/C vssd1 vssd1 vccd1 vccd1 _16625_/A sky130_fd_sc_hd__a21oi_2
XFILLER_143_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17498_ fanout932/X _17498_/D vssd1 vssd1 vccd1 vccd1 _17498_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16449_ _16536_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16450_/B sky130_fd_sc_hd__nand2_4
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout404 _17529_/Q vssd1 vssd1 vccd1 vccd1 _09025_/C sky130_fd_sc_hd__buf_4
Xfanout415 _09407_/B vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__buf_2
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout426 _14777_/A vssd1 vssd1 vccd1 vccd1 _17397_/A sky130_fd_sc_hd__buf_6
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09823_ _09827_/A _09822_/B _09822_/A vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__o21ba_2
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout437 _16209_/C vssd1 vssd1 vccd1 vccd1 _13405_/B sky130_fd_sc_hd__buf_6
Xfanout448 _11791_/B vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__buf_6
XFILLER_87_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout459 _17523_/Q vssd1 vssd1 vccd1 vccd1 _17389_/A sky130_fd_sc_hd__buf_6
XFILLER_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09754_ _09754_/A _09758_/A _09754_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__or3_4
XFILLER_101_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09685_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__nor2_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _10459_/A _10459_/Y _10336_/Y _10353_/X vssd1 vssd1 vccd1 vccd1 _10463_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_149_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09119_ _09119_/A _09119_/B _09119_/C _09119_/D vssd1 vssd1 vccd1 vccd1 _09119_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_135_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10391_ _10391_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__xnor2_4
XFILLER_129_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12130_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12343_/B sky130_fd_sc_hd__nor2_1
XFILLER_151_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _14911_/B _12061_/B vssd1 vssd1 vccd1 vccd1 _12061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _10962_/A _10920_/B _10720_/A _10718_/Y vssd1 vssd1 vccd1 vccd1 _11013_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15820_ _15820_/A _16025_/A _15820_/C _16030_/B vssd1 vssd1 vccd1 vccd1 _15821_/D
+ sky130_fd_sc_hd__or4_1
XTAP_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15751_/A _15751_/B vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__xor2_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ _17419_/A _17417_/A _13434_/D _13321_/D vssd1 vssd1 vccd1 vccd1 _12964_/B
+ sky130_fd_sc_hd__and4_1
XTAP_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _14729_/B vssd1 vssd1 vccd1 vccd1 _14702_/Y sky130_fd_sc_hd__inv_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11914_ _11915_/A _11915_/B _12148_/B _11913_/X vssd1 vssd1 vccd1 vccd1 _11914_/X
+ sky130_fd_sc_hd__a2bb2o_2
X_15682_ _15769_/B _15682_/B _15682_/C vssd1 vssd1 vccd1 vccd1 _15690_/A sky130_fd_sc_hd__nor3_4
XFILLER_79_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12894_ _12895_/A _12895_/B vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__and2b_1
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17421_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__or2_1
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14633_/A _14633_/B vssd1 vssd1 vccd1 vccd1 _14638_/B sky130_fd_sc_hd__nand2_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11845_ _11822_/X _11844_/X _14421_/S vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__mux2_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _13908_/B _17354_/A2 _17351_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17505_/D
+ sky130_fd_sc_hd__o211a_1
X_14564_ _14565_/A _14612_/A _14564_/C vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__and3_1
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11775_/A _11773_/A _11773_/B _11774_/Y vssd1 vssd1 vccd1 vccd1 _17138_/B
+ sky130_fd_sc_hd__a31o_4
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16302_/A _16302_/B _16302_/C vssd1 vssd1 vccd1 vccd1 _16304_/C sky130_fd_sc_hd__a21oi_1
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13515_ _14756_/A1 _13513_/Y _13619_/B _13391_/Y _13394_/X vssd1 vssd1 vccd1 vccd1
+ _17587_/D sky130_fd_sc_hd__a32o_1
X_17283_ _17571_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17283_/X sky130_fd_sc_hd__and2_1
X_10727_ _10721_/X _10725_/X _10714_/X _10715_/Y vssd1 vssd1 vccd1 vccd1 _10728_/B
+ sky130_fd_sc_hd__o211ai_4
X_14495_ _14495_/A _14495_/B vssd1 vssd1 vccd1 vccd1 _14497_/C sky130_fd_sc_hd__nor2_1
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16234_ _16410_/A _16662_/D _16234_/C vssd1 vssd1 vccd1 vccd1 _16339_/A sky130_fd_sc_hd__or3_2
XFILLER_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13446_ _13329_/A _13330_/B _13444_/A _13445_/Y vssd1 vssd1 vccd1 vccd1 _13607_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_174_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10658_ _15126_/A _10755_/D _14956_/A vssd1 vssd1 vccd1 vccd1 _10658_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16165_ _16165_/A _16165_/B _16454_/A vssd1 vssd1 vccd1 vccd1 _16279_/A sky130_fd_sc_hd__and3_2
X_13377_ _13246_/A _13249_/C _13500_/A _13376_/X vssd1 vssd1 vccd1 vccd1 _13500_/B
+ sky130_fd_sc_hd__a211oi_4
X_10589_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10589_/X sky130_fd_sc_hd__and2_2
XFILLER_86_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15116_ _15116_/A _15116_/B _15796_/B vssd1 vssd1 vccd1 vccd1 _15117_/B sky130_fd_sc_hd__or3_1
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12328_ _12795_/A _12637_/C _12328_/C vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__nand3_2
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16096_ _16096_/A _16096_/B _16096_/C vssd1 vssd1 vccd1 vccd1 _16203_/A sky130_fd_sc_hd__nor3_2
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15047_ _11595_/B _15804_/A2 _15713_/B1 _14792_/B vssd1 vssd1 vccd1 vccd1 _15047_/X
+ sky130_fd_sc_hd__a22o_1
X_12259_ _12259_/A _12259_/B vssd1 vssd1 vccd1 vccd1 _12261_/B sky130_fd_sc_hd__xnor2_4
XFILLER_123_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16998_ _16880_/A _09424_/X _16743_/C _16937_/A vssd1 vssd1 vccd1 vccd1 _17000_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15949_ _16055_/A _16168_/B _16533_/B _16056_/A vssd1 vssd1 vccd1 vccd1 _15949_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09470_ _09470_/A _09470_/B _09928_/D _10309_/B vssd1 vssd1 vccd1 vccd1 _09602_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout201 _12854_/Y vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__buf_4
Xfanout212 _11800_/Y vssd1 vssd1 vccd1 vccd1 _14911_/B sky130_fd_sc_hd__buf_6
Xfanout223 _17156_/B vssd1 vssd1 vccd1 vccd1 _15309_/B sky130_fd_sc_hd__buf_4
XFILLER_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout234 _14928_/Y vssd1 vssd1 vccd1 vccd1 _16580_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout245 _16015_/A vssd1 vssd1 vccd1 vccd1 _16115_/A sky130_fd_sc_hd__buf_4
XFILLER_115_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout256 _15011_/B vssd1 vssd1 vccd1 vccd1 _16389_/A sky130_fd_sc_hd__buf_12
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__and2_1
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout267 _14939_/X vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__buf_4
Xfanout278 _12021_/A vssd1 vssd1 vccd1 vccd1 _17363_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout289 _12862_/S vssd1 vssd1 vccd1 vccd1 _15384_/S sky130_fd_sc_hd__buf_8
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09737_ _09724_/X _09725_/Y _09732_/X _09868_/A vssd1 vssd1 vccd1 vccd1 _09740_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09668_ _09668_/A _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09668_/Y sky130_fd_sc_hd__nand3_4
XFILLER_28_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09480_/A _09480_/B _09480_/C vssd1 vssd1 vccd1 vccd1 _09599_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11630_/A _14792_/B vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__nand2_4
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ _11561_/A _11561_/B _11561_/C _11561_/D vssd1 vssd1 vccd1 vccd1 _11564_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_168_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13300_ _13658_/A _17389_/A _13300_/C _13300_/D vssd1 vssd1 vccd1 vccd1 _13301_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10512_ _10970_/A _10745_/D _10415_/A _10413_/Y vssd1 vssd1 vccd1 vccd1 _10513_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14280_ _14121_/X _14281_/B _14279_/Y _14204_/A vssd1 vssd1 vccd1 vccd1 _14280_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11492_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11493_/C sky130_fd_sc_hd__xnor2_4
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _13232_/A _13232_/B vssd1 vssd1 vccd1 vccd1 _13361_/A sky130_fd_sc_hd__and2b_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10443_ _10407_/Y _10442_/Y _10319_/Y _10354_/X vssd1 vssd1 vccd1 vccd1 _10459_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13162_ _13295_/B _13162_/B vssd1 vssd1 vccd1 vccd1 _13165_/C sky130_fd_sc_hd__nand2_2
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10374_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10375_/B sky130_fd_sc_hd__or3_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _12113_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__xnor2_1
XFILLER_123_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13093_ _13093_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__nor2_1
X_16921_ _16921_/A _16921_/B vssd1 vssd1 vccd1 vccd1 _16922_/B sky130_fd_sc_hd__xnor2_1
X_12044_ _12700_/D _12044_/B vssd1 vssd1 vccd1 vccd1 _12044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16852_ _16786_/A _16853_/A _16786_/B vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_172_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout790 _17490_/Q vssd1 vssd1 vccd1 vccd1 _13321_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15803_ _15801_/B _15899_/A2 _16008_/B1 _15811_/A _16008_/C1 vssd1 vssd1 vccd1 vccd1
+ _15803_/X sky130_fd_sc_hd__a221o_1
X_16783_ _16784_/A _16784_/B _16784_/C vssd1 vssd1 vccd1 vccd1 _16850_/A sky130_fd_sc_hd__a21oi_2
X_13995_ _17409_/A _14545_/D vssd1 vssd1 vccd1 vccd1 _13997_/B sky130_fd_sc_hd__and2_1
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15734_ _15734_/A _15734_/B _16039_/B _16150_/B vssd1 vssd1 vccd1 vccd1 _15735_/B
+ sky130_fd_sc_hd__or4_4
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12946_ _12946_/A _13085_/B vssd1 vssd1 vccd1 vccd1 _12947_/C sky130_fd_sc_hd__nor2_1
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _15666_/A _15666_/B vssd1 vssd1 vccd1 vccd1 _15665_/Y sky130_fd_sc_hd__nand2_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _17397_/A _17395_/A _14153_/C _14215_/B vssd1 vssd1 vccd1 vccd1 _13040_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14658_/A _14616_/B vssd1 vssd1 vccd1 vccd1 _14618_/B sky130_fd_sc_hd__nor2_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ input48/X _17422_/A2 _17403_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17530_/D
+ sky130_fd_sc_hd__o211a_1
X_11828_ _12618_/D _12463_/D _12060_/S vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__mux2_1
X_15596_ _16281_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _15598_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ input46/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17335_/X sky130_fd_sc_hd__or3_1
X_14547_ _14548_/A _14601_/A _14548_/C vssd1 vssd1 vccd1 vccd1 _14549_/A sky130_fd_sc_hd__o21a_1
XFILLER_147_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ _11759_/A _11762_/A vssd1 vssd1 vccd1 vccd1 _16641_/A sky130_fd_sc_hd__xor2_4
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17266_ _17456_/Q _17266_/A2 _17264_/X _17265_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17456_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14478_ _14479_/A _14479_/B vssd1 vssd1 vccd1 vccd1 _14478_/X sky130_fd_sc_hd__or2_1
XFILLER_174_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16217_ _14859_/B _16115_/B _16216_/Y vssd1 vssd1 vccd1 vccd1 _16221_/B sky130_fd_sc_hd__o21a_1
X_13429_ _13428_/A _13428_/B _13427_/X vssd1 vssd1 vccd1 vccd1 _13430_/B sky130_fd_sc_hd__o21bai_1
XFILLER_128_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17197_ _17198_/C _17185_/X _17231_/A2 _17575_/Q _17231_/B1 vssd1 vssd1 vccd1 vccd1
+ _17197_/X sky130_fd_sc_hd__a221o_1
XFILLER_161_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ _16032_/A _16034_/B _16032_/B vssd1 vssd1 vccd1 vccd1 _16155_/A sky130_fd_sc_hd__o21ba_4
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _16080_/A _16080_/B _16080_/C vssd1 vssd1 vccd1 vccd1 _16081_/A sky130_fd_sc_hd__o21ai_4
X_08970_ _09780_/A _08968_/B _12700_/C vssd1 vssd1 vccd1 vccd1 _08971_/C sky130_fd_sc_hd__a21oi_4
XFILLER_130_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput1 buttons vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09522_ _09522_/A _09522_/B _09634_/A vssd1 vssd1 vccd1 vccd1 _09523_/B sky130_fd_sc_hd__nor3_2
XFILLER_37_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09453_ _09440_/X _09441_/Y _09448_/X _09579_/A vssd1 vssd1 vccd1 vccd1 _09455_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09384_ _09385_/B _09385_/A vssd1 vssd1 vccd1 vccd1 _09384_/X sky130_fd_sc_hd__and2b_1
XFILLER_40_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1001 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10090_ _10090_/A _10101_/A vssd1 vssd1 vccd1 vccd1 _10091_/C sky130_fd_sc_hd__nor2_2
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ _12800_/A _12950_/B vssd1 vssd1 vccd1 vccd1 _12801_/B sky130_fd_sc_hd__nand2_2
X_13780_ _13676_/A _13678_/B _13676_/B vssd1 vssd1 vccd1 vccd1 _13781_/B sky130_fd_sc_hd__o21ba_1
XFILLER_56_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ _15126_/A _10899_/D _10657_/C vssd1 vssd1 vccd1 vccd1 _10992_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12577_/A _12579_/B _12577_/B vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__o21ba_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15450_ _15450_/A _15796_/B _15396_/A vssd1 vssd1 vccd1 vccd1 _15453_/B sky130_fd_sc_hd__or3b_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12662_ _12662_/A _12662_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__nor3_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14401_ _14401_/A vssd1 vssd1 vccd1 vccd1 _14466_/B sky130_fd_sc_hd__inv_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11613_/A _11646_/A vssd1 vssd1 vccd1 vccd1 _11614_/C sky130_fd_sc_hd__nand2_1
X_15381_ _15381_/A _15381_/B vssd1 vssd1 vccd1 vccd1 _15381_/Y sky130_fd_sc_hd__nor2_1
X_12593_ _12593_/A _12775_/A vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__or2_2
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17120_ _17119_/A _17081_/A _17038_/B _17038_/C _17086_/A vssd1 vssd1 vccd1 vccd1
+ _17121_/B sky130_fd_sc_hd__o41a_1
X_14332_ _14333_/A _14333_/B vssd1 vssd1 vccd1 vccd1 _14332_/X sky130_fd_sc_hd__or2_4
XFILLER_168_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11544_ _11460_/B _11460_/C _11460_/A vssd1 vssd1 vccd1 vccd1 _11544_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_183_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17051_ _17052_/A _17052_/B _17050_/X vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__o21ba_1
X_14263_ _14265_/A _14265_/B vssd1 vssd1 vccd1 vccd1 _14266_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ _11475_/A _11475_/B _11475_/C vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__and3_4
XFILLER_13_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16002_ _15891_/X _15892_/Y _15890_/X vssd1 vssd1 vccd1 vccd1 _16004_/B sky130_fd_sc_hd__a21boi_2
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__o21ai_2
X_10426_ _10427_/B _10427_/C _10427_/A vssd1 vssd1 vccd1 vccd1 _10437_/A sky130_fd_sc_hd__a21o_1
X_14194_ _14194_/A _14195_/B _14102_/B vssd1 vssd1 vccd1 vccd1 _14270_/B sky130_fd_sc_hd__or3b_2
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145_ _17371_/A _13145_/B vssd1 vssd1 vccd1 vccd1 _13145_/Y sky130_fd_sc_hd__nor2_1
X_10357_ _10262_/A _10262_/C _10262_/B vssd1 vssd1 vccd1 vccd1 _10357_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _12933_/B _12935_/A _13074_/X _13075_/Y vssd1 vssd1 vccd1 vccd1 _13121_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_140_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10288_ _10288_/A _10296_/A _10288_/C vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__or3_1
X_16904_ _16905_/A _16905_/B vssd1 vssd1 vccd1 vccd1 _17008_/A sky130_fd_sc_hd__nand2_1
X_12027_ _12024_/Y _12026_/Y _15038_/A vssd1 vssd1 vccd1 vccd1 _12027_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16835_ _16835_/A _16835_/B _16835_/C vssd1 vssd1 vccd1 vccd1 _16836_/B sky130_fd_sc_hd__nor3_1
XFILLER_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _13978_/A _13978_/B vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__nor2_2
X_16766_ _16767_/A _16767_/B vssd1 vssd1 vccd1 vccd1 _16768_/A sky130_fd_sc_hd__and2_1
XFILLER_53_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15717_ _14924_/A _12401_/A _13273_/X _15716_/X vssd1 vssd1 vccd1 vccd1 _15717_/Y
+ sky130_fd_sc_hd__o31ai_1
X_12929_ _13117_/A _12929_/B vssd1 vssd1 vccd1 vccd1 _12931_/B sky130_fd_sc_hd__and2_1
X_16697_ _16697_/A _16697_/B _16697_/C vssd1 vssd1 vccd1 vccd1 _16698_/B sky130_fd_sc_hd__or3_1
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15648_ _15648_/A _15648_/B vssd1 vssd1 vccd1 vccd1 _15651_/A sky130_fd_sc_hd__xnor2_4
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15579_ _16056_/A _15774_/B _15578_/B vssd1 vssd1 vccd1 vccd1 _15580_/B sky130_fd_sc_hd__a21oi_2
XFILLER_187_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17318_ _13067_/D _17322_/A2 _17317_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17488_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17249_ _17592_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08953_ _08953_/A _08959_/A _08953_/C vssd1 vssd1 vccd1 vccd1 _08962_/B sky130_fd_sc_hd__or3_1
XFILLER_103_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08884_ _11026_/A _10647_/D vssd1 vssd1 vccd1 vccd1 _16315_/A sky130_fd_sc_hd__nand2_8
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09505_ _09786_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__and2_4
XFILLER_53_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09577_/A vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__nand2_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09370_/B _09367_/B vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__and2_2
XFILLER_184_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09298_ _09298_/A _09298_/B vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__nor2_1
XANTENNA_50 _15101_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_61 _15872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_72 i_wb_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_83 _17441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_94 fanout757/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ _11261_/A _11259_/Y _11260_/C _11563_/D vssd1 vssd1 vccd1 vccd1 _11304_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_192_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10211_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10211_/Y sky130_fd_sc_hd__nand2_1
X_11191_ _11222_/A _11190_/C _11190_/A vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__o21a_2
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _10392_/A _10738_/D vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__nand2_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__xor2_2
XFILLER_82_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14950_ _15038_/A _14949_/Y _14948_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14950_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_102_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13901_ _13900_/B _13901_/B vssd1 vssd1 vccd1 vccd1 _13902_/B sky130_fd_sc_hd__nand2b_4
XFILLER_130_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14881_ _14876_/X _14880_/X _15143_/A vssd1 vssd1 vccd1 vccd1 _14881_/X sky130_fd_sc_hd__a21o_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16620_ _16620_/A _16774_/A vssd1 vssd1 vccd1 vccd1 _16622_/C sky130_fd_sc_hd__and2_1
XFILLER_46_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13832_ _14839_/A _13832_/B vssd1 vssd1 vccd1 vccd1 _13832_/Y sky130_fd_sc_hd__nor2_1
X_16551_ _16636_/A _16551_/B vssd1 vssd1 vccd1 vccd1 _16554_/A sky130_fd_sc_hd__nand2_2
X_13763_ _14050_/B _13764_/C _13764_/D _14050_/A vssd1 vssd1 vccd1 vccd1 _13765_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10975_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _11024_/B sky130_fd_sc_hd__and2_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15594_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15504_/B sky130_fd_sc_hd__nor2_4
X_12714_ _17403_/A _17399_/A _13564_/C _13450_/D vssd1 vssd1 vccd1 vccd1 _12715_/B
+ sky130_fd_sc_hd__and4_1
X_16482_ _16390_/Y _16395_/Y _16481_/X vssd1 vssd1 vccd1 vccd1 _16482_/Y sky130_fd_sc_hd__o21ai_2
X_13694_ _13694_/A _13793_/B vssd1 vssd1 vccd1 vccd1 _13695_/C sky130_fd_sc_hd__nor2_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15433_ _15433_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15436_/A sky130_fd_sc_hd__xor2_4
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12645_ _12795_/A _12645_/B _12645_/C vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__nand3_4
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15364_ _15296_/A _15296_/B _15294_/Y vssd1 vssd1 vccd1 vccd1 _15365_/B sky130_fd_sc_hd__o21ai_1
X_12576_ _17391_/A _17389_/A _12576_/C _12576_/D vssd1 vssd1 vccd1 vccd1 _12577_/B
+ sky130_fd_sc_hd__and4_1
X_14315_ _14315_/A _14315_/B vssd1 vssd1 vccd1 vccd1 _14316_/B sky130_fd_sc_hd__nand2_1
X_17103_ _17156_/B _17103_/B _17102_/X vssd1 vssd1 vccd1 vccd1 _17103_/X sky130_fd_sc_hd__or3b_1
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11527_ _11527_/A _11527_/B _11526_/Y vssd1 vssd1 vccd1 vccd1 _11534_/B sky130_fd_sc_hd__or3b_4
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15295_ _15295_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _15296_/B sky130_fd_sc_hd__xor2_4
XFILLER_116_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17034_ _17021_/Y _17022_/X _17024_/X _17169_/A1 vssd1 vssd1 vccd1 vccd1 _17035_/C
+ sky130_fd_sc_hd__o22a_1
X_14246_ _14245_/A _14245_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14330_/A sky130_fd_sc_hd__o21ai_4
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11458_ _11458_/A _11458_/B _11458_/C vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__and3_2
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _10402_/A _10402_/Y _10408_/Y _10315_/X vssd1 vssd1 vccd1 vccd1 _10453_/A
+ sky130_fd_sc_hd__a211o_4
X_14177_ _14177_/A _14177_/B vssd1 vssd1 vccd1 vccd1 _14180_/A sky130_fd_sc_hd__xor2_4
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11389_ _11629_/A _11480_/C vssd1 vssd1 vccd1 vccd1 _11389_/X sky130_fd_sc_hd__and2_1
XFILLER_139_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13258_/A _13125_/X _12980_/X _12984_/A vssd1 vssd1 vccd1 vccd1 _13128_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13060_/A _13060_/B vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__and2b_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16818_ _16818_/A _16818_/B vssd1 vssd1 vccd1 vccd1 _16888_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16749_ _16883_/C _16749_/B vssd1 vssd1 vccd1 vccd1 _16750_/B sky130_fd_sc_hd__xnor2_2
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _09221_/A _09221_/B _09221_/C vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__nor3_2
XFILLER_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09152_ _09152_/A vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09083_ _09084_/A _09084_/C vssd1 vssd1 vccd1 vccd1 _09088_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput70 reset vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_4
XFILLER_174_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09985_ _10115_/A _10241_/B _10491_/B _10490_/C vssd1 vssd1 vccd1 vccd1 _09986_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08936_ _11932_/A _12595_/C _08936_/C _08936_/D vssd1 vssd1 vccd1 vccd1 _08953_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_190_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08867_ _08867_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08869_/C sky130_fd_sc_hd__or2_2
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08798_ _08798_/A _08821_/A _08798_/C vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__or3_1
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10760_ _10760_/A _10760_/B _10760_/C vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__and3_2
XFILLER_73_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ _09434_/B _09434_/C _09434_/A vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__a21o_2
X_10691_ _10678_/A _10677_/C _10677_/B vssd1 vssd1 vccd1 vccd1 _10691_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12430_ _12607_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__nor2_4
XFILLER_185_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _12526_/B _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__nand3_2
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14100_ _14011_/A _14115_/B _14010_/B _13990_/B _13990_/A vssd1 vssd1 vccd1 vccd1
+ _14102_/B sky130_fd_sc_hd__a32o_2
XFILLER_148_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11312_ _11311_/A _11311_/C _11311_/B vssd1 vssd1 vccd1 vccd1 _11312_/Y sky130_fd_sc_hd__o21ai_4
X_15080_ _15278_/A _15647_/A vssd1 vssd1 vccd1 vccd1 _15157_/A sky130_fd_sc_hd__nand2_4
X_12292_ _12289_/Y _12290_/X _12122_/A _12122_/Y vssd1 vssd1 vccd1 vccd1 _12312_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14031_ _14029_/Y _14031_/B vssd1 vssd1 vccd1 vccd1 _14122_/B sky130_fd_sc_hd__nand2b_1
X_11243_ _11306_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__and2_2
XFILLER_153_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11176_/C sky130_fd_sc_hd__xor2_4
XFILLER_84_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10125_ _10125_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__xnor2_4
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15982_ _16281_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _15983_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10056_ _10029_/A _10029_/B _10029_/C vssd1 vssd1 vccd1 vccd1 _10057_/C sky130_fd_sc_hd__o21ai_4
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14933_ _14933_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14933_/Y sky130_fd_sc_hd__nor2_4
XFILLER_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14864_ _14864_/A _14864_/B vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__and2_2
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16603_ _16758_/B _16809_/C _16165_/B _16604_/B vssd1 vssd1 vccd1 vccd1 _16603_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13815_ _13925_/A _13815_/B vssd1 vssd1 vccd1 vccd1 _13817_/B sky130_fd_sc_hd__and2_2
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14795_ _14794_/A _14794_/B _15008_/B _11651_/A vssd1 vssd1 vccd1 vccd1 _14796_/D
+ sky130_fd_sc_hd__a22o_1
X_17583_ fanout936/X _17583_/D vssd1 vssd1 vccd1 vccd1 _17583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13746_ _13746_/A _13858_/A vssd1 vssd1 vccd1 vccd1 _13747_/A sky130_fd_sc_hd__or2_1
X_16534_ _16534_/A _16622_/A vssd1 vssd1 vccd1 vccd1 _16537_/A sky130_fd_sc_hd__nor2_4
XFILLER_188_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _11005_/A _10957_/D _10955_/Y _10957_/B vssd1 vssd1 vccd1 vccd1 _10961_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16465_ _16466_/A _16466_/B vssd1 vssd1 vccd1 vccd1 _16557_/B sky130_fd_sc_hd__nor2_1
X_13677_ _14226_/A _14141_/D vssd1 vssd1 vccd1 vccd1 _13678_/B sky130_fd_sc_hd__nand2_1
XFILLER_189_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10889_ _10899_/C _11132_/C _11131_/B vssd1 vssd1 vccd1 vccd1 _10891_/C sky130_fd_sc_hd__and3_1
XFILLER_176_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15416_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15416_/Y sky130_fd_sc_hd__nor2_1
X_12628_ _12629_/B _12629_/A vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__nand2b_1
X_16396_ _16396_/A _16396_/B vssd1 vssd1 vccd1 vccd1 _16396_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15347_ _15428_/A _15428_/B vssd1 vssd1 vccd1 vccd1 _15429_/A sky130_fd_sc_hd__nand2_2
XFILLER_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _12235_/C _12869_/C _12557_/X vssd1 vssd1 vccd1 vccd1 _12560_/B sky130_fd_sc_hd__a21bo_2
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15278_ _15278_/A _15397_/A vssd1 vssd1 vccd1 vccd1 _15279_/B sky130_fd_sc_hd__nand2_2
XFILLER_176_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14229_ _14229_/A _14229_/B _14229_/C vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__nor3_1
X_17017_ _14766_/A _17134_/C _17028_/A vssd1 vssd1 vccd1 vccd1 _17018_/A sky130_fd_sc_hd__a21bo_1
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _12442_/B vssd1 vssd1 vccd1 vccd1 _12592_/C sky130_fd_sc_hd__buf_8
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout619 _13300_/C vssd1 vssd1 vccd1 vccd1 _14181_/B sky130_fd_sc_hd__buf_6
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09770_ _09812_/C vssd1 vssd1 vccd1 vccd1 _09770_/Y sky130_fd_sc_hd__clkinv_2
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _12845_/S vssd1 vssd1 vccd1 vccd1 _08721_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09204_ _09637_/B _09937_/B _09803_/B _09942_/A vssd1 vssd1 vccd1 vccd1 _09204_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_50_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__nor2_2
XFILLER_120_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__and2_2
XFILLER_136_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _09968_/A _09968_/B _09970_/A vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__or3_4
XTAP_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _17375_/A _12734_/D vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__nand2_1
XTAP_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _14789_/A _10171_/B _10543_/B _10657_/B vssd1 vssd1 vccd1 vccd1 _10034_/A
+ sky130_fd_sc_hd__and4_2
XTAP_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ _17373_/A _11930_/B _12752_/B _12270_/C vssd1 vssd1 vccd1 vccd1 _11931_/B
+ sky130_fd_sc_hd__and4_1
XTAP_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _12237_/A _12068_/D vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__nand2_4
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13601_/B sky130_fd_sc_hd__and2_1
XFILLER_26_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _10812_/A _10823_/A vssd1 vssd1 vccd1 vccd1 _10814_/B sky130_fd_sc_hd__nor2_2
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14627_/B _14580_/B vssd1 vssd1 vccd1 vccd1 _14583_/C sky130_fd_sc_hd__or2_1
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _16809_/A _16136_/A _15262_/A vssd1 vssd1 vccd1 vccd1 _14888_/C sky130_fd_sc_hd__or3_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _13641_/A _13745_/B _13948_/D _13844_/D vssd1 vssd1 vccd1 vccd1 _13532_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10743_ _10933_/A _10933_/B _10743_/C _11132_/C vssd1 vssd1 vccd1 vccd1 _10746_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_186_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16250_ _16250_/A _16250_/B _16250_/C vssd1 vssd1 vccd1 vccd1 _16251_/B sky130_fd_sc_hd__nor3_2
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _13462_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13463_/B sky130_fd_sc_hd__and3_1
XFILLER_186_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10674_ _10769_/A _10675_/B vssd1 vssd1 vccd1 vccd1 _10674_/Y sky130_fd_sc_hd__nor2_1
XFILLER_167_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _15726_/A _16536_/A vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__nand2_4
XFILLER_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12413_ _17395_/A _12565_/D _13094_/B _17397_/A vssd1 vssd1 vccd1 vccd1 _12415_/A
+ sky130_fd_sc_hd__a22oi_4
X_16181_ _16181_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _16183_/C sky130_fd_sc_hd__xnor2_2
XFILLER_159_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13393_ _14666_/S _13393_/B vssd1 vssd1 vccd1 vccd1 _13393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ _15119_/Y _15120_/X _15106_/Y vssd1 vssd1 vccd1 vccd1 _15132_/X sky130_fd_sc_hd__o21a_1
XFILLER_153_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ _12344_/A _12344_/B vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15063_ _15131_/A _15063_/B vssd1 vssd1 vccd1 vccd1 _15063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ _12275_/A _17383_/A _12578_/B _12576_/C vssd1 vssd1 vccd1 vccd1 _12276_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14014_ _14015_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14016_/B sky130_fd_sc_hd__nor2_1
X_11226_ _11195_/A _11194_/B _11194_/A vssd1 vssd1 vccd1 vccd1 _11228_/B sky130_fd_sc_hd__o21bai_4
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11157_ _11157_/A _11157_/B vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__and2_4
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _10113_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__nor2_2
X_15965_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__a21oi_2
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__xnor2_4
XFILLER_64_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10039_ _10039_/A _10151_/A vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__nor2_2
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14916_ _14958_/A _14913_/Y _14915_/Y _14912_/Y vssd1 vssd1 vccd1 vccd1 _14916_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15896_ _16933_/A _15895_/B _15895_/C vssd1 vssd1 vccd1 vccd1 _15897_/C sky130_fd_sc_hd__a21oi_1
XFILLER_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14847_ _15116_/B _15110_/B vssd1 vssd1 vccd1 vccd1 _14848_/C sky130_fd_sc_hd__and2_1
XFILLER_17_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17566_ fanout945/X _17566_/D vssd1 vssd1 vccd1 vccd1 _17566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14778_ _16209_/C _14859_/B vssd1 vssd1 vccd1 vccd1 _14778_/X sky130_fd_sc_hd__or2_2
X_16517_ _16517_/A _16517_/B vssd1 vssd1 vccd1 vccd1 _16519_/C sky130_fd_sc_hd__xnor2_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13729_ _13514_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__nand2b_2
XFILLER_189_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17497_ fanout932/X _17497_/D vssd1 vssd1 vccd1 vccd1 _17497_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16448_ _16533_/A _16165_/B _16533_/C _16447_/Y vssd1 vssd1 vccd1 vccd1 _16450_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16379_ _16285_/A _16285_/B _16287_/Y vssd1 vssd1 vccd1 vccd1 _16381_/B sky130_fd_sc_hd__a21bo_2
XFILLER_145_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout405 _17529_/Q vssd1 vssd1 vccd1 vccd1 _12237_/A sky130_fd_sc_hd__buf_4
Xfanout416 _17528_/Q vssd1 vssd1 vccd1 vccd1 _09407_/B sky130_fd_sc_hd__clkbuf_4
Xfanout427 _13641_/A vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__buf_6
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout438 _17526_/Q vssd1 vssd1 vccd1 vccd1 _16209_/C sky130_fd_sc_hd__buf_6
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout449 _17391_/A vssd1 vssd1 vccd1 vccd1 _13658_/A sky130_fd_sc_hd__buf_6
XFILLER_63_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09753_ _09754_/A _09754_/C vssd1 vssd1 vccd1 vccd1 _09758_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _09626_/A _09629_/B _09626_/C vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _09119_/A _09119_/D vssd1 vssd1 vccd1 vccd1 _09257_/B sky130_fd_sc_hd__nand2_2
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10390_ _10390_/A _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__nand3_4
XFILLER_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _09050_/A _09049_/B _09049_/C vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__nand3_4
XFILLER_191_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12060_ _17302_/A1 _10321_/C _12060_/S vssd1 vssd1 vccd1 vccd1 _12061_/B sky130_fd_sc_hd__mux2_1
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _11025_/B _11025_/A vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__nand2b_4
XFILLER_89_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _16165_/A _16352_/B _15751_/A vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__and3_1
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12962_ _17417_/A _13434_/D _13321_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _12964_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _14701_/A _14701_/B vssd1 vssd1 vccd1 vccd1 _14729_/B sky130_fd_sc_hd__nor2_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _12148_/A _11911_/Y _08863_/X _08867_/A vssd1 vssd1 vccd1 vccd1 _11913_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_46_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15588_/A _15588_/B _15563_/Y vssd1 vssd1 vccd1 vccd1 _15682_/C sky130_fd_sc_hd__a21oi_4
X_12893_ _13043_/B _12893_/B vssd1 vssd1 vccd1 vccd1 _12895_/B sky130_fd_sc_hd__nor2_2
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ input56/X _17422_/A2 _17419_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17538_/D
+ sky130_fd_sc_hd__o211a_1
X_14632_ _14633_/A _14633_/B vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__or2_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _11827_/X _11832_/X _11838_/X _11843_/X _12865_/S _17369_/A vssd1 vssd1 vccd1
+ vccd1 _11844_/X sky130_fd_sc_hd__mux4_2
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14612_/A _14564_/C vssd1 vssd1 vccd1 vccd1 _14565_/B sky130_fd_sc_hd__and2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ input55/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17351_/X sky130_fd_sc_hd__or3_1
XFILLER_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11775_ _11775_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11775_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16302_/A _16302_/B _16302_/C vssd1 vssd1 vccd1 vccd1 _16304_/B sky130_fd_sc_hd__and3_1
X_10726_ _10714_/X _10715_/Y _10721_/X _10725_/X vssd1 vssd1 vccd1 vccd1 _10728_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_41_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13514_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13619_/B sky130_fd_sc_hd__or2_1
X_14494_ _16965_/C _14708_/D _14493_/C vssd1 vssd1 vccd1 vccd1 _14495_/B sky130_fd_sc_hd__a21oi_1
X_17282_ _17603_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__a21o_1
XFILLER_41_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16233_ _11791_/C _16317_/B _15209_/Y _16743_/C vssd1 vssd1 vccd1 vccd1 _16235_/A
+ sky130_fd_sc_hd__a22o_1
X_13445_ _13443_/A _13443_/B _13443_/C vssd1 vssd1 vccd1 vccd1 _13445_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ _15126_/A _10657_/B _10657_/C vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__and3_2
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16164_ _16165_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13376_ _13494_/B _13374_/X _13249_/A _13249_/Y vssd1 vssd1 vccd1 vccd1 _13376_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_186_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10588_ _10500_/Y _10519_/C _10519_/B vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__o21a_1
XFILLER_115_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12327_ _12327_/A _12498_/A vssd1 vssd1 vccd1 vccd1 _12328_/C sky130_fd_sc_hd__and2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15115_ _15116_/A _15796_/B _15116_/B vssd1 vssd1 vccd1 vccd1 _15117_/A sky130_fd_sc_hd__o21ai_2
XFILLER_181_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16095_ _16095_/A _16095_/B vssd1 vssd1 vccd1 vccd1 _16096_/C sky130_fd_sc_hd__xnor2_4
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15046_ _15008_/A _15008_/B _14792_/B vssd1 vssd1 vccd1 vccd1 _15046_/Y sky130_fd_sc_hd__a21oi_1
X_12258_ _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__nand2_4
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11209_ _11168_/A _11168_/Y _11719_/A _11208_/Y vssd1 vssd1 vccd1 vccd1 _11719_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_141_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12189_ _12189_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12190_/B sky130_fd_sc_hd__nand2_2
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16997_ _16997_/A _17052_/A vssd1 vssd1 vccd1 vccd1 _17000_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15948_ _15948_/A _16827_/C vssd1 vssd1 vccd1 vccd1 _16361_/A sky130_fd_sc_hd__or2_4
XFILLER_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15879_ _15773_/B _15775_/B _15773_/A vssd1 vssd1 vccd1 vccd1 _15881_/B sky130_fd_sc_hd__o21ba_1
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17549_ fanout934/X _17549_/D vssd1 vssd1 vccd1 vccd1 _17549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout202 _12401_/A vssd1 vssd1 vccd1 vccd1 _15457_/B sky130_fd_sc_hd__buf_4
XFILLER_132_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout213 _17362_/C vssd1 vssd1 vccd1 vccd1 _17327_/B sky130_fd_sc_hd__clkbuf_4
Xfanout224 _14938_/X vssd1 vssd1 vccd1 vccd1 _17156_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_141_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout235 _14928_/Y vssd1 vssd1 vccd1 vccd1 _15899_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout246 _14844_/X vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__buf_2
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09805_ _09805_/A _09805_/B _09939_/A vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__or3_1
Xfanout257 _17429_/C vssd1 vssd1 vccd1 vccd1 _17327_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout268 _14939_/X vssd1 vssd1 vccd1 vccd1 _16108_/B sky130_fd_sc_hd__buf_2
Xfanout279 _12054_/A vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09736_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__and2_2
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ _09628_/A _09628_/B _09628_/C vssd1 vssd1 vccd1 vccd1 _09668_/C sky130_fd_sc_hd__o21ai_4
XFILLER_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09624_/B _09624_/C _09624_/A vssd1 vssd1 vccd1 vccd1 _09627_/A sky130_fd_sc_hd__o21a_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ _11565_/A _11565_/B vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__xnor2_2
XFILLER_183_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _11444_/Y _11466_/X _11487_/A _11527_/A vssd1 vssd1 vccd1 vccd1 _11493_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_137_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13230_ _13230_/A _13230_/B vssd1 vssd1 vccd1 vccd1 _13232_/B sky130_fd_sc_hd__xnor2_2
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10442_ _10473_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10442_/Y sky130_fd_sc_hd__nor2_2
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13161_ _13161_/A _13161_/B vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__or2_1
XFILLER_164_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__o21ai_4
XFILLER_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ _12113_/B _12113_/A vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__and2b_2
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ _13092_/A _13092_/B _13092_/C vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__and3_1
XFILLER_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16920_ _10784_/A _10784_/B _11766_/X vssd1 vssd1 vccd1 vccd1 _16921_/B sky130_fd_sc_hd__o21ai_1
X_12043_ _12770_/D _12618_/D _12060_/S vssd1 vssd1 vccd1 vccd1 _12044_/B sky130_fd_sc_hd__mux2_1
XFILLER_137_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16851_ _16851_/A _16851_/B vssd1 vssd1 vccd1 vccd1 _16931_/A sky130_fd_sc_hd__nand2_1
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout780 _09030_/D vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__buf_6
Xfanout791 _17489_/Q vssd1 vssd1 vccd1 vccd1 _12158_/C sky130_fd_sc_hd__clkbuf_16
XFILLER_93_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15802_ _15802_/A _15802_/B vssd1 vssd1 vccd1 vccd1 _15802_/Y sky130_fd_sc_hd__xnor2_1
X_16782_ _16846_/B _16782_/B vssd1 vssd1 vccd1 vccd1 _16784_/C sky130_fd_sc_hd__or2_1
X_13994_ _16864_/A _16918_/A _13991_/X vssd1 vssd1 vccd1 vccd1 _13997_/A sky130_fd_sc_hd__o21a_1
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15733_ _15647_/A _16604_/B _16758_/B _16226_/B vssd1 vssd1 vccd1 vccd1 _15735_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12945_/A _13085_/A _12945_/C vssd1 vssd1 vccd1 vccd1 _13085_/B sky130_fd_sc_hd__nor3_2
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15664_ _16410_/A _16446_/A vssd1 vssd1 vccd1 vccd1 _15666_/B sky130_fd_sc_hd__nor2_8
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _17395_/A _14153_/C _14215_/B _17397_/A vssd1 vssd1 vccd1 vccd1 _12878_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17403_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17403_/X sky130_fd_sc_hd__or2_1
X_14615_ _14614_/B _14615_/B vssd1 vssd1 vccd1 vccd1 _14616_/B sky130_fd_sc_hd__and2b_1
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _11824_/Y _11826_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _15595_/A _15595_/B vssd1 vssd1 vccd1 vccd1 _15598_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _12950_/B _17360_/A2 _17333_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17496_/D
+ sky130_fd_sc_hd__o211a_1
X_14546_ _14676_/A _14641_/D vssd1 vssd1 vccd1 vccd1 _14548_/C sky130_fd_sc_hd__nand2_1
X_11758_ _11758_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__nor2_4
XFILLER_18_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10709_ _10709_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__xor2_4
X_17265_ _17565_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17265_/X sky130_fd_sc_hd__and2_1
X_14477_ _14533_/A _14419_/B _14414_/A vssd1 vssd1 vccd1 vccd1 _14479_/B sky130_fd_sc_hd__a21oi_1
XFILLER_159_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11689_ _15302_/A _15302_/B vssd1 vssd1 vccd1 vccd1 _15303_/A sky130_fd_sc_hd__nand2_1
X_16216_ _14859_/B _16115_/B _16652_/A vssd1 vssd1 vccd1 vccd1 _16216_/Y sky130_fd_sc_hd__a21oi_1
X_13428_ _13428_/A _13428_/B _13427_/X vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__or3b_4
XFILLER_128_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17196_ input29/X _17196_/B _17196_/C vssd1 vssd1 vccd1 vccd1 _17196_/X sky130_fd_sc_hd__or3_4
XFILLER_128_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16147_ _16040_/A _16040_/B _16043_/A vssd1 vssd1 vccd1 vccd1 _16157_/A sky130_fd_sc_hd__a21bo_4
XFILLER_154_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13359_ _13360_/B _13360_/A vssd1 vssd1 vccd1 vccd1 _13477_/B sky130_fd_sc_hd__and2b_1
XFILLER_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16078_ _16183_/B _16078_/B vssd1 vssd1 vccd1 vccd1 _16080_/C sky130_fd_sc_hd__nor2_2
XFILLER_143_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15029_ _15820_/A _15687_/A _15028_/A vssd1 vssd1 vccd1 vccd1 _15030_/D sky130_fd_sc_hd__o21ai_2
XFILLER_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 clk vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_16
XFILLER_110_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09522_/B _09634_/A _09522_/A vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__o21a_1
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__and2_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09383_ _09383_/A _09511_/A vssd1 vssd1 vccd1 vccd1 _09385_/B sky130_fd_sc_hd__nor2_4
XFILLER_178_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1013 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09719_ _09720_/A _09719_/B _09719_/C vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__nand3_1
X_10991_ _15126_/A _11841_/B _10991_/C vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__and3_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12730_ _12730_/A _12730_/B _12730_/C vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__nand3_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12661_ _12662_/A _12662_/B _12662_/C vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__o21a_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _14400_/A _14466_/A _14400_/C vssd1 vssd1 vccd1 vccd1 _14401_/A sky130_fd_sc_hd__and3_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11612_ _11613_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__nand3_1
XFILLER_187_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15102_/Y _15123_/Y _15125_/Y _15131_/Y _15130_/S _15116_/A vssd1 vssd1 vccd1
+ vccd1 _15380_/X sky130_fd_sc_hd__mux4_2
X_12592_ _12592_/A _12592_/B _12592_/C _12752_/B vssd1 vssd1 vccd1 vccd1 _12775_/A
+ sky130_fd_sc_hd__and4_1
X_14331_ _14409_/A _14331_/B vssd1 vssd1 vccd1 vccd1 _14333_/B sky130_fd_sc_hd__or2_1
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11543_ _11543_/A _11543_/B _11542_/X vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__or3b_2
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ _14262_/A _14340_/A _14262_/C vssd1 vssd1 vccd1 vccd1 _14265_/B sky130_fd_sc_hd__or3_4
XFILLER_167_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17050_ _17088_/B _17050_/B vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__or2_1
XFILLER_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ _11430_/A _11430_/C _11430_/B vssd1 vssd1 vccd1 vccd1 _11475_/C sky130_fd_sc_hd__o21ai_4
XFILLER_167_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13213_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__or3_1
X_16001_ _16001_/A _16001_/B vssd1 vssd1 vccd1 vccd1 _16004_/A sky130_fd_sc_hd__nand2_1
X_10425_ _10427_/B _10427_/C _10427_/A vssd1 vssd1 vccd1 vccd1 _10425_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_183_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14193_ _14270_/A _14193_/B vssd1 vssd1 vccd1 vccd1 _14195_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ _12028_/X _12056_/X _13627_/S vssd1 vssd1 vccd1 vccd1 _13145_/B sky130_fd_sc_hd__mux2_1
X_10356_ _10283_/X _10356_/B vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__nand2b_4
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13075_ _13075_/A _13075_/B _13075_/C vssd1 vssd1 vccd1 vccd1 _13075_/Y sky130_fd_sc_hd__nand3_4
X_10287_ _10187_/X _10285_/Y _10283_/C _10266_/X vssd1 vssd1 vccd1 vccd1 _10287_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_151_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16903_ _16838_/A _16838_/B _16836_/A vssd1 vssd1 vccd1 vccd1 _16905_/B sky130_fd_sc_hd__a21o_2
X_12026_ _14949_/A _14948_/C _12031_/A vssd1 vssd1 vccd1 vccd1 _12026_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_39_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16834_ _16835_/A _16835_/B _16835_/C vssd1 vssd1 vccd1 vccd1 _16836_/A sky130_fd_sc_hd__o21a_1
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16765_ _16765_/A _16765_/B vssd1 vssd1 vccd1 vccd1 _16767_/B sky130_fd_sc_hd__or2_1
X_13977_ _14599_/A _13977_/B _14213_/C _14213_/D vssd1 vssd1 vccd1 vccd1 _13978_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15716_ _14963_/X _15715_/X _15714_/Y _15712_/X _15710_/X vssd1 vssd1 vccd1 vccd1
+ _15716_/X sky130_fd_sc_hd__o2111a_1
X_12928_ _12928_/A _12928_/B _12928_/C vssd1 vssd1 vccd1 vccd1 _12929_/B sky130_fd_sc_hd__or3_1
X_16696_ _16697_/A _16697_/B _16697_/C vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15647_ _15647_/A _16246_/A vssd1 vssd1 vccd1 vccd1 _15648_/B sky130_fd_sc_hd__nand2_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _13837_/A _12857_/X _12858_/Y _13837_/C vssd1 vssd1 vccd1 vccd1 _15457_/C
+ sky130_fd_sc_hd__o22a_2
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15578_ _16056_/A _15578_/B _15774_/B vssd1 vssd1 vccd1 vccd1 _15580_/A sky130_fd_sc_hd__and3_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17317_ input37/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__or3_1
X_14529_ _14583_/B _14529_/B vssd1 vssd1 vccd1 vccd1 _14531_/C sky130_fd_sc_hd__and2_1
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17248_ _17450_/Q _17290_/A2 _17246_/X _17247_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17450_/D sky130_fd_sc_hd__o221a_1
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17179_ input10/X input13/X input12/X input16/X vssd1 vssd1 vccd1 vccd1 _17180_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08952_ _08953_/A _08953_/C vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08883_ _08883_/A _08883_/B _08889_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__or3_2
XFILLER_9_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _09504_/A _09504_/B vssd1 vssd1 vccd1 vccd1 _09657_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _09436_/A _09435_/B _09435_/C vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__nand3_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__nand3_1
XFILLER_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_40 _11791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09297_ _12907_/A _11881_/D _09061_/A _09059_/Y vssd1 vssd1 vccd1 vccd1 _09298_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_51 _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_62 _15996_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 _17562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_95 fanout757/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10210_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__xnor2_2
X_11190_ _11190_/A _11222_/A _11190_/C vssd1 vssd1 vccd1 vccd1 _11222_/B sky130_fd_sc_hd__nor3_4
XFILLER_106_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10141_ _10392_/A _10738_/D vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__and2_4
XFILLER_0_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10072_ _10560_/B _12127_/C _10073_/A vssd1 vssd1 vccd1 vccd1 _10072_/Y sky130_fd_sc_hd__nand3_4
XFILLER_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _13901_/B _13900_/B vssd1 vssd1 vccd1 vccd1 _13902_/A sky130_fd_sc_hd__nand2b_1
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14880_ _17612_/Q _15262_/D _14877_/Y vssd1 vssd1 vccd1 vccd1 _14880_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _12844_/X _12852_/B _17164_/A vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16550_ _16550_/A _16550_/B _16550_/C vssd1 vssd1 vccd1 vccd1 _16551_/B sky130_fd_sc_hd__nand3_1
XFILLER_62_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13762_ _13762_/A _13762_/B vssd1 vssd1 vccd1 vccd1 _13768_/A sky130_fd_sc_hd__nor2_4
XFILLER_44_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _10974_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__xnor2_4
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ _15501_/A _15501_/B _15501_/C vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__nor3_2
XFILLER_16_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12713_ _17399_/A _13564_/C _13450_/D _17403_/A vssd1 vssd1 vccd1 vccd1 _12715_/A
+ sky130_fd_sc_hd__a22oi_2
X_16481_ _16481_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _16481_/X sky130_fd_sc_hd__and2_1
XFILLER_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13693_ _16796_/A _13693_/B _13793_/A vssd1 vssd1 vccd1 vccd1 _13793_/B sky130_fd_sc_hd__nor3_2
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15432_ _15433_/A _15433_/B vssd1 vssd1 vccd1 vccd1 _15514_/B sky130_fd_sc_hd__nand2_1
XFILLER_188_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12644_ _12644_/A _12798_/A vssd1 vssd1 vccd1 vccd1 _12645_/C sky130_fd_sc_hd__and2_2
XFILLER_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _17389_/A _12576_/C _12576_/D _17391_/A vssd1 vssd1 vccd1 vccd1 _12577_/A
+ sky130_fd_sc_hd__a22oi_2
X_15363_ _15363_/A _15363_/B vssd1 vssd1 vccd1 vccd1 _15366_/B sky130_fd_sc_hd__xnor2_1
XFILLER_178_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17102_ _17064_/X _17067_/Y _17099_/A _17100_/X vssd1 vssd1 vccd1 vccd1 _17102_/X
+ sky130_fd_sc_hd__a211o_1
X_14314_ _14315_/A _14315_/B vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__or2_2
XFILLER_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ _11526_/A _11526_/B vssd1 vssd1 vccd1 vccd1 _11526_/Y sky130_fd_sc_hd__nand2_1
XFILLER_102_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15294_ _15295_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _15294_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17033_ _17033_/A _17033_/B _17033_/C _17033_/D vssd1 vssd1 vccd1 vccd1 _17035_/B
+ sky130_fd_sc_hd__and4_1
X_14245_ _14245_/A _14245_/B _14245_/C vssd1 vssd1 vccd1 vccd1 _14247_/A sky130_fd_sc_hd__or3_1
X_11457_ _11456_/B _11456_/C _11456_/A vssd1 vssd1 vccd1 vccd1 _11458_/C sky130_fd_sc_hd__o21bai_4
XFILLER_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ _10315_/A _10315_/B _10315_/C vssd1 vssd1 vccd1 vccd1 _10408_/Y sky130_fd_sc_hd__a21oi_4
X_14176_ _14326_/A _14318_/C _14177_/A vssd1 vssd1 vccd1 vccd1 _14252_/B sky130_fd_sc_hd__nand3_2
XFILLER_139_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11388_ _11630_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11436_/A sky130_fd_sc_hd__nand2_2
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _10215_/B _10228_/Y _10336_/A _10336_/Y vssd1 vssd1 vccd1 vccd1 _10340_/B
+ sky130_fd_sc_hd__a211o_1
X_13127_ _12980_/X _12984_/A _13258_/A _13125_/X vssd1 vssd1 vccd1 vccd1 _13127_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13058_ _13199_/A _13058_/B vssd1 vssd1 vccd1 vccd1 _13060_/B sky130_fd_sc_hd__nor2_4
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12009_ _12009_/A vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__clkinv_2
XFILLER_61_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16817_ _16818_/A _16818_/B vssd1 vssd1 vccd1 vccd1 _16819_/A sky130_fd_sc_hd__or2_1
XFILLER_93_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16748_ _16814_/A _16938_/D _16748_/C vssd1 vssd1 vccd1 vccd1 _16749_/B sky130_fd_sc_hd__or3_2
XFILLER_47_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16679_ _16807_/A _16760_/B _16603_/X _16604_/X vssd1 vssd1 vccd1 vccd1 _16688_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09220_ _09220_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _09221_/C sky130_fd_sc_hd__nor2_1
XFILLER_50_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09151_ _09153_/A _09153_/B _09153_/C vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__o21ai_2
XFILLER_148_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09082_ _11932_/A _11813_/B _08957_/C _08957_/D vssd1 vssd1 vccd1 vccd1 _09084_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput60 i_wb_data[31] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _10241_/B _10491_/B _10490_/C _10115_/A vssd1 vssd1 vccd1 vccd1 _09986_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ _11930_/B _12102_/D _12734_/C _09470_/A vssd1 vssd1 vccd1 vccd1 _08936_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__nor2_1
XFILLER_111_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08797_ _08798_/A _08821_/A _08798_/C vssd1 vssd1 vccd1 vccd1 _11911_/B sky130_fd_sc_hd__o21ai_2
XFILLER_38_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09418_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09434_/C sky130_fd_sc_hd__nand2_1
XFILLER_164_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__xor2_4
XFILLER_185_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09349_ _10542_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _14982_/B sky130_fd_sc_hd__and2_2
XFILLER_166_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12360_ _12360_/A _12360_/B vssd1 vssd1 vccd1 vccd1 _12361_/C sky130_fd_sc_hd__nand2_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ _11311_/A _11311_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__or3_4
XFILLER_180_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _12122_/A _12122_/Y _12289_/Y _12290_/X vssd1 vssd1 vccd1 vccd1 _12312_/A
+ sky130_fd_sc_hd__a211o_2
X_14030_ _14030_/A _14030_/B _14030_/C vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__nand3_1
X_11242_ _11242_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__nor2_4
XFILLER_141_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ _11202_/A _11171_/Y _10988_/Y _10999_/X vssd1 vssd1 vccd1 vccd1 _11186_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ _10125_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__nand2b_2
XFILLER_122_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15981_ _15981_/A _15981_/B vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__nor2_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10055_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14932_ _16207_/B _14931_/X _11841_/A vssd1 vssd1 vccd1 vccd1 _14932_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14863_ _14863_/A _14863_/B _16652_/B vssd1 vssd1 vccd1 vccd1 _14864_/B sky130_fd_sc_hd__and3_1
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16602_ _16517_/A _16517_/B _16515_/B vssd1 vssd1 vccd1 vccd1 _16611_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13814_ _13814_/A _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13815_/B sky130_fd_sc_hd__or3_1
XFILLER_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17582_ fanout934/X _17582_/D vssd1 vssd1 vccd1 vccd1 _17582_/Q sky130_fd_sc_hd__dfxtp_1
X_14794_ _14794_/A _14794_/B vssd1 vssd1 vccd1 vccd1 _14796_/C sky130_fd_sc_hd__or2_2
XFILLER_169_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16533_ _16533_/A _16533_/B _16533_/C vssd1 vssd1 vccd1 vccd1 _16622_/A sky130_fd_sc_hd__and3_2
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ _13852_/A _13745_/B _13948_/C _13745_/D vssd1 vssd1 vccd1 vccd1 _13858_/A
+ sky130_fd_sc_hd__and4_1
X_10957_ _11010_/A _10957_/B _11005_/A _10957_/D vssd1 vssd1 vccd1 vccd1 _11010_/B
+ sky130_fd_sc_hd__and4b_2
XFILLER_73_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16464_ _16362_/A _16362_/B _16365_/A vssd1 vssd1 vccd1 vccd1 _16466_/B sky130_fd_sc_hd__a21oi_4
X_13676_ _13676_/A _13676_/B vssd1 vssd1 vccd1 vccd1 _13678_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ _10891_/B _10888_/B vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__nor2_2
XFILLER_188_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15415_ _15415_/A _16041_/A vssd1 vssd1 vccd1 vccd1 _15417_/B sky130_fd_sc_hd__or2_4
X_12627_ _12820_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__nand2_2
X_16395_ _16394_/A _16394_/B _16396_/A vssd1 vssd1 vccd1 vccd1 _16395_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_185_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15346_ _15346_/A _15346_/B vssd1 vssd1 vccd1 vccd1 _15428_/B sky130_fd_sc_hd__xnor2_4
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _14774_/A _16571_/A vssd1 vssd1 vccd1 vccd1 _12869_/C sky130_fd_sc_hd__and2_4
XFILLER_89_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11509_ _11506_/X _11509_/B _11553_/B _14792_/B vssd1 vssd1 vccd1 vccd1 _11555_/A
+ sky130_fd_sc_hd__and4b_1
X_15277_ _15277_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__xor2_4
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12489_ _12490_/A _12642_/A _12490_/C vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__o21a_1
X_17016_ _17063_/A _17016_/B _17016_/C vssd1 vssd1 vccd1 vccd1 _17035_/A sky130_fd_sc_hd__or3_1
X_14228_ _14229_/A _14229_/B _14229_/C vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__o21a_1
XFILLER_176_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14159_ _14159_/A _14159_/B vssd1 vssd1 vccd1 vccd1 _14161_/A sky130_fd_sc_hd__nor2_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout609 _08969_/B vssd1 vssd1 vccd1 vccd1 _12442_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_112_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _10647_/C vssd1 vssd1 vccd1 vccd1 _08720_/Y sky130_fd_sc_hd__inv_2
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _09942_/A _09637_/B _09937_/B _09803_/B vssd1 vssd1 vccd1 vccd1 _09206_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09134_ _09172_/A _10067_/B _10446_/B _09360_/A vssd1 vssd1 vccd1 vccd1 _09135_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09065_ _09065_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__nor2_1
XFILLER_191_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09967_ _09969_/A _09969_/B _09969_/C vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__o21a_2
XFILLER_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08918_ _08918_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09902_/A _09898_/C vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__or3_1
XTAP_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08849_ _17375_/A _12734_/C _08846_/Y _08996_/A vssd1 vssd1 vccd1 vccd1 _08850_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_73_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _11860_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__nor2_2
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10812_/A _10810_/Y _10962_/A _11005_/B vssd1 vssd1 vccd1 vccd1 _10823_/A
+ sky130_fd_sc_hd__and4bb_2
X_11791_ _15069_/A _11791_/B _11791_/C _12578_/A vssd1 vssd1 vccd1 vccd1 _15262_/D
+ sky130_fd_sc_hd__or4_2
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13530_ _13745_/B _13948_/D _13844_/D _13641_/A vssd1 vssd1 vccd1 vccd1 _13532_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_41_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10742_ _10742_/A _10747_/A _10742_/C vssd1 vssd1 vccd1 vccd1 _10750_/B sky130_fd_sc_hd__or3_2
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13461_ _13462_/A _13462_/B _13462_/C vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__a21oi_2
X_10673_ _10673_/A _10673_/B vssd1 vssd1 vccd1 vccd1 _10675_/B sky130_fd_sc_hd__xnor2_4
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15200_ _14887_/B _15198_/X _14924_/A vssd1 vssd1 vccd1 vccd1 _16262_/A sky130_fd_sc_hd__a21bo_4
XFILLER_138_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__xor2_4
X_16180_ _16279_/C _16180_/B vssd1 vssd1 vccd1 vccd1 _16181_/B sky130_fd_sc_hd__nor2_1
XFILLER_167_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _12387_/X _12391_/X _17369_/A vssd1 vssd1 vccd1 vccd1 _13393_/B sky130_fd_sc_hd__mux2_1
XFILLER_166_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15131_ _15131_/A _15131_/B vssd1 vssd1 vccd1 vccd1 _15131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12343_ _12343_/A _12343_/B _12343_/C vssd1 vssd1 vccd1 vccd1 _12344_/B sky130_fd_sc_hd__nor3_1
XFILLER_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12274_ _17383_/A _12578_/B _12576_/C _12275_/A vssd1 vssd1 vccd1 vccd1 _12276_/A
+ sky130_fd_sc_hd__a22oi_2
X_15062_ _17302_/A1 _11629_/C _14848_/B _14848_/A _15062_/S0 _12398_/S vssd1 vssd1
+ vccd1 vccd1 _15063_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14013_ _14013_/A _14013_/B _14013_/C vssd1 vssd1 vccd1 vccd1 _14015_/C sky130_fd_sc_hd__and3_1
X_11225_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__xnor2_4
XFILLER_49_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ _11155_/A _11234_/A _11232_/A vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__o21ai_4
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10107_ _09981_/C _17469_/D _09982_/A _09980_/Y vssd1 vssd1 vccd1 vccd1 _10113_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15964_ _15964_/A _15964_/B vssd1 vssd1 vccd1 vccd1 _15966_/C sky130_fd_sc_hd__xnor2_2
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11087_ _11087_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10038_ _10039_/A _10037_/Y _10970_/A _10755_/D vssd1 vssd1 vccd1 vccd1 _10151_/A
+ sky130_fd_sc_hd__and4bb_2
X_14915_ _14958_/A _14915_/B vssd1 vssd1 vccd1 vccd1 _14915_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15895_ _16933_/A _15895_/B _15895_/C vssd1 vssd1 vccd1 vccd1 _15897_/B sky130_fd_sc_hd__and3_1
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14846_ _15274_/A _14846_/B vssd1 vssd1 vccd1 vccd1 _15110_/B sky130_fd_sc_hd__nor2_2
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17565_ fanout945/X _17565_/D vssd1 vssd1 vccd1 vccd1 _17565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14777_ _14777_/A _16298_/A vssd1 vssd1 vccd1 vccd1 _16302_/B sky130_fd_sc_hd__or2_2
X_11989_ _11990_/A _11990_/B _11990_/C vssd1 vssd1 vccd1 vccd1 _12155_/A sky130_fd_sc_hd__a21oi_4
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16516_ _16938_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16517_/B sky130_fd_sc_hd__nand2_1
XFILLER_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ _13619_/A _13616_/Y _13617_/X vssd1 vssd1 vccd1 vccd1 _13728_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ fanout930/X _17496_/D vssd1 vssd1 vccd1 vccd1 _17496_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16447_ _16533_/A _16355_/B _16352_/C vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__a21oi_4
X_13659_ _13659_/A _13659_/B vssd1 vssd1 vccd1 vccd1 _13662_/C sky130_fd_sc_hd__xnor2_2
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16378_ _16378_/A _16378_/B vssd1 vssd1 vccd1 vccd1 _16381_/A sky130_fd_sc_hd__xnor2_4
XFILLER_191_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ _15553_/A _15553_/B _15752_/B vssd1 vssd1 vccd1 vccd1 _15331_/B sky130_fd_sc_hd__or3_4
XFILLER_144_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout406 _09981_/C vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _09819_/A _09819_/B _09819_/C vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__o21a_1
XFILLER_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout417 _14776_/A vssd1 vssd1 vccd1 vccd1 _17399_/A sky130_fd_sc_hd__buf_8
Xfanout428 _14777_/A vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__buf_4
Xfanout439 _12079_/A vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__buf_12
XFILLER_101_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09752_ _15537_/A _09928_/D _09746_/A _09612_/Y vssd1 vssd1 vccd1 vccd1 _09754_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09683_ _09668_/A _09668_/C _09668_/B vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09117_ _08930_/X _09018_/Y _09071_/A _09259_/A vssd1 vssd1 vccd1 vccd1 _09119_/D
+ sky130_fd_sc_hd__a211o_2
XFILLER_109_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09048_ _09048_/A _09048_/B _09048_/C vssd1 vssd1 vccd1 vccd1 _09049_/C sky130_fd_sc_hd__nand3_2
XFILLER_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11010_ _11010_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout940 fanout944/X vssd1 vssd1 vccd1 vccd1 fanout940/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12961_ _12771_/A _12773_/B _12771_/B vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__o21ba_2
XTAP_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _14701_/A _14701_/B vssd1 vssd1 vccd1 vccd1 _14700_/Y sky130_fd_sc_hd__nand2_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _08863_/X _08867_/A _12148_/A _11911_/Y vssd1 vssd1 vccd1 vccd1 _12148_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _15772_/B _15679_/C _15679_/A vssd1 vssd1 vccd1 vccd1 _15682_/B sky130_fd_sc_hd__a21oi_4
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _17387_/A _13169_/D _12889_/Y _13043_/A vssd1 vssd1 vccd1 vccd1 _12893_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14631_ _14631_/A _14631_/B vssd1 vssd1 vccd1 vccd1 _14633_/B sky130_fd_sc_hd__or2_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11843_ _11840_/Y _11842_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__mux2_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _13903_/B _17354_/A2 _17349_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17504_/D
+ sky130_fd_sc_hd__o211a_1
X_14562_ _14562_/A _14562_/B _14562_/C vssd1 vssd1 vccd1 vccd1 _14564_/C sky130_fd_sc_hd__nand3_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _10347_/X _11775_/B _11775_/A vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16301_/A _16301_/B vssd1 vssd1 vccd1 vccd1 _16301_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13513_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13513_/Y sky130_fd_sc_hd__nand2_1
X_17281_ _17461_/Q _17290_/A2 _17279_/X _17280_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17461_/D sky130_fd_sc_hd__o221a_1
XFILLER_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10725_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _10725_/X sky130_fd_sc_hd__and2_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14493_ _16965_/C _14708_/D _14493_/C vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__and3_1
X_16232_ _16232_/A _16232_/B vssd1 vssd1 vccd1 vccd1 _16239_/A sky130_fd_sc_hd__xor2_2
X_13444_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13444_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10656_ _11629_/B _11841_/B vssd1 vssd1 vccd1 vccd1 _10657_/C sky130_fd_sc_hd__and2_4
XFILLER_167_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16163_ _16044_/A _16044_/B _16045_/X vssd1 vssd1 vccd1 vccd1 _16177_/A sky130_fd_sc_hd__a21oi_2
X_10587_ _10555_/A _10555_/C _10555_/B vssd1 vssd1 vccd1 vccd1 _10587_/Y sky130_fd_sc_hd__o21ai_4
X_13375_ _13249_/A _13249_/Y _13494_/B _13374_/X vssd1 vssd1 vccd1 vccd1 _13500_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_166_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15114_ _14790_/A _16735_/A _12230_/B _15113_/X vssd1 vssd1 vccd1 vccd1 _15114_/X
+ sky130_fd_sc_hd__o31a_1
X_12326_ _12325_/A _12325_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__o21ai_1
X_16094_ _16095_/B _16095_/A vssd1 vssd1 vccd1 vccd1 _16200_/B sky130_fd_sc_hd__nand2b_2
XFILLER_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _15041_/X _15042_/X _15043_/X _15309_/B vssd1 vssd1 vccd1 vccd1 _15045_/X
+ sky130_fd_sc_hd__a31o_1
X_12257_ _12257_/A _12257_/B vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__nor2_2
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11208_ _10761_/A _11206_/Y _11178_/Y _11175_/Y vssd1 vssd1 vccd1 vccd1 _11208_/Y
+ sky130_fd_sc_hd__o211ai_4
X_12188_ _12188_/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12189_/B sky130_fd_sc_hd__or2_1
XFILLER_68_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _11139_/A _11139_/B _11139_/C vssd1 vssd1 vccd1 vccd1 _11255_/A sky130_fd_sc_hd__and3_4
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16996_ _16995_/B _16996_/B vssd1 vssd1 vccd1 vccd1 _17052_/A sky130_fd_sc_hd__and2b_1
XFILLER_96_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15947_ _16880_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16827_/C sky130_fd_sc_hd__nand2_4
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15878_ _15992_/A _15878_/B vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__nand2b_1
XFILLER_58_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14829_ _17134_/A _14829_/B vssd1 vssd1 vccd1 vccd1 _14829_/X sky130_fd_sc_hd__or2_4
XFILLER_24_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17548_ fanout946/X _17548_/D vssd1 vssd1 vccd1 vccd1 _17548_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_189_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17479_ fanout926/X _17479_/D vssd1 vssd1 vccd1 vccd1 _17479_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_165_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout203 _11853_/Y vssd1 vssd1 vccd1 vccd1 _12401_/A sky130_fd_sc_hd__buf_6
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout214 _17196_/X vssd1 vssd1 vccd1 vccd1 _17362_/C sky130_fd_sc_hd__buf_6
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _15454_/A vssd1 vssd1 vccd1 vccd1 _16917_/A sky130_fd_sc_hd__buf_6
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout236 _14926_/B vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__buf_4
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09804_ _09805_/B _09939_/A _09805_/A vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__o21ai_4
XFILLER_59_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout247 _16304_/A vssd1 vssd1 vccd1 vccd1 _17169_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout258 _17295_/X vssd1 vssd1 vccd1 vccd1 _17429_/C sky130_fd_sc_hd__buf_4
Xfanout269 _16644_/B vssd1 vssd1 vccd1 vccd1 _17134_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09735_ _09735_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__nor2_1
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09666_ _09666_/A _09666_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__and2_2
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09597_/A _09597_/B _09686_/B vssd1 vssd1 vccd1 vccd1 _09624_/C sky130_fd_sc_hd__and3_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _10511_/B _10511_/A vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__and2b_2
X_11490_ _11456_/A _11456_/C _11456_/B vssd1 vssd1 vccd1 vccd1 _11490_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10441_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__xnor2_4
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13160_ _13161_/A _13161_/B vssd1 vssd1 vccd1 vccd1 _13295_/B sky130_fd_sc_hd__nand2_2
X_10372_ _10372_/A _10372_/B vssd1 vssd1 vccd1 vccd1 _10374_/C sky130_fd_sc_hd__xnor2_2
XFILLER_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _11901_/A _11903_/B _11901_/B vssd1 vssd1 vccd1 vccd1 _12113_/B sky130_fd_sc_hd__o21ba_2
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13091_ _13092_/A _13092_/B _13092_/C vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__a21oi_1
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _12700_/D _12042_/B vssd1 vssd1 vccd1 vccd1 _12042_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16850_ _16850_/A _16850_/B vssd1 vssd1 vccd1 vccd1 _16851_/B sky130_fd_sc_hd__or2_1
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout770 _13196_/B vssd1 vssd1 vccd1 vccd1 _12637_/D sky130_fd_sc_hd__buf_12
X_15801_ _15801_/A _15801_/B vssd1 vssd1 vccd1 vccd1 _15802_/B sky130_fd_sc_hd__and2_1
XFILLER_59_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout781 _09030_/D vssd1 vssd1 vccd1 vccd1 _12659_/B sky130_fd_sc_hd__buf_12
X_16781_ _16781_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16782_/B sky130_fd_sc_hd__and2_1
XFILLER_19_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout792 _17489_/Q vssd1 vssd1 vccd1 vccd1 _09414_/C sky130_fd_sc_hd__buf_6
X_13993_ _16913_/C _14865_/B vssd1 vssd1 vccd1 vccd1 _16918_/A sky130_fd_sc_hd__nand2_4
XFILLER_46_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15732_ _15732_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15741_/A sky130_fd_sc_hd__xnor2_4
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12944_ _12945_/A _13085_/A _12945_/C vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__o21a_1
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _15663_/A _15663_/B vssd1 vssd1 vccd1 vccd1 _15673_/A sky130_fd_sc_hd__xnor2_4
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12875_/A _12875_/B vssd1 vssd1 vccd1 vccd1 _12884_/A sky130_fd_sc_hd__xor2_4
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ input46/X _17422_/A2 _17401_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17529_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14614_ _14615_/B _14614_/B vssd1 vssd1 vccd1 vccd1 _14658_/A sky130_fd_sc_hd__and2b_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _12700_/D _11826_/B vssd1 vssd1 vccd1 vccd1 _11826_/Y sky130_fd_sc_hd__nand2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15594_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15595_/B sky130_fd_sc_hd__or2_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ input45/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17333_/X sky130_fd_sc_hd__or3_1
X_14545_ _14593_/A _14593_/B _14545_/C _14545_/D vssd1 vssd1 vccd1 vccd1 _14601_/A
+ sky130_fd_sc_hd__and4_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11757_ _11732_/Y _11733_/X _11737_/Y _11753_/A vssd1 vssd1 vccd1 vccd1 _11758_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17264_ _17597_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17264_/X sky130_fd_sc_hd__a21o_1
XFILLER_140_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__xnor2_4
XFILLER_174_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14476_ _14533_/B _14533_/C vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11688_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _15302_/B sky130_fd_sc_hd__xor2_1
X_16215_ _08760_/Y _14778_/X _14813_/X _16304_/A _16214_/Y vssd1 vssd1 vccd1 vccd1
+ _16215_/X sky130_fd_sc_hd__a311o_1
X_13427_ _13304_/A _13304_/B _13305_/Y vssd1 vssd1 vccd1 vccd1 _13427_/X sky130_fd_sc_hd__a21bo_1
X_17195_ _17195_/A _17195_/B _17195_/C vssd1 vssd1 vccd1 vccd1 _17196_/C sky130_fd_sc_hd__or3_1
X_10639_ _11258_/B _10933_/D _10970_/B _11314_/A vssd1 vssd1 vccd1 vccd1 _10639_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_155_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _16146_/A _16146_/B vssd1 vssd1 vccd1 vccd1 _16158_/A sky130_fd_sc_hd__xnor2_4
X_13358_ _13228_/A _13230_/B _13228_/B vssd1 vssd1 vccd1 vccd1 _13360_/B sky130_fd_sc_hd__o21ba_1
XFILLER_182_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ _12309_/A _12309_/B _12309_/C vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__and3_1
X_16077_ _16077_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16078_/B sky130_fd_sc_hd__nor2_1
X_13289_ _13643_/A _13844_/D _13286_/Y _13417_/A vssd1 vssd1 vccd1 vccd1 _13290_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_142_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15028_ _15028_/A _15687_/A vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__or2_2
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16979_ _17169_/A1 _16971_/Y _16972_/Y _15794_/A _16978_/X vssd1 vssd1 vccd1 vccd1
+ _16979_/X sky130_fd_sc_hd__o221a_1
Xinput3 i_wb_addr[0] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09520_ _10067_/A _09791_/B _09520_/C vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__and3_1
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09451_ _09451_/A _09451_/B vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ _10067_/A _12770_/D _09382_/C vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__and3_2
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ _09718_/A _09718_/B _09718_/C vssd1 vssd1 vccd1 vccd1 _09719_/C sky130_fd_sc_hd__nand3_1
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__nand3_2
XFILLER_142_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _09969_/B _09649_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__nor2_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _12662_/C sky130_fd_sc_hd__xnor2_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11617_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _11612_/C sky130_fd_sc_hd__and2_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _12592_/A _12592_/C vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__nand2_1
XFILLER_169_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14330_ _14330_/A _14330_/B _14330_/C vssd1 vssd1 vccd1 vccd1 _14331_/B sky130_fd_sc_hd__and3_1
XFILLER_184_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _11542_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__or2_1
XFILLER_156_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14261_ _14340_/A _14262_/C _14262_/A vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__o21ai_1
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11473_ _11469_/X _11471_/X _11472_/A vssd1 vssd1 vccd1 vccd1 _11475_/B sky130_fd_sc_hd__a21o_2
XFILLER_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16000_ _16014_/A _17153_/B _16317_/A vssd1 vssd1 vccd1 vccd1 _16001_/B sky130_fd_sc_hd__or3b_1
XFILLER_171_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13212_ _13212_/A _13339_/B vssd1 vssd1 vccd1 vccd1 _13213_/C sky130_fd_sc_hd__nor2_1
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10424_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10427_/C sky130_fd_sc_hd__nand2_2
XFILLER_171_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14192_ _14192_/A _14192_/B _14192_/C vssd1 vssd1 vccd1 vccd1 _14193_/B sky130_fd_sc_hd__nand3_1
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13143_ _15457_/B _13142_/X _17165_/A1 vssd1 vssd1 vccd1 vccd1 _13143_/Y sky130_fd_sc_hd__o21ai_1
X_10355_ _10283_/B _10283_/C _10283_/D _10283_/A vssd1 vssd1 vccd1 vccd1 _10356_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10266_/X _10283_/C _10285_/Y _10187_/X vssd1 vssd1 vccd1 vccd1 _10330_/A
+ sky130_fd_sc_hd__a211o_4
X_13074_ _13075_/A _13075_/B _13075_/C vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__a21o_2
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16902_ _16902_/A _16902_/B vssd1 vssd1 vccd1 vccd1 _16905_/A sky130_fd_sc_hd__nor2_4
X_12025_ _17363_/A _12025_/B vssd1 vssd1 vccd1 vccd1 _14948_/C sky130_fd_sc_hd__and2_1
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16833_ _16833_/A _16897_/B vssd1 vssd1 vccd1 vccd1 _16835_/C sky130_fd_sc_hd__nor2_1
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16764_ _16763_/B _16764_/B vssd1 vssd1 vccd1 vccd1 _16765_/B sky130_fd_sc_hd__and2b_1
XFILLER_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13976_ _13977_/B _14213_/C _14213_/D _14599_/A vssd1 vssd1 vccd1 vccd1 _13978_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15715_ _16011_/A _15715_/B vssd1 vssd1 vccd1 vccd1 _15715_/X sky130_fd_sc_hd__or2_4
X_12927_ _12928_/A _12928_/B _12928_/C vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__o21ai_2
X_16695_ _16695_/A _16695_/B _16695_/C vssd1 vssd1 vccd1 vccd1 _16697_/C sky130_fd_sc_hd__and3_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15646_ _15734_/A _15645_/B _16150_/B _15644_/X vssd1 vssd1 vccd1 vccd1 _15648_/A
+ sky130_fd_sc_hd__o31a_4
X_12858_ _15537_/A _15384_/S vssd1 vssd1 vccd1 vccd1 _12858_/Y sky130_fd_sc_hd__nand2_8
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11809_ _09652_/C _14982_/C _14912_/B vssd1 vssd1 vccd1 vccd1 _11809_/Y sky130_fd_sc_hd__o21ai_2
X_15577_ _16056_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15577_/Y sky130_fd_sc_hd__nand2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12790_/A _12947_/A _12790_/C vssd1 vssd1 vccd1 vccd1 _12791_/A sky130_fd_sc_hd__o21a_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _12923_/D _17328_/A2 _17315_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17487_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_193_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14528_ _14528_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _14529_/B sky130_fd_sc_hd__nand2_1
XFILLER_175_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17247_ _17559_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17247_/X sky130_fd_sc_hd__and2_1
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14459_ _14518_/A _14459_/B _14459_/C vssd1 vssd1 vccd1 vccd1 _14518_/B sky130_fd_sc_hd__nand3_4
XFILLER_190_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17178_ input6/X input9/X input8/X input11/X vssd1 vssd1 vccd1 vccd1 _17180_/C sky130_fd_sc_hd__or4_1
XFILLER_190_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16129_ _16226_/B _16129_/B vssd1 vssd1 vccd1 vccd1 _16130_/B sky130_fd_sc_hd__nand2_2
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08951_ _11932_/A _12595_/C _08936_/C _08936_/D vssd1 vssd1 vccd1 vccd1 _08953_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ _08882_/A _09027_/A vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__nor2_4
XFILLER_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1026 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09503_ _09502_/A _09944_/D _09497_/A _09361_/Y vssd1 vssd1 vccd1 vccd1 _09504_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_112_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09434_ _09434_/A _09434_/B _09434_/C vssd1 vssd1 vccd1 vccd1 _09435_/C sky130_fd_sc_hd__nand3_2
XFILLER_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _09497_/A _09504_/A _09497_/C vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__o21a_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 _17439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _09296_/A _09296_/B _09296_/C vssd1 vssd1 vccd1 vccd1 _09296_/Y sky130_fd_sc_hd__nand3_2
XANTENNA_41 _11902_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_52 _12659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 _17560_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_74 _17476_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_85 _10640_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_96 _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10071_ _10560_/B _12127_/C vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__nand2_1
XFILLER_153_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _13936_/B _13830_/B vssd1 vssd1 vccd1 vccd1 _13830_/X sky130_fd_sc_hd__or2_1
XFILLER_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13762_/B sky130_fd_sc_hd__and2_1
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10973_ _10973_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__nor2_2
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15500_ _15501_/A _15501_/B _15501_/C vssd1 vssd1 vccd1 vccd1 _15594_/A sky130_fd_sc_hd__o21a_2
XFILLER_44_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12712_ _12698_/Y _12699_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _17581_/D sky130_fd_sc_hd__o21ai_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _16480_/A _17153_/B _14775_/A vssd1 vssd1 vccd1 vccd1 _16481_/B sky130_fd_sc_hd__or3b_1
XFILLER_188_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13692_ _13693_/B _13793_/A _16796_/A vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__o21a_1
XFILLER_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ _15431_/A _15431_/B vssd1 vssd1 vccd1 vccd1 _15433_/B sky130_fd_sc_hd__xnor2_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12643_ _12642_/A _12642_/B _12642_/C vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__o21ai_4
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15362_ _15362_/A _15362_/B vssd1 vssd1 vccd1 vccd1 _15363_/B sky130_fd_sc_hd__xnor2_2
X_12574_ _12415_/A _12417_/B _12415_/B vssd1 vssd1 vccd1 vccd1 _12581_/A sky130_fd_sc_hd__o21ba_1
X_17101_ _17099_/A _17100_/X _17064_/X _17067_/Y vssd1 vssd1 vccd1 vccd1 _17103_/B
+ sky130_fd_sc_hd__o211a_1
X_14313_ _14381_/A _14313_/B vssd1 vssd1 vccd1 vccd1 _14315_/B sky130_fd_sc_hd__or2_1
XFILLER_178_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ _11526_/A _11525_/B _11525_/C vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__nand3_4
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15293_ _15159_/A _15159_/B _15221_/B _15226_/A _15226_/B vssd1 vssd1 vccd1 vccd1
+ _15295_/B sky130_fd_sc_hd__a32o_4
XFILLER_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17032_ _16653_/A _14636_/B _16582_/A _15715_/X vssd1 vssd1 vccd1 vccd1 _17033_/D
+ sky130_fd_sc_hd__o22a_1
X_14244_ _14244_/A _14244_/B vssd1 vssd1 vccd1 vccd1 _14245_/C sky130_fd_sc_hd__xnor2_2
XFILLER_137_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11456_ _11456_/A _11456_/B _11456_/C vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__or3_4
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10407_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10407_/Y sky130_fd_sc_hd__nor2_4
X_14175_ _14326_/A _14175_/B vssd1 vssd1 vccd1 vccd1 _14177_/B sky130_fd_sc_hd__nand2_2
XFILLER_178_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11387_ _11480_/A _11480_/C _11387_/C vssd1 vssd1 vccd1 vccd1 _11393_/B sky130_fd_sc_hd__and3_1
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13126_ _12980_/X _12984_/A _13258_/A _13125_/X vssd1 vssd1 vccd1 vccd1 _13258_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10338_ _10451_/A _10334_/B _10332_/X vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__a21o_2
XFILLER_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13057_ _13057_/A _13057_/B _13057_/C vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__nor3_2
XFILLER_140_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10269_ _15262_/B _15624_/A vssd1 vssd1 vccd1 vccd1 _10269_/X sky130_fd_sc_hd__and2_1
X_12008_ _12800_/A _11961_/B _09230_/A _09228_/A vssd1 vssd1 vccd1 vccd1 _12009_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16816_ _16816_/A _16888_/A _16816_/C vssd1 vssd1 vccd1 vccd1 _16818_/B sky130_fd_sc_hd__and3_1
XFILLER_66_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13959_ _14044_/B _13959_/B vssd1 vssd1 vccd1 vccd1 _13961_/C sky130_fd_sc_hd__nor2_1
X_16747_ _16747_/A _16813_/B vssd1 vssd1 vccd1 vccd1 _16883_/C sky130_fd_sc_hd__nor2_4
XFILLER_4_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1032 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16678_ _16770_/A _16678_/B vssd1 vssd1 vccd1 vccd1 _16690_/A sky130_fd_sc_hd__or2_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15629_ _15037_/X _15039_/X _15057_/X _15059_/Y _15130_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15629_/X sky130_fd_sc_hd__mux4_1
XFILLER_148_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09153_/C sky130_fd_sc_hd__xnor2_2
XFILLER_188_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09081_ _09081_/A _09306_/A vssd1 vssd1 vccd1 vccd1 _09088_/A sky130_fd_sc_hd__nor2_1
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 i_wb_data[22] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput61 i_wb_data[3] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09983_ _09983_/A _09983_/B _09989_/B vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__or3_4
X_08934_ _08937_/A vssd1 vssd1 vccd1 vccd1 _08936_/C sky130_fd_sc_hd__inv_2
XFILLER_130_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08865_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__and2_2
XFILLER_184_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08796_ _08796_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _08798_/C sky130_fd_sc_hd__xor2_2
XFILLER_72_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09417_ _09417_/A _09417_/B vssd1 vssd1 vccd1 vccd1 _09546_/B sky130_fd_sc_hd__xnor2_4
XFILLER_38_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09348_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _09355_/A sky130_fd_sc_hd__nor2_2
XFILLER_139_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__xnor2_4
X_11310_ _11285_/A _11285_/B _11285_/C vssd1 vssd1 vccd1 vccd1 _11311_/C sky130_fd_sc_hd__a21oi_2
XFILLER_193_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12290_ _12267_/Y _12268_/X _12476_/B _12290_/D vssd1 vssd1 vccd1 vccd1 _12290_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_107_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11241_ _10962_/A _11097_/D _11098_/A _11096_/Y vssd1 vssd1 vccd1 vccd1 _11242_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _10988_/Y _10999_/X _11202_/A _11171_/Y vssd1 vssd1 vccd1 vccd1 _11202_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10125_/B sky130_fd_sc_hd__xnor2_4
XFILLER_121_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15980_ _15980_/A _15980_/B _15980_/C vssd1 vssd1 vccd1 vccd1 _15981_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__nor2_4
XFILLER_94_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14931_ _17476_/D _17477_/D _14836_/B vssd1 vssd1 vccd1 vccd1 _14931_/X sky130_fd_sc_hd__or3b_4
XFILLER_94_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14862_ _16651_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16652_/B sky130_fd_sc_hd__and2_2
XFILLER_48_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16601_ _16601_/A _16601_/B vssd1 vssd1 vccd1 vccd1 _16614_/A sky130_fd_sc_hd__nand2_1
X_13813_ _13814_/A _13814_/B _13814_/C vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__o21ai_2
XFILLER_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17581_ fanout925/X _17581_/D vssd1 vssd1 vccd1 vccd1 _17581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14793_ _14794_/A _14794_/B vssd1 vssd1 vccd1 vccd1 _14793_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16532_ _16533_/C _16695_/C vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__and2b_1
X_13744_ _13852_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10956_ _11006_/B _11097_/D _11027_/C _11006_/A vssd1 vssd1 vccd1 vccd1 _10957_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16463_ _16557_/A _16463_/B vssd1 vssd1 vccd1 vccd1 _16466_/A sky130_fd_sc_hd__nand2b_4
X_13675_ _14153_/A _14153_/B _14050_/D _13866_/C vssd1 vssd1 vccd1 vccd1 _13676_/B
+ sky130_fd_sc_hd__and4_1
X_10887_ _11629_/B _09712_/B _15206_/A _15130_/S vssd1 vssd1 vccd1 vccd1 _10888_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15414_ _15414_/A _15414_/B vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__xor2_4
X_12626_ _12626_/A _12626_/B _12626_/C vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__nand3_1
XFILLER_188_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16394_ _16394_/A _16394_/B vssd1 vssd1 vccd1 vccd1 _16396_/B sky130_fd_sc_hd__and2_1
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15345_ _15345_/A _15345_/B vssd1 vssd1 vccd1 vccd1 _15346_/B sky130_fd_sc_hd__xnor2_4
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _17399_/A _13564_/D _13966_/D _17403_/A vssd1 vssd1 vccd1 vccd1 _12557_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11508_ _11553_/A _14794_/B _11553_/D _11506_/A vssd1 vssd1 vccd1 vccd1 _11509_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15276_ _15277_/A _15277_/B vssd1 vssd1 vccd1 vccd1 _15276_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12488_ _12488_/A _12637_/C vssd1 vssd1 vccd1 vccd1 _12490_/C sky130_fd_sc_hd__nand2_2
XFILLER_89_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17015_ _17014_/A _17014_/C _17014_/B vssd1 vssd1 vccd1 vccd1 _17016_/C sky130_fd_sc_hd__a21oi_1
X_14227_ _14227_/A _16970_/A vssd1 vssd1 vccd1 vccd1 _14229_/C sky130_fd_sc_hd__xnor2_1
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11439_ _11440_/A _11438_/Y _11520_/C _11480_/C vssd1 vssd1 vccd1 vccd1 _11479_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_171_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14158_ _14158_/A _14158_/B _14158_/C vssd1 vssd1 vccd1 vccd1 _14159_/B sky130_fd_sc_hd__nor3_2
XFILLER_171_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _13109_/A _13109_/B vssd1 vssd1 vccd1 vccd1 _13110_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14326_/A _14089_/B vssd1 vssd1 vccd1 vccd1 _14090_/B sky130_fd_sc_hd__nand2_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09202_ _09202_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09133_ _09502_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09064_ _17375_/A _12258_/B _08950_/A _08948_/Y vssd1 vssd1 vccd1 vccd1 _09065_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09966_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09969_/C sky130_fd_sc_hd__xnor2_1
XFILLER_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08917_ _08918_/B _08918_/A vssd1 vssd1 vccd1 vccd1 _08917_/X sky130_fd_sc_hd__and2b_2
XTAP_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09898_/A _09898_/C vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__nor2_1
XTAP_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _08846_/Y _08996_/A _17375_/A _12734_/C vssd1 vssd1 vccd1 vccd1 _08996_/B
+ sky130_fd_sc_hd__and4bb_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__xor2_4
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10810_ _11240_/A _10957_/D _11097_/D _10963_/A vssd1 vssd1 vccd1 vccd1 _10810_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11791_/C _16136_/A vssd1 vssd1 vccd1 vccd1 _11790_/X sky130_fd_sc_hd__or2_1
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ _10742_/A _10742_/C vssd1 vssd1 vccd1 vccd1 _10747_/B sky130_fd_sc_hd__nor2_2
XFILLER_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _13576_/B _13460_/B vssd1 vssd1 vccd1 vccd1 _13462_/C sky130_fd_sc_hd__nand2_1
XFILLER_186_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10672_ _10672_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10673_/B sky130_fd_sc_hd__and2_4
XFILLER_167_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__and2_1
X_13391_ _12401_/A _13390_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _13391_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15130_ _15131_/B _15129_/X _15130_/S vssd1 vssd1 vccd1 vccd1 _15130_/X sky130_fd_sc_hd__mux2_1
X_12342_ _12343_/A _12343_/B _12343_/C vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__o21a_1
XFILLER_193_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _15131_/A _15061_/B vssd1 vssd1 vccd1 vccd1 _15061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _12273_/A _12273_/B vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14012_ _14013_/A _14013_/B _14013_/C vssd1 vssd1 vccd1 vccd1 _14015_/B sky130_fd_sc_hd__a21oi_1
X_11224_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11224_/X sky130_fd_sc_hd__and2b_1
XFILLER_175_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11155_ _11155_/A _11234_/A vssd1 vssd1 vccd1 vccd1 _11232_/B sky130_fd_sc_hd__nor2_2
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__xnor2_4
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15963_ _15963_/A _15963_/B vssd1 vssd1 vccd1 vccd1 _15964_/B sky130_fd_sc_hd__xor2_4
X_11086_ _11069_/X _11070_/Y _11084_/A _11090_/A vssd1 vssd1 vccd1 vccd1 _11087_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10037_ _10036_/B _10534_/D _10647_/D _10525_/A vssd1 vssd1 vccd1 vccd1 _10037_/Y
+ sky130_fd_sc_hd__a22oi_2
X_14914_ _10013_/B _09712_/B _14942_/A vssd1 vssd1 vccd1 vccd1 _14915_/B sky130_fd_sc_hd__mux2_1
X_15894_ _15890_/X _15891_/X _15892_/Y _15893_/Y _17156_/B vssd1 vssd1 vccd1 vccd1
+ _15894_/X sky130_fd_sc_hd__a311o_1
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14845_ _15008_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _14846_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17564_ fanout945/X _17564_/D vssd1 vssd1 vccd1 vccd1 _17564_/Q sky130_fd_sc_hd__dfxtp_1
X_14776_ _14776_/A _16399_/A vssd1 vssd1 vccd1 vccd1 _16397_/B sky130_fd_sc_hd__or2_1
X_11988_ _11988_/A _11988_/B vssd1 vssd1 vccd1 vccd1 _11990_/C sky130_fd_sc_hd__xnor2_2
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16515_ _16515_/A _16515_/B vssd1 vssd1 vccd1 vccd1 _16517_/A sky130_fd_sc_hd__nand2_1
X_13727_ _13727_/A _13727_/B vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__or2_2
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ _10940_/A _10940_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__nand2_2
XFILLER_31_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17495_ fanout937/X _17495_/D vssd1 vssd1 vccd1 vccd1 _17495_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16446_ _16446_/A _16619_/A _16681_/C _16681_/D vssd1 vssd1 vccd1 vccd1 _16446_/X
+ sky130_fd_sc_hd__or4_2
X_13658_ _13658_/A _13948_/C _13658_/C vssd1 vssd1 vccd1 vccd1 _13659_/B sky130_fd_sc_hd__and3_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12610_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__or2_1
X_16377_ _16378_/B _16378_/A vssd1 vssd1 vccd1 vccd1 _16470_/B sky130_fd_sc_hd__nand2b_1
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ _13589_/A _13589_/B vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__xor2_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15328_ _14899_/X _14968_/X _15752_/B _11675_/B vssd1 vssd1 vccd1 vccd1 _15404_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15259_ _15233_/X _15234_/Y _15258_/X vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout407 _09409_/C vssd1 vssd1 vccd1 vccd1 _09981_/C sky130_fd_sc_hd__buf_2
X_09820_ _09524_/A _09523_/B _09523_/A vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__o21ba_4
Xfanout418 _13948_/B vssd1 vssd1 vccd1 vccd1 _13844_/B sky130_fd_sc_hd__buf_6
XFILLER_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout429 _17527_/Q vssd1 vssd1 vccd1 vccd1 _14777_/A sky130_fd_sc_hd__buf_8
XFILLER_154_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09751_ _09751_/A _09880_/A vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__nor2_2
XFILLER_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09682_ _09674_/B _09670_/X _09631_/Y _09666_/B vssd1 vssd1 vccd1 vccd1 _09819_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _09119_/B _09119_/C vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__nand2_2
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09047_ _09047_/A _09047_/B vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__xnor2_4
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout930 fanout931/X vssd1 vssd1 vccd1 vccd1 fanout930/X sky130_fd_sc_hd__clkbuf_4
Xfanout941 fanout942/X vssd1 vssd1 vccd1 vccd1 fanout941/X sky130_fd_sc_hd__clkbuf_4
X_09949_ _10560_/A _12127_/D _10061_/B vssd1 vssd1 vccd1 vccd1 _09951_/C sky130_fd_sc_hd__and3_1
XFILLER_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ _12960_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _12979_/A sky130_fd_sc_hd__and2_2
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _11911_/A _11911_/B _11911_/C vssd1 vssd1 vccd1 vccd1 _11911_/Y sky130_fd_sc_hd__nand3_2
XFILLER_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12889_/Y _13043_/A _17387_/A _13169_/D vssd1 vssd1 vccd1 vccd1 _13043_/B
+ sky130_fd_sc_hd__and4bb_2
XFILLER_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14585_/A _14582_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14631_/B sky130_fd_sc_hd__a21oi_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _10897_/C _11841_/X _14911_/B vssd1 vssd1 vccd1 vccd1 _11842_/Y sky130_fd_sc_hd__o21ai_4
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14562_/A _14562_/B _14562_/C vssd1 vssd1 vccd1 vccd1 _14612_/A sky130_fd_sc_hd__a21o_1
XFILLER_14_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11773_/A _11773_/B vssd1 vssd1 vccd1 vccd1 _17105_/B sky130_fd_sc_hd__and2_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16300_/A _16300_/B vssd1 vssd1 vccd1 vccd1 _16301_/B sky130_fd_sc_hd__nor2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13010_/B _13511_/X _13510_/X vssd1 vssd1 vccd1 vccd1 _13514_/B sky130_fd_sc_hd__a21oi_2
X_17280_ _17570_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17280_/X sky130_fd_sc_hd__and2_1
X_10724_ _10724_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _11174_/B sky130_fd_sc_hd__nor2_4
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/A _14492_/B vssd1 vssd1 vccd1 vccd1 _14493_/C sky130_fd_sc_hd__xor2_1
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _16232_/A _16232_/B vssd1 vssd1 vccd1 vccd1 _16231_/Y sky130_fd_sc_hd__nand2_1
X_13443_ _13443_/A _13443_/B _13443_/C vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__and3_2
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10655_ _10655_/A _10655_/B vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__nor2_4
XFILLER_186_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16162_ _16068_/A _16068_/B _16069_/Y vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__a21bo_1
XFILLER_127_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13374_ _13494_/A _13373_/B _13496_/B _13373_/D vssd1 vssd1 vccd1 vccd1 _13374_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_177_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10586_ _10586_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__xnor2_4
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15113_ _16115_/A _14848_/C _15110_/Y _15112_/Y _15109_/X vssd1 vssd1 vccd1 vccd1
+ _15113_/X sky130_fd_sc_hd__o311a_1
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12325_ _12325_/A _12325_/B _12325_/C vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__or3_1
XFILLER_103_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16093_ _15981_/B _15983_/B _15979_/Y vssd1 vssd1 vccd1 vccd1 _16095_/B sky130_fd_sc_hd__o21a_2
XFILLER_177_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15044_ _15041_/X _15042_/X _15043_/X vssd1 vssd1 vccd1 vccd1 _15044_/Y sky130_fd_sc_hd__a21oi_2
X_12256_ _12256_/A _12256_/B _12567_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12257_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_170_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11207_ _11175_/Y _11178_/Y _11206_/Y _10761_/A vssd1 vssd1 vccd1 vccd1 _11719_/A
+ sky130_fd_sc_hd__a211o_2
X_12187_ _12188_/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__nand2_2
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11138_ _11293_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11139_/C sky130_fd_sc_hd__and2_2
X_16995_ _16996_/B _16995_/B vssd1 vssd1 vccd1 vccd1 _16997_/A sky130_fd_sc_hd__and2b_1
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15946_ _16683_/A _16020_/B vssd1 vssd1 vccd1 vccd1 _16533_/B sky130_fd_sc_hd__and2_4
X_11069_ _11069_/A _11069_/B _11069_/C vssd1 vssd1 vccd1 vccd1 _11069_/X sky130_fd_sc_hd__or3_4
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15877_ _15877_/A _15877_/B _15875_/Y vssd1 vssd1 vccd1 vccd1 _15878_/B sky130_fd_sc_hd__or3b_1
XFILLER_23_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14828_ _14492_/A _14826_/X _14827_/Y _14597_/B vssd1 vssd1 vccd1 vccd1 _14828_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_184_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17547_ fanout934/X _17547_/D vssd1 vssd1 vccd1 vccd1 _17547_/Q sky130_fd_sc_hd__dfxtp_1
X_14759_ _14755_/A _14755_/B _14751_/A vssd1 vssd1 vccd1 vccd1 _14762_/A sky130_fd_sc_hd__o21a_1
XFILLER_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17478_ fanout926/X _17478_/D vssd1 vssd1 vccd1 vccd1 _17478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16429_ _16747_/A _16827_/B _16938_/B _16827_/A vssd1 vssd1 vccd1 vccd1 _16431_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout204 _17165_/A1 vssd1 vssd1 vccd1 vccd1 _16653_/A sky130_fd_sc_hd__buf_4
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout215 _17196_/X vssd1 vssd1 vccd1 vccd1 _17359_/B sky130_fd_sc_hd__buf_4
Xfanout226 _14933_/Y vssd1 vssd1 vccd1 vccd1 _16974_/B sky130_fd_sc_hd__buf_4
X_09803_ _10067_/A _09803_/B _09803_/C vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__and3_2
Xfanout237 _16218_/C1 vssd1 vssd1 vccd1 vccd1 _17074_/C1 sky130_fd_sc_hd__buf_4
XFILLER_141_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout248 _16007_/A vssd1 vssd1 vccd1 vccd1 _16304_/A sky130_fd_sc_hd__buf_6
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout259 _17295_/X vssd1 vssd1 vccd1 vccd1 _17359_/C sky130_fd_sc_hd__buf_4
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09734_ _09750_/C _10308_/B _09607_/A _09605_/Y vssd1 vssd1 vccd1 vccd1 _09735_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__xnor2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _10440_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__nand2_4
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10371_ _10383_/B _10383_/C _10383_/A vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__a21o_4
XFILLER_163_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12110_/A _12110_/B vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__xnor2_2
XFILLER_124_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _13220_/B _13090_/B vssd1 vssd1 vccd1 vccd1 _13092_/C sky130_fd_sc_hd__nand2_1
XFILLER_151_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ _15314_/A _14848_/A _12060_/S vssd1 vssd1 vccd1 vccd1 _12042_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout760 _10645_/C vssd1 vssd1 vccd1 vccd1 _10745_/D sky130_fd_sc_hd__buf_4
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout771 _10412_/C vssd1 vssd1 vccd1 vccd1 _10743_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_93_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15800_ _15797_/Y _15798_/Y _15799_/Y vssd1 vssd1 vccd1 vccd1 _15800_/Y sky130_fd_sc_hd__o21ai_1
Xfanout782 _10791_/D vssd1 vssd1 vccd1 vccd1 _09030_/D sky130_fd_sc_hd__buf_8
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16780_ _16781_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16846_/B sky130_fd_sc_hd__nor2_1
X_13992_ _14450_/A _14485_/D vssd1 vssd1 vccd1 vccd1 _14080_/C sky130_fd_sc_hd__and2_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout793 _13067_/C vssd1 vssd1 vccd1 vccd1 _13194_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_120_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15731_ _15732_/A _15732_/B vssd1 vssd1 vccd1 vccd1 _15731_/X sky130_fd_sc_hd__or2_1
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ _14771_/A _13866_/D vssd1 vssd1 vccd1 vccd1 _12945_/C sky130_fd_sc_hd__nand2_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15662_ _15662_/A _15774_/B vssd1 vssd1 vccd1 vccd1 _15663_/B sky130_fd_sc_hd__nand2_2
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _12875_/B _12875_/A vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__nand2b_2
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17401_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17401_/X sky130_fd_sc_hd__or2_1
X_14613_ _14567_/A _14567_/B _14566_/A vssd1 vssd1 vccd1 vccd1 _14615_/B sky130_fd_sc_hd__a21oi_1
X_11825_ _11841_/A _14848_/A _11595_/A vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__a21bo_2
X_15593_ _15594_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15595_/A sky130_fd_sc_hd__nand2_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14544_ _14593_/B _14545_/C _14545_/D _14593_/A vssd1 vssd1 vccd1 vccd1 _14548_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _12795_/B _17360_/A2 _17331_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17495_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _16568_/B sky130_fd_sc_hd__xor2_4
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10707_ _10708_/B _10708_/A vssd1 vssd1 vccd1 vccd1 _10715_/B sky130_fd_sc_hd__nand2b_2
X_14475_ _14475_/A vssd1 vssd1 vccd1 vccd1 _14533_/C sky130_fd_sc_hd__inv_2
X_17263_ _17455_/Q _17290_/A2 _17261_/X _17262_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1
+ _17455_/D sky130_fd_sc_hd__o221a_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11687_ _11688_/A _11688_/B vssd1 vssd1 vccd1 vccd1 _11692_/B sky130_fd_sc_hd__nand2_1
X_13426_ _13421_/Y _13422_/X _13308_/A _13309_/B vssd1 vssd1 vccd1 vccd1 _13428_/B
+ sky130_fd_sc_hd__o211a_1
X_16214_ _08760_/Y _14778_/X _14813_/X vssd1 vssd1 vccd1 vccd1 _16214_/Y sky130_fd_sc_hd__a21oi_1
X_17194_ input6/X input11/X input13/X input12/X vssd1 vssd1 vccd1 vccd1 _17195_/C
+ sky130_fd_sc_hd__or4_1
X_10638_ _11314_/A _11258_/B _10933_/D _10970_/B vssd1 vssd1 vccd1 vccd1 _10641_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16145_ _16146_/B _16146_/A vssd1 vssd1 vccd1 vccd1 _16145_/Y sky130_fd_sc_hd__nand2b_1
X_13357_ _13357_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__xnor2_2
X_10569_ _10672_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__and2_1
XFILLER_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12308_ _12309_/A _12309_/B _12309_/C vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__a21oi_4
XFILLER_115_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16076_ _16077_/A _16077_/B vssd1 vssd1 vccd1 vccd1 _16183_/B sky130_fd_sc_hd__and2_1
XFILLER_154_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13288_ _13286_/Y _13417_/A _17393_/A _13844_/D vssd1 vssd1 vccd1 vccd1 _13417_/B
+ sky130_fd_sc_hd__and4bb_2
X_15027_ _15024_/Y _15025_/Y _11480_/A vssd1 vssd1 vccd1 vccd1 _15687_/A sky130_fd_sc_hd__o21ai_4
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ _12239_/A _12239_/B vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__nor2_2
XFILLER_111_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16978_ _17140_/A _17028_/B _16973_/Y _16977_/X vssd1 vssd1 vccd1 vccd1 _16978_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 i_wb_addr[10] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_15929_ _15726_/A _15918_/A _16743_/C _17043_/B _15821_/X vssd1 vssd1 vccd1 vccd1
+ _15937_/A sky130_fd_sc_hd__a41o_1
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09450_ _09750_/C _10309_/B _09328_/A _09320_/Y vssd1 vssd1 vccd1 vccd1 _09451_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_188_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09381_ _09381_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__xnor2_1
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09717_ _09717_/A _09717_/B vssd1 vssd1 vccd1 vccd1 _09719_/B sky130_fd_sc_hd__xnor2_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _10560_/B _09647_/B _09647_/C vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__a21oi_2
XFILLER_167_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09579_ _09579_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09581_/C sky130_fd_sc_hd__or2_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__nand2_1
XFILLER_169_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12590_ _12592_/B _12592_/C _17139_/A _12592_/A vssd1 vssd1 vccd1 vccd1 _12593_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11541_ _11541_/A _11542_/A _11541_/C vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nor3_4
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _14257_/Y _14258_/X _14164_/X _14186_/A vssd1 vssd1 vccd1 vccd1 _14262_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_109_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11472_ _11472_/A _11472_/B _11471_/X vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__or3b_4
XFILLER_184_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13211_ _13211_/A _13339_/A _13211_/C vssd1 vssd1 vccd1 vccd1 _13339_/B sky130_fd_sc_hd__nor3_2
XFILLER_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ _10423_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__xnor2_4
X_14191_ _14192_/A _14192_/B _14192_/C vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__a21o_1
XFILLER_167_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ _13837_/A _12047_/X _12063_/C _12858_/Y vssd1 vssd1 vccd1 vccd1 _13142_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _10330_/B _10319_/C _10319_/D _10319_/A vssd1 vssd1 vccd1 vccd1 _10354_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_48_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13073_ _13244_/A _13073_/B vssd1 vssd1 vccd1 vccd1 _13075_/C sky130_fd_sc_hd__nor2_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10285_ _10188_/A _10188_/B _10188_/C vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__a21oi_4
X_16901_ _16900_/A _16900_/B _16900_/C vssd1 vssd1 vccd1 vccd1 _16902_/B sky130_fd_sc_hd__a21oi_2
X_12024_ _14952_/A _14949_/B _12053_/A vssd1 vssd1 vccd1 vccd1 _12024_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16832_ _16832_/A _16832_/B vssd1 vssd1 vccd1 vccd1 _16897_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout590 _12214_/A vssd1 vssd1 vccd1 vccd1 _12398_/S sky130_fd_sc_hd__buf_6
XFILLER_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16763_ _16764_/B _16763_/B vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__and2b_1
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13975_ _13867_/A _13869_/B _13867_/B vssd1 vssd1 vccd1 vccd1 _13982_/A sky130_fd_sc_hd__o21ba_4
XFILLER_47_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15714_ _10145_/B _15804_/A2 _15713_/X vssd1 vssd1 vccd1 vccd1 _15714_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12926_ _12926_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12928_/C sky130_fd_sc_hd__xnor2_2
X_16694_ _16777_/A _16694_/B vssd1 vssd1 vccd1 vccd1 _16701_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15645_ _15734_/A _15645_/B _16150_/B vssd1 vssd1 vccd1 vccd1 _15645_/Y sky130_fd_sc_hd__nor3_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _12382_/X _12398_/X _16011_/B vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__mux2_1
XFILLER_181_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _12021_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _14982_/C sky130_fd_sc_hd__and2_1
X_15576_ _15393_/B _15205_/B _15617_/A vssd1 vssd1 vccd1 vccd1 _16168_/B sky130_fd_sc_hd__a21bo_4
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _14771_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _12790_/C sky130_fd_sc_hd__nand2_1
XFILLER_187_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ input67/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17315_/X sky130_fd_sc_hd__or3_1
X_14527_ _14528_/A _14528_/B vssd1 vssd1 vccd1 vccd1 _14583_/B sky130_fd_sc_hd__or2_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11739_ _11739_/A _11739_/B _11739_/C vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__or3_4
XFILLER_187_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17246_ _17591_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17246_/X sky130_fd_sc_hd__a21o_1
X_14458_ _14528_/A _14458_/B vssd1 vssd1 vccd1 vccd1 _14459_/C sky130_fd_sc_hd__and2_2
XFILLER_128_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13409_ _13409_/A _13409_/B vssd1 vssd1 vccd1 vccd1 _13411_/C sky130_fd_sc_hd__xor2_4
X_14389_ _14389_/A _14389_/B vssd1 vssd1 vccd1 vccd1 _14456_/B sky130_fd_sc_hd__or2_2
XFILLER_128_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17177_ input30/X input32/X input31/X input34/X vssd1 vssd1 vccd1 vccd1 _17180_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_116_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16128_ _16807_/A _16127_/X _16126_/X vssd1 vssd1 vccd1 vccd1 _16130_/A sky130_fd_sc_hd__a21o_2
XFILLER_142_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08950_ _08950_/A _09065_/A vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__nor2_2
XFILLER_170_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16059_ _16165_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16060_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08881_ _08882_/A _08880_/Y _09025_/C _09555_/C vssd1 vssd1 vccd1 vccd1 _09027_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09502_ _09502_/A _17466_/D _09502_/C vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__and3_1
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__xnor2_4
XFILLER_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09364_/A _09364_/B vssd1 vssd1 vccd1 vccd1 _09497_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 _17444_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09295_ _09296_/A _09296_/B _09296_/C vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__a21o_4
XFILLER_178_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_31 _17443_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 _12592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _10839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_64 _17575_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_75 _17475_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_86 _10640_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_97 _13196_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__and2_2
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ _13761_/A _13761_/B vssd1 vssd1 vccd1 vccd1 _13762_/A sky130_fd_sc_hd__nor2_2
XFILLER_56_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ _10971_/A _10971_/B _14806_/A vssd1 vssd1 vccd1 vccd1 _10973_/B sky130_fd_sc_hd__a21oi_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _11849_/A _12707_/X _12710_/X _17165_/A1 vssd1 vssd1 vccd1 vccd1 _12711_/X
+ sky130_fd_sc_hd__a22o_2
X_13691_ _13895_/A _14318_/B _16722_/A _14213_/D vssd1 vssd1 vccd1 vccd1 _13793_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_44_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12642_ _12642_/A _12642_/B _12642_/C vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__or3_1
X_15430_ _16281_/A _15667_/B vssd1 vssd1 vccd1 vccd1 _15431_/B sky130_fd_sc_hd__nand2_2
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15361_ _15362_/B _15362_/A vssd1 vssd1 vccd1 vccd1 _15361_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12573_ _12425_/A _12427_/B _12425_/B vssd1 vssd1 vccd1 vccd1 _12583_/A sky130_fd_sc_hd__o21ba_2
XFILLER_178_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17100_ _14867_/A _17134_/C _17421_/A vssd1 vssd1 vccd1 vccd1 _17100_/X sky130_fd_sc_hd__and3b_1
X_14312_ _14312_/A _14312_/B vssd1 vssd1 vccd1 vccd1 _14313_/B sky130_fd_sc_hd__and2_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11524_ _11514_/A _11514_/C _11558_/A vssd1 vssd1 vccd1 vccd1 _11525_/C sky130_fd_sc_hd__o21ai_4
X_15292_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15295_/A sky130_fd_sc_hd__xnor2_4
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14243_ _14387_/A _14318_/C vssd1 vssd1 vccd1 vccd1 _14244_/B sky130_fd_sc_hd__nand2_2
X_17031_ _17023_/A _17163_/A2 _17030_/X vssd1 vssd1 vccd1 vccd1 _17033_/C sky130_fd_sc_hd__o21ba_1
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ _11451_/A _11451_/B _11495_/A vssd1 vssd1 vccd1 vccd1 _11456_/C sky130_fd_sc_hd__o21ba_4
XFILLER_184_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10406_ _10405_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10441_/B sky130_fd_sc_hd__and2b_4
X_14174_ _14252_/A _14174_/B vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__and2_4
XFILLER_152_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _11386_/A _11386_/B vssd1 vssd1 vccd1 vccd1 _11393_/A sky130_fd_sc_hd__xnor2_1
XFILLER_125_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13125_ _13125_/A _13125_/B _13125_/C vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__and3_4
XFILLER_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10337_ _10336_/A _10336_/Y _10215_/B _10228_/Y vssd1 vssd1 vccd1 vccd1 _10337_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13057_/A _13057_/B _13057_/C vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__o21a_2
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__xnor2_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12007_ _12007_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__xor2_4
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10199_ _10067_/A _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__a21oi_1
XFILLER_39_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _16108_/C _16589_/B _16813_/Y vssd1 vssd1 vccd1 vccd1 _16816_/C sky130_fd_sc_hd__a21o_1
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16746_ _16746_/A _16746_/B vssd1 vssd1 vccd1 vccd1 _16750_/A sky130_fd_sc_hd__xnor2_2
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _13958_/A _13958_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _13959_/B sky130_fd_sc_hd__nor3_1
XFILLER_46_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1044 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12909_ _12910_/A _12910_/B _12910_/C vssd1 vssd1 vccd1 vccd1 _13060_/A sky130_fd_sc_hd__o21ai_4
XFILLER_185_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16677_ _16676_/B _16677_/B vssd1 vssd1 vccd1 vccd1 _16678_/B sky130_fd_sc_hd__and2b_1
X_13889_ _13990_/A _13889_/B vssd1 vssd1 vccd1 vccd1 _13891_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15628_ _16012_/S _15628_/B vssd1 vssd1 vccd1 vccd1 _15628_/X sky130_fd_sc_hd__and2_1
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15559_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15675_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09080_ _09081_/A _09079_/Y _09750_/C _10180_/B vssd1 vssd1 vccd1 vccd1 _09306_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 i_wb_data[13] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
X_17229_ _17553_/Q _17229_/B vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__and2_1
XFILLER_190_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput51 i_wb_data[23] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_2
Xinput62 i_wb_data[4] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_2
XFILLER_162_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09982_ _09982_/A _10113_/A vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__nor2_4
XFILLER_171_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08933_ _09470_/A _09470_/B _12102_/D _12734_/C vssd1 vssd1 vccd1 vccd1 _08937_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _08796_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _11911_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09416_ _16983_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__xnor2_4
XFILLER_164_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09347_ _12546_/B _09350_/B _09161_/Y _09163_/B vssd1 vssd1 vccd1 vccd1 _09354_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_139_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09278_ _16982_/A _09273_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__o21ba_4
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _11240_/A _14785_/A _11423_/C _11605_/B vssd1 vssd1 vccd1 vccd1 _11306_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _11168_/Y _11169_/X _11021_/X _11041_/A vssd1 vssd1 vccd1 vccd1 _11171_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_162_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10122_ _10116_/A _10118_/B _10116_/B vssd1 vssd1 vccd1 vccd1 _10125_/A sky130_fd_sc_hd__o21ba_4
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10053_ _10053_/A _10053_/B _10053_/C vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__and3_4
XFILLER_88_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14930_ _17476_/D _17477_/D _14836_/B vssd1 vssd1 vccd1 vccd1 _14930_/Y sky130_fd_sc_hd__nor3b_2
X_14861_ _16571_/A _17497_/Q _16400_/B vssd1 vssd1 vccd1 vccd1 _16651_/B sky130_fd_sc_hd__and3_1
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16600_ _16600_/A _16600_/B vssd1 vssd1 vccd1 vccd1 _16601_/B sky130_fd_sc_hd__or2_1
X_13812_ _13812_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13814_/C sky130_fd_sc_hd__xor2_2
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17580_ fanout936/X _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14792_ _14792_/A _14792_/B vssd1 vssd1 vccd1 vccd1 _14796_/B sky130_fd_sc_hd__or2_2
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16531_ _16533_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16695_/C sky130_fd_sc_hd__nand2_1
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13743_ _13745_/B _13948_/C _13745_/D _13852_/A vssd1 vssd1 vccd1 vccd1 _13746_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10955_ _11010_/A vssd1 vssd1 vccd1 vccd1 _10955_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16462_ _16462_/A _16462_/B _16460_/Y vssd1 vssd1 vccd1 vccd1 _16463_/B sky130_fd_sc_hd__or3b_2
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ _14153_/B _16480_/A _13866_/C _14153_/A vssd1 vssd1 vccd1 vccd1 _13676_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ _11630_/A _11132_/C vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__nand2_1
X_15413_ _15660_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _15414_/B sky130_fd_sc_hd__nand2_4
XFILLER_176_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ _12626_/A _12626_/B _12626_/C vssd1 vssd1 vccd1 vccd1 _12820_/A sky130_fd_sc_hd__a21o_2
X_16393_ _16300_/A _16300_/B _16299_/B vssd1 vssd1 vccd1 vccd1 _16394_/B sky130_fd_sc_hd__o21ai_2
XFILLER_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12556_ _17401_/A _13450_/D vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__nand2_8
X_15344_ _15662_/A _15667_/B vssd1 vssd1 vccd1 vccd1 _15345_/B sky130_fd_sc_hd__nand2_4
XFILLER_157_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11507_ _11553_/A _14794_/B _11553_/D _11506_/A vssd1 vssd1 vccd1 vccd1 _11507_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15275_ _14881_/X _14889_/X _16595_/A _11841_/A vssd1 vssd1 vccd1 vccd1 _15277_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12487_ _12487_/A _12487_/B _12637_/D _12659_/B vssd1 vssd1 vccd1 vccd1 _12642_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_184_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17014_ _17014_/A _17014_/B _17014_/C vssd1 vssd1 vccd1 vccd1 _17016_/B sky130_fd_sc_hd__and3_1
X_14226_ _14226_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _16970_/A sky130_fd_sc_hd__nand2_8
XFILLER_176_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11438_ _11561_/B _11391_/B _11518_/C _11629_/A vssd1 vssd1 vccd1 vccd1 _11438_/Y
+ sky130_fd_sc_hd__a22oi_2
X_14157_ _14158_/A _14158_/B _14158_/C vssd1 vssd1 vccd1 vccd1 _14159_/A sky130_fd_sc_hd__o21a_1
X_11369_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__xnor2_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13109_/A _13109_/B vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__or2_2
X_14088_ _14088_/A _14088_/B vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__nand2_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13039_ _13040_/A _13040_/B _13040_/C vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__o21ai_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16729_ _13459_/A _16729_/B vssd1 vssd1 vccd1 vccd1 _16730_/B sky130_fd_sc_hd__nand2b_1
XFILLER_179_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09201_ _12488_/A _12338_/D _09196_/B _09193_/Y vssd1 vssd1 vccd1 vccd1 _09202_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_179_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09132_ _09360_/A _09172_/A _10067_/B _10446_/B vssd1 vssd1 vccd1 vccd1 _09135_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09063_ _09063_/A _09063_/B vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__xnor2_1
XFILLER_163_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09965_ _09966_/B _09966_/A vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__and2b_2
XFILLER_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08916_ _08916_/A _09057_/A vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _15537_/A _10309_/B _09890_/A _09756_/Y vssd1 vssd1 vccd1 vccd1 _09898_/C
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08847_ _11895_/A _12270_/B _12734_/D _12258_/B vssd1 vssd1 vccd1 vccd1 _08996_/A
+ sky130_fd_sc_hd__and4_2
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _12245_/A _11867_/D vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__nand2_2
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ _10647_/C _10647_/D _10648_/A _10646_/Y vssd1 vssd1 vccd1 vccd1 _10742_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _10671_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10672_/B sky130_fd_sc_hd__nand2_1
XFILLER_185_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12410_ _17401_/A _13866_/D _12238_/A _12236_/B vssd1 vssd1 vccd1 vccd1 _12412_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13390_ _12384_/X _12400_/B _13390_/S vssd1 vssd1 vccd1 vccd1 _13390_/X sky130_fd_sc_hd__mux2_4
XFILLER_154_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12341_ _12341_/A _12341_/B vssd1 vssd1 vccd1 vccd1 _12343_/C sky130_fd_sc_hd__xnor2_1
XFILLER_182_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ _15314_/A _15381_/A _15463_/A _15541_/A _15062_/S0 _12398_/S vssd1 vssd1
+ vccd1 vccd1 _15061_/B sky130_fd_sc_hd__mux4_1
X_12272_ _17375_/A _12752_/B vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__nand2_1
XFILLER_154_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _14011_/A _14011_/B vssd1 vssd1 vccd1 vccd1 _14013_/C sky130_fd_sc_hd__xnor2_2
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ _11223_/A _11223_/B vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__xor2_4
XFILLER_88_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11154_ _11154_/A _11155_/A _11154_/C vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__nor3_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10105_ _10005_/A _10005_/C _10005_/B vssd1 vssd1 vccd1 vccd1 _10105_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15962_ _15963_/A _15963_/B vssd1 vssd1 vccd1 vccd1 _15962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11085_ _11084_/A _11090_/A _11069_/X _11070_/Y vssd1 vssd1 vccd1 vccd1 _11087_/A
+ sky130_fd_sc_hd__o211a_1
X_10036_ _10525_/A _10036_/B _10534_/D _10036_/D vssd1 vssd1 vccd1 vccd1 _10039_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14913_ _12054_/A _10791_/C _10991_/C vssd1 vssd1 vccd1 vccd1 _14913_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15893_ _15890_/X _15891_/X _15892_/Y vssd1 vssd1 vccd1 vccd1 _15893_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14844_ _14929_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _14844_/X sky130_fd_sc_hd__or2_1
XFILLER_17_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17563_ fanout941/X _17563_/D vssd1 vssd1 vccd1 vccd1 _17563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14775_ _14775_/A _17497_/Q vssd1 vssd1 vccd1 vccd1 _14775_/X sky130_fd_sc_hd__or2_2
X_11987_ _11987_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _11988_/B sky130_fd_sc_hd__nor2_4
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _16827_/B _16938_/B _16514_/C vssd1 vssd1 vccd1 vccd1 _16515_/B sky130_fd_sc_hd__or3_1
XFILLER_1_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13726_ _13726_/A _13726_/B vssd1 vssd1 vccd1 vccd1 _13727_/B sky130_fd_sc_hd__and2_1
XFILLER_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10938_ _10938_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10940_/B sky130_fd_sc_hd__xor2_4
X_17494_ fanout930/X _17494_/D vssd1 vssd1 vccd1 vccd1 _17494_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16445_ _16619_/A _16681_/D vssd1 vssd1 vccd1 vccd1 _16533_/C sky130_fd_sc_hd__nor2_1
X_13657_ _13541_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13658_/C sky130_fd_sc_hd__nand2b_1
X_10869_ _14787_/A _11561_/C _15175_/B _14786_/A vssd1 vssd1 vccd1 vccd1 _10870_/B
+ sky130_fd_sc_hd__a22oi_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12608_ _12778_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12610_/B sky130_fd_sc_hd__nand2_2
X_16376_ _16280_/B _16282_/B _16280_/A vssd1 vssd1 vccd1 vccd1 _16378_/B sky130_fd_sc_hd__o21ba_2
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _13469_/A _13471_/B _13469_/B vssd1 vssd1 vccd1 vccd1 _13589_/B sky130_fd_sc_hd__o21ba_2
XFILLER_185_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15327_ _14882_/X _15325_/X _17377_/A vssd1 vssd1 vccd1 vccd1 _15327_/X sky130_fd_sc_hd__a21o_1
X_12539_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12539_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15258_ _16389_/A _15235_/Y _15236_/X _15257_/X vssd1 vssd1 vccd1 vccd1 _15258_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14209_ _12388_/X _12401_/B _14839_/A vssd1 vssd1 vccd1 vccd1 _14209_/X sky130_fd_sc_hd__mux2_2
XFILLER_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15189_ _15131_/A _14921_/X _15254_/S vssd1 vssd1 vccd1 vccd1 _15189_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout408 _17529_/Q vssd1 vssd1 vccd1 vccd1 _09409_/C sky130_fd_sc_hd__buf_2
Xfanout419 _14776_/A vssd1 vssd1 vccd1 vccd1 _13948_/B sky130_fd_sc_hd__buf_4
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _09751_/A _09749_/Y _09750_/C _10657_/B vssd1 vssd1 vccd1 vccd1 _09880_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09681_ _09681_/A _09681_/B vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__or2_2
XFILLER_95_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09115_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09119_/C sky130_fd_sc_hd__or3_4
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_967 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ _09047_/B _09047_/A vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__nand2b_2
XFILLER_191_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout920 _08730_/Y vssd1 vssd1 vccd1 vccd1 _17322_/C1 sky130_fd_sc_hd__buf_4
XFILLER_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout931 fanout937/X vssd1 vssd1 vccd1 vccd1 fanout931/X sky130_fd_sc_hd__clkbuf_4
Xfanout942 fanout943/X vssd1 vssd1 vccd1 vccd1 fanout942/X sky130_fd_sc_hd__buf_4
X_09948_ _09948_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__xnor2_2
XTAP_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09879_ _09750_/C _10657_/B _09751_/A _09749_/Y vssd1 vssd1 vccd1 vccd1 _09880_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11911_/A _11911_/B _11911_/C vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__a21o_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _13658_/A _13298_/A _13908_/B _13903_/B vssd1 vssd1 vccd1 vccd1 _13043_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__and2_2
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _14560_/A _14560_/B vssd1 vssd1 vccd1 vccd1 _14562_/C sky130_fd_sc_hd__xor2_2
X_11772_ _11771_/A _16972_/A _16972_/B _11770_/Y vssd1 vssd1 vccd1 vccd1 _11773_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10723_ _11260_/C _10640_/D _10641_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _10724_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13511_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13511_/X sky130_fd_sc_hd__and2_2
X_14491_ _14599_/B _14641_/C vssd1 vssd1 vccd1 vccd1 _14492_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16126_/X _16130_/B _16127_/X _16807_/A vssd1 vssd1 vccd1 vccd1 _16232_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_13442_ _13442_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13443_/C sky130_fd_sc_hd__xnor2_2
X_10654_ _10993_/C _10545_/D _10546_/A _10544_/Y vssd1 vssd1 vccd1 vccd1 _10655_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_186_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _16161_/A _16161_/B vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__xnor2_4
X_13373_ _13494_/A _13373_/B _13496_/B _13373_/D vssd1 vssd1 vccd1 vccd1 _13494_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_186_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ _10573_/X _10574_/Y _10567_/A _10572_/A vssd1 vssd1 vccd1 vccd1 _10585_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_177_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ _14791_/X _15899_/A2 _15111_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15112_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12324_ _12324_/A _12492_/B vssd1 vssd1 vccd1 vccd1 _12325_/C sky130_fd_sc_hd__nor2_1
XFILLER_186_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16092_ _16092_/A _16092_/B vssd1 vssd1 vccd1 vccd1 _16095_/A sky130_fd_sc_hd__xnor2_4
XFILLER_103_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12255_ _12088_/B _12567_/B _12565_/C _12256_/A vssd1 vssd1 vccd1 vccd1 _12257_/A
+ sky130_fd_sc_hd__a22oi_4
X_15043_ _14941_/X _15003_/X _15002_/X vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__a21bo_2
XFILLER_108_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11206_ _10760_/A _10760_/B _10760_/C vssd1 vssd1 vccd1 vccd1 _11206_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12186_ _12186_/A _12186_/B vssd1 vssd1 vccd1 vccd1 _12188_/B sky130_fd_sc_hd__xor2_2
XFILLER_79_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11137_ _11137_/A _11137_/B _11137_/C vssd1 vssd1 vccd1 vccd1 _11138_/B sky130_fd_sc_hd__or3_1
XFILLER_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16994_ _16994_/A _16994_/B vssd1 vssd1 vccd1 vccd1 _16995_/B sky130_fd_sc_hd__and2_1
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15945_ _15859_/A _15859_/B _15857_/X vssd1 vssd1 vccd1 vccd1 _15969_/A sky130_fd_sc_hd__o21ai_1
XFILLER_62_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11068_ _11055_/X _11056_/Y _11065_/B _11065_/Y vssd1 vssd1 vccd1 vccd1 _11069_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10019_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__xnor2_4
XFILLER_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15876_ _15877_/A _15877_/B _15875_/Y vssd1 vssd1 vccd1 vccd1 _15992_/A sky130_fd_sc_hd__o21ba_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14827_ _17421_/A _14867_/A vssd1 vssd1 vccd1 vccd1 _14827_/Y sky130_fd_sc_hd__nor2_2
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17546_ fanout946/X _17546_/D vssd1 vssd1 vccd1 vccd1 _17546_/Q sky130_fd_sc_hd__dfxtp_4
X_14758_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14758_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13709_ _13706_/Y _13707_/X _13594_/X _13598_/A vssd1 vssd1 vccd1 vccd1 _13710_/D
+ sky130_fd_sc_hd__a211oi_4
X_17477_ fanout929/X _17477_/D vssd1 vssd1 vccd1 vccd1 _17477_/Q sky130_fd_sc_hd__dfxtp_4
X_14689_ _14717_/A _14689_/B vssd1 vssd1 vccd1 vccd1 _14691_/B sky130_fd_sc_hd__nand2_1
X_16428_ _16324_/A _16326_/B _16324_/B vssd1 vssd1 vccd1 vccd1 _16436_/A sky130_fd_sc_hd__a21bo_4
XFILLER_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _16443_/A _16359_/B vssd1 vssd1 vccd1 vccd1 _16361_/B sky130_fd_sc_hd__and2_2
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 _11849_/Y vssd1 vssd1 vccd1 vccd1 _17165_/A1 sky130_fd_sc_hd__buf_4
Xfanout216 _17196_/X vssd1 vssd1 vccd1 vccd1 _17355_/B sky130_fd_sc_hd__buf_2
XFILLER_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09802_ _09805_/B _09802_/B vssd1 vssd1 vccd1 vccd1 _09803_/C sky130_fd_sc_hd__nor2_1
Xfanout227 _14933_/Y vssd1 vssd1 vccd1 vccd1 _16733_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 _16218_/C1 vssd1 vssd1 vccd1 vccd1 _14944_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_87_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout249 _15108_/A vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__buf_6
XFILLER_87_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09733_ _09733_/A _09733_/B vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09664_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__or2_1
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09595_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ _10709_/A _10370_/B _10370_/C vssd1 vssd1 vccd1 vccd1 _10383_/C sky130_fd_sc_hd__or3_4
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09029_ _11867_/B _12637_/D _09030_/D _09030_/A vssd1 vssd1 vccd1 vccd1 _09031_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_123_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ _14911_/B _12040_/B vssd1 vssd1 vccd1 vccd1 _12040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout750 _10899_/D vssd1 vssd1 vccd1 vccd1 _10647_/D sky130_fd_sc_hd__buf_6
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout761 _10897_/B vssd1 vssd1 vccd1 vccd1 _10645_/C sky130_fd_sc_hd__buf_6
Xfanout772 _13196_/B vssd1 vssd1 vccd1 vccd1 _10412_/C sky130_fd_sc_hd__clkbuf_4
X_13991_ _13895_/B _14485_/D _16859_/A _13895_/A vssd1 vssd1 vccd1 vccd1 _13991_/X
+ sky130_fd_sc_hd__a22o_1
Xfanout783 _10791_/D vssd1 vssd1 vccd1 vccd1 _11132_/C sky130_fd_sc_hd__buf_6
XFILLER_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout794 _17489_/Q vssd1 vssd1 vccd1 vccd1 _13067_/C sky130_fd_sc_hd__buf_6
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15730_ _15730_/A _15730_/B vssd1 vssd1 vccd1 vccd1 _15732_/B sky130_fd_sc_hd__xnor2_4
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _17413_/A _17411_/A _13229_/B _13100_/B vssd1 vssd1 vccd1 vccd1 _13085_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15661_ _15661_/A _15661_/B vssd1 vssd1 vccd1 vccd1 _15663_/A sky130_fd_sc_hd__xnor2_4
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12715_/A _12717_/B _12715_/B vssd1 vssd1 vccd1 vccd1 _12875_/B sky130_fd_sc_hd__o21ba_2
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ input45/X _17422_/A2 _17399_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17528_/D
+ sky130_fd_sc_hd__o211a_1
X_14612_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14614_/B sky130_fd_sc_hd__xnor2_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11824_ _12700_/D _11824_/B vssd1 vssd1 vccd1 vccd1 _11824_/Y sky130_fd_sc_hd__nand2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15278_/A _16812_/A _15498_/A _15496_/A vssd1 vssd1 vccd1 vccd1 _15594_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ input44/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17331_/X sky130_fd_sc_hd__or3_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _16653_/A _14543_/B vssd1 vssd1 vccd1 vccd1 _14543_/Y sky130_fd_sc_hd__nand2_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11759_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11756_/B sky130_fd_sc_hd__and2b_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17564_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__and2_1
XFILLER_144_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ _11030_/A _10705_/B _10705_/A vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__o21ba_2
X_14474_ _14473_/A _14473_/B _14473_/C vssd1 vssd1 vccd1 vccd1 _14475_/A sky130_fd_sc_hd__a21oi_4
XFILLER_187_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _11686_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__xnor2_2
XFILLER_146_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16213_ _16107_/Y _16111_/B _16210_/Y _16917_/A vssd1 vssd1 vccd1 vccd1 _16213_/X
+ sky130_fd_sc_hd__o31a_1
X_13425_ _13428_/A vssd1 vssd1 vccd1 vccd1 _13425_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_186_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17193_ input32/X input31/X input33/X input7/X vssd1 vssd1 vccd1 vccd1 _17195_/B
+ sky130_fd_sc_hd__or4_1
X_10637_ _10637_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__xnor2_4
XFILLER_167_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _16035_/A _16035_/B _16027_/Y vssd1 vssd1 vccd1 vccd1 _16146_/B sky130_fd_sc_hd__o21a_4
XFILLER_128_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _13357_/A _13357_/B vssd1 vssd1 vccd1 vccd1 _13477_/A sky130_fd_sc_hd__and2b_1
X_10568_ _10672_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__nor2_4
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _12307_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12309_/C sky130_fd_sc_hd__xnor2_4
X_16075_ _16075_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _16077_/B sky130_fd_sc_hd__xnor2_1
XFILLER_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13287_ _13852_/A _13745_/B _14002_/B _13523_/B vssd1 vssd1 vccd1 vccd1 _13417_/A
+ sky130_fd_sc_hd__and4_2
X_10499_ _10499_/A vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _15024_/Y _15025_/Y _11480_/A vssd1 vssd1 vccd1 vccd1 _15872_/A sky130_fd_sc_hd__o21a_4
XFILLER_142_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12238_ _12238_/A _12238_/B vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__xnor2_4
XFILLER_151_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12169_ _12169_/A _12169_/B _12169_/C vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__and3_1
XFILLER_25_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16977_ _16977_/A _16977_/B _16977_/C vssd1 vssd1 vccd1 vccd1 _16977_/X sky130_fd_sc_hd__and3_1
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 i_wb_addr[11] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15928_ _15832_/A _15829_/X _15831_/B vssd1 vssd1 vccd1 vccd1 _15939_/A sky130_fd_sc_hd__o21ai_1
XFILLER_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15859_ _15859_/A _15859_/B vssd1 vssd1 vccd1 vccd1 _15861_/B sky130_fd_sc_hd__xor2_4
XFILLER_149_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09380_ _09381_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__and2b_1
XFILLER_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17529_ fanout932/X _17529_/D vssd1 vssd1 vccd1 vccd1 _17529_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09716_ _09717_/B _09717_/A vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__nand2b_2
XFILLER_68_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09647_ _10560_/B _09647_/B _09647_/C vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__and3_2
XFILLER_167_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__nor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11540_ _11539_/A _11539_/B _11538_/X vssd1 vssd1 vccd1 vccd1 _11541_/C sky130_fd_sc_hd__o21ba_2
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11471_ _11553_/A _14792_/B _11506_/C _11506_/A vssd1 vssd1 vccd1 vccd1 _11471_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ _13211_/A _13339_/A _13211_/C vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__o21a_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10422_ _10422_/A _10531_/A vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__or2_4
X_14190_ _14190_/A _14190_/B vssd1 vssd1 vccd1 vccd1 _14192_/C sky130_fd_sc_hd__xnor2_1
XFILLER_167_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10353_ _10336_/A _10336_/C _10336_/B vssd1 vssd1 vccd1 vccd1 _10353_/X sky130_fd_sc_hd__o21a_2
X_13141_ _16922_/A _13139_/X _13140_/Y _13013_/Y _13016_/X vssd1 vssd1 vccd1 vccd1
+ _17584_/D sky130_fd_sc_hd__a32o_1
XFILLER_174_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13072_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13073_/B sky130_fd_sc_hd__nor3_1
XFILLER_151_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10284_ _10263_/X _10283_/X _10157_/Y _10230_/X vssd1 vssd1 vccd1 vccd1 _10319_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_970 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16900_ _16900_/A _16900_/B _16900_/C vssd1 vssd1 vccd1 vccd1 _16902_/A sky130_fd_sc_hd__and3_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12023_ _17363_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _14949_/B sky130_fd_sc_hd__and2_1
X_16831_ _16832_/A _16832_/B vssd1 vssd1 vccd1 vccd1 _16833_/A sky130_fd_sc_hd__and2_1
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout580 _14922_/S vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__buf_4
Xfanout591 _14794_/A vssd1 vssd1 vccd1 vccd1 _10993_/C sky130_fd_sc_hd__buf_4
X_16762_ _16762_/A _16762_/B vssd1 vssd1 vccd1 vccd1 _16763_/B sky130_fd_sc_hd__xor2_1
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13974_ _13974_/A _13974_/B vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__xnor2_4
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15713_ _15707_/B _15899_/A2 _15713_/B1 _15709_/A _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15713_/X sky130_fd_sc_hd__a221o_1
X_12925_ _17421_/A _13067_/C vssd1 vssd1 vccd1 vccd1 _12926_/B sky130_fd_sc_hd__nand2_2
X_16693_ _16692_/B _16693_/B vssd1 vssd1 vccd1 vccd1 _16694_/B sky130_fd_sc_hd__nand2b_1
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15644_ _15821_/A _16604_/B _15551_/Y _15918_/A vssd1 vssd1 vccd1 vccd1 _15644_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _12856_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _17582_/D sky130_fd_sc_hd__nand2_1
XFILLER_62_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _14912_/B _11807_/B vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__nand2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15575_ _15393_/B _15205_/B _15617_/A vssd1 vssd1 vccd1 vccd1 _15575_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _14769_/A _14770_/A _13100_/B _13551_/D vssd1 vssd1 vccd1 vccd1 _12947_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _12770_/D _17328_/A2 _17313_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17486_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14526_ _14583_/A _14526_/B vssd1 vssd1 vccd1 vccd1 _14528_/B sky130_fd_sc_hd__nand2_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11738_ _11736_/A _11736_/B _11735_/Y vssd1 vssd1 vccd1 vccd1 _11739_/C sky130_fd_sc_hd__o21ba_1
XFILLER_175_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17245_ _17449_/Q _17290_/A2 _17243_/X _17244_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17449_/D sky130_fd_sc_hd__o221a_1
XFILLER_31_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ _14456_/A _14456_/B _14456_/C vssd1 vssd1 vccd1 vccd1 _14458_/B sky130_fd_sc_hd__a21o_1
XFILLER_70_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11669_ _15524_/C _11670_/C vssd1 vssd1 vccd1 vccd1 _11690_/B sky130_fd_sc_hd__and2b_1
XFILLER_128_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ _13408_/A _13408_/B vssd1 vssd1 vccd1 vccd1 _13409_/B sky130_fd_sc_hd__xnor2_4
XFILLER_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17176_ input33/X input5/X input4/X input7/X vssd1 vssd1 vccd1 vccd1 _17180_/A sky130_fd_sc_hd__or4_1
X_14388_ _14388_/A _14388_/B vssd1 vssd1 vccd1 vccd1 _14456_/A sky130_fd_sc_hd__xnor2_4
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16127_ _16127_/A _16127_/B _17119_/C vssd1 vssd1 vccd1 vccd1 _16127_/X sky130_fd_sc_hd__and3_1
X_13339_ _13339_/A _13339_/B _13339_/C vssd1 vssd1 vccd1 vccd1 _13341_/A sky130_fd_sc_hd__or3_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16058_ _16058_/A _16058_/B vssd1 vssd1 vccd1 vccd1 _16060_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15009_ _15248_/C _14846_/B _15008_/X _16008_/B1 _15008_/A vssd1 vssd1 vccd1 vccd1
+ _15009_/X sky130_fd_sc_hd__a32o_1
XFILLER_29_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08880_ _09023_/B _09414_/C _09509_/B _09023_/A vssd1 vssd1 vccd1 vccd1 _08880_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_9_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09501_ _09502_/A _10062_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09432_ _09433_/B _09433_/A vssd1 vssd1 vccd1 vccd1 _09441_/B sky130_fd_sc_hd__nand2b_2
XFILLER_25_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _09502_/A _10067_/B _09357_/A _09174_/Y vssd1 vssd1 vccd1 vccd1 _09364_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09294_ _09294_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09296_/C sky130_fd_sc_hd__or2_2
XANTENNA_10 _17534_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_21 _17446_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _16352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 _15396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 _11268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_65 _17575_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_76 _17542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_87 _08969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10971_ _10971_/A _10971_/B _14806_/A vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__and3_1
XFILLER_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _15457_/B _12710_/B vssd1 vssd1 vccd1 vccd1 _12710_/X sky130_fd_sc_hd__or2_1
XFILLER_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ _14318_/B _16722_/A _14213_/D _13895_/A vssd1 vssd1 vccd1 vccd1 _13693_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_188_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12641_/A _12792_/B vssd1 vssd1 vccd1 vccd1 _12642_/C sky130_fd_sc_hd__nor2_2
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15360_ _15292_/A _15292_/B _15286_/Y vssd1 vssd1 vccd1 vccd1 _15362_/B sky130_fd_sc_hd__a21oi_2
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12572_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__or3_2
XFILLER_184_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14311_ _14312_/A _14312_/B vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__nor2_1
XFILLER_178_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _11523_/A _11523_/B vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__xnor2_4
XFILLER_156_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15291_ _15291_/A _15291_/B vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__xnor2_4
XFILLER_184_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17030_ _17023_/B _17162_/A2 _16974_/B _17028_/A _17170_/B1 vssd1 vssd1 vccd1 vccd1
+ _17030_/X sky130_fd_sc_hd__a221o_1
X_14242_ _14242_/A _14242_/B vssd1 vssd1 vccd1 vccd1 _14244_/A sky130_fd_sc_hd__nor2_1
X_11454_ _11460_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11456_/B sky130_fd_sc_hd__nand2_4
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _10405_/A _10405_/B _10405_/C _10405_/D vssd1 vssd1 vccd1 vccd1 _10406_/B
+ sky130_fd_sc_hd__or4_4
X_14173_ _14173_/A _14173_/B _14173_/C vssd1 vssd1 vccd1 vccd1 _14174_/B sky130_fd_sc_hd__or3_1
X_11385_ _11395_/B _11435_/A _11395_/A vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__a21o_1
XFILLER_139_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13124_ _13125_/A _13125_/B _13125_/C vssd1 vssd1 vccd1 vccd1 _13258_/A sky130_fd_sc_hd__a21oi_4
X_10336_ _10336_/A _10336_/B _10336_/C vssd1 vssd1 vccd1 vccd1 _10336_/Y sky130_fd_sc_hd__nor3_4
XFILLER_180_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13055_ _13055_/A _13055_/B vssd1 vssd1 vccd1 vccd1 _13057_/C sky130_fd_sc_hd__xor2_2
X_10267_ _10267_/A _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10267_/Y sky130_fd_sc_hd__nand3_2
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12006_ _12007_/A _12007_/B vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__and2_1
XFILLER_79_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10198_ _10198_/A _10322_/A _10198_/C vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__or3_1
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814_ _16814_/A _16814_/B _16938_/D _16883_/C vssd1 vssd1 vccd1 vccd1 _16888_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16745_ _16938_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16746_/B sky130_fd_sc_hd__nand2_1
X_13957_ _13958_/A _13958_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _14044_/B sky130_fd_sc_hd__o21a_1
X_12908_ _12908_/A _12908_/B vssd1 vssd1 vccd1 vccd1 _12910_/C sky130_fd_sc_hd__xnor2_4
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16676_ _16677_/B _16676_/B vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__and2b_1
XFILLER_146_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13888_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _13889_/B sky130_fd_sc_hd__and2_1
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15627_ _16011_/A _15627_/B vssd1 vssd1 vccd1 vccd1 _15628_/B sky130_fd_sc_hd__or2_2
X_12839_ _12689_/A _12691_/A _13001_/B _12837_/Y vssd1 vssd1 vccd1 vccd1 _12840_/B
+ sky130_fd_sc_hd__o211ai_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15558_ _15559_/A _15559_/B vssd1 vssd1 vccd1 vccd1 _15558_/Y sky130_fd_sc_hd__nor2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14509_ _14509_/A _14509_/B _14509_/C vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__nor3_2
XFILLER_159_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15489_ _15489_/A _15489_/B vssd1 vssd1 vccd1 vccd1 _15499_/A sky130_fd_sc_hd__xor2_4
X_17228_ _17585_/Q _17270_/A2 _17270_/B1 vssd1 vssd1 vccd1 vccd1 _17228_/X sky130_fd_sc_hd__a21o_1
Xinput30 i_wb_addr[5] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput41 i_wb_data[14] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput52 i_wb_data[24] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput63 i_wb_data[5] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17159_ _11778_/Y _17157_/Y _17158_/Y vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__o21ai_4
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09981_ _09982_/A _09980_/Y _09981_/C _17469_/D vssd1 vssd1 vccd1 vccd1 _10113_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08932_ _08872_/X _08874_/X _08930_/A _08929_/Y vssd1 vssd1 vccd1 vccd1 _09016_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08863_ _08864_/B _08864_/A vssd1 vssd1 vccd1 vccd1 _08863_/X sky130_fd_sc_hd__and2b_2
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08794_ _11878_/B _08794_/B vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__nor2_2
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09415_ _09415_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__nor2_2
XFILLER_52_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__or2_2
XFILLER_139_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _09290_/B _09290_/C _09290_/A vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__a21o_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11170_ _11021_/X _11041_/A _11168_/Y _11169_/X vssd1 vssd1 vccd1 vccd1 _11202_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_134_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10121_ _10133_/B _10133_/C _10133_/A vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__a21o_4
XFILLER_171_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10052_ _10074_/B _10052_/B vssd1 vssd1 vccd1 vccd1 _10053_/C sky130_fd_sc_hd__and2_2
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14860_ _16399_/A _16399_/B vssd1 vssd1 vccd1 vccd1 _16400_/B sky130_fd_sc_hd__and2_2
XFILLER_76_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _13812_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13921_/B sky130_fd_sc_hd__or2_1
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14791_ _14791_/A _15116_/B vssd1 vssd1 vccd1 vccd1 _14791_/X sky130_fd_sc_hd__or2_2
XFILLER_29_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16530_ _16437_/A _16437_/B _16435_/X vssd1 vssd1 vccd1 vccd1 _16543_/A sky130_fd_sc_hd__a21o_1
X_13742_ _13742_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__nor2_4
X_10954_ _11006_/A _11006_/B _11097_/D _11027_/C vssd1 vssd1 vccd1 vccd1 _11010_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16461_ _16462_/A _16462_/B _16460_/Y vssd1 vssd1 vccd1 vccd1 _16557_/A sky130_fd_sc_hd__o21ba_2
X_13673_ _13670_/Y _13770_/B _13558_/A _13559_/Y vssd1 vssd1 vccd1 vccd1 _13710_/B
+ sky130_fd_sc_hd__o211a_2
X_10885_ _11561_/A _11629_/B _10932_/B _11135_/B vssd1 vssd1 vccd1 vccd1 _10891_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15412_ _15948_/A _15932_/A vssd1 vssd1 vccd1 vccd1 _15414_/A sky130_fd_sc_hd__nor2_4
X_12624_ _12780_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _12626_/C sky130_fd_sc_hd__nand2_1
X_16392_ _14776_/A _16391_/Y _16390_/Y vssd1 vssd1 vccd1 vccd1 _16396_/A sky130_fd_sc_hd__a21o_1
XFILLER_106_1010 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15343_ _15342_/A _15661_/A _15340_/X vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__a21oi_4
X_12555_ _12542_/Y _12555_/B vssd1 vssd1 vccd1 vccd1 _17580_/D sky130_fd_sc_hd__nand2b_1
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1054 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A _11553_/A _11506_/C _11553_/D vssd1 vssd1 vccd1 vccd1 _11506_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_129_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15274_ _15274_/A _15948_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__or3b_4
XFILLER_157_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12486_ _12487_/B _12637_/D _12659_/B _12487_/A vssd1 vssd1 vccd1 vccd1 _12490_/A
+ sky130_fd_sc_hd__a22oi_4
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _17014_/C sky130_fd_sc_hd__clkinv_2
X_14225_ _14225_/A _14225_/B vssd1 vssd1 vccd1 vccd1 _14227_/A sky130_fd_sc_hd__nor2_1
X_11437_ _11629_/A _11437_/B _14897_/A _11518_/C vssd1 vssd1 vccd1 vccd1 _11440_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_171_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14156_ _14156_/A _14156_/B vssd1 vssd1 vccd1 vccd1 _14158_/C sky130_fd_sc_hd__xnor2_2
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11368_ _11367_/A _11367_/C _11448_/A vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _13107_/A _13107_/B vssd1 vssd1 vccd1 vccd1 _13109_/B sky130_fd_sc_hd__nor2_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10319_/A _10330_/B _10319_/C _10319_/D vssd1 vssd1 vccd1 vccd1 _10319_/Y
+ sky130_fd_sc_hd__nand4_4
X_14087_ _14086_/B _14087_/B vssd1 vssd1 vccd1 vccd1 _14088_/B sky130_fd_sc_hd__nand2b_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11299_ _11299_/A _11299_/B _11299_/C vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__or3_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13038_/A _13038_/B vssd1 vssd1 vccd1 vccd1 _13040_/C sky130_fd_sc_hd__xnor2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14989_ _14986_/Y _14988_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _14989_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16728_ _16727_/B _16728_/B vssd1 vssd1 vccd1 vccd1 _16728_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_62_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16659_ _17063_/A _16639_/Y _16658_/X vssd1 vssd1 vccd1 vccd1 _16659_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09200_ _09227_/B _09200_/B vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__and2_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09131_ _09167_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__and2_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09062_ _09063_/B _09063_/A vssd1 vssd1 vccd1 vccd1 _09062_/X sky130_fd_sc_hd__and2b_2
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09964_ _09964_/A _10091_/A vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__nor2_1
XFILLER_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ _08916_/A _08914_/Y _17381_/A _12565_/D vssd1 vssd1 vccd1 vccd1 _09057_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _09895_/A _10021_/A vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _12270_/B _12734_/D _12258_/B _11895_/A vssd1 vssd1 vccd1 vccd1 _08846_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__nor2_4
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10670_ _10670_/A _10670_/B vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__nand2_4
XFILLER_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09332_/B _09329_/B vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__and2_1
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _12659_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__nand2_1
X_12271_ _12271_/A _12271_/B vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__nor2_1
XFILLER_182_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _14115_/B _14010_/B vssd1 vssd1 vccd1 vccd1 _14011_/B sky130_fd_sc_hd__and2_1
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11222_ _11222_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11223_/B sky130_fd_sc_hd__or2_4
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1003 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11153_ _11153_/A _11153_/B _11153_/C vssd1 vssd1 vccd1 vccd1 _11154_/C sky130_fd_sc_hd__nor3_2
XFILLER_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10104_ _10027_/B _10027_/C _10025_/Y _10028_/A vssd1 vssd1 vccd1 vccd1 _10104_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_95_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15961_ _15855_/A _15855_/B _15852_/Y vssd1 vssd1 vccd1 vccd1 _15963_/B sky130_fd_sc_hd__o21a_2
X_11084_ _11084_/A _11084_/B _11084_/C vssd1 vssd1 vccd1 vccd1 _11090_/A sky130_fd_sc_hd__nor3_4
XFILLER_89_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10035_ _10035_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14912_ _12104_/A _14912_/B vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_103_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15892_ _15797_/Y _15798_/Y _15797_/A vssd1 vssd1 vccd1 vccd1 _15892_/Y sky130_fd_sc_hd__o21ai_2
X_14843_ _14929_/A _14938_/B vssd1 vssd1 vccd1 vccd1 _15248_/C sky130_fd_sc_hd__nor2_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17562_ fanout945/X _17562_/D vssd1 vssd1 vccd1 vccd1 _17562_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _14774_/A _16571_/A vssd1 vssd1 vccd1 vccd1 _16576_/B sky130_fd_sc_hd__or2_1
X_11986_ _11985_/B _11986_/B vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__and2b_1
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16513_ _16827_/B _16938_/B _16514_/C vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__o21ai_1
XFILLER_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13725_ _13726_/A _13726_/B vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10937_ _10938_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__nand2_2
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17493_ fanout930/X _17493_/D vssd1 vssd1 vccd1 vccd1 _17493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16444_ _16444_/A _16444_/B vssd1 vssd1 vccd1 vccd1 _16455_/A sky130_fd_sc_hd__or2_2
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13656_ _13654_/X _13656_/B vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__nand2b_1
X_10868_ _14788_/A _15314_/A vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__nand2_4
XFILLER_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ _12607_/A _12607_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__or3_1
X_16375_ _16375_/A _16375_/B vssd1 vssd1 vccd1 vccd1 _16378_/A sky130_fd_sc_hd__xnor2_4
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13587_ _13587_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13589_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10799_ _14787_/A _15381_/A vssd1 vssd1 vccd1 vccd1 _10799_/Y sky130_fd_sc_hd__nand2_2
X_15326_ _14882_/X _15325_/X _17377_/A vssd1 vssd1 vccd1 vccd1 _16695_/A sky130_fd_sc_hd__a21oi_4
XFILLER_118_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12538_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15257_ _15257_/A _15257_/B _15257_/C _15256_/X vssd1 vssd1 vccd1 vccd1 _15257_/X
+ sky130_fd_sc_hd__or4b_2
X_12469_ _12271_/A _12273_/B _12271_/B vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__o21ba_2
X_14208_ _14763_/S _14206_/Y _14207_/X _14129_/Y vssd1 vssd1 vccd1 vccd1 _17594_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_99_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15188_ _15188_/A _15188_/B vssd1 vssd1 vccd1 vccd1 _15188_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14139_ _14221_/A _14139_/B vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__or2_1
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout409 _14775_/A vssd1 vssd1 vccd1 vccd1 _13950_/A sky130_fd_sc_hd__buf_6
XFILLER_99_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09680_ _09678_/B _09675_/C _09675_/B vssd1 vssd1 vccd1 vccd1 _09681_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09114_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09114_/Y sky130_fd_sc_hd__nor3_4
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09045_ _17387_/A _12795_/B _09044_/B _09041_/Y vssd1 vssd1 vccd1 vccd1 _09047_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xmax_cap193 _15209_/Y vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__buf_6
XFILLER_81_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout910 _17290_/A2 vssd1 vssd1 vccd1 vccd1 _17293_/A2 sky130_fd_sc_hd__buf_4
Xfanout921 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17426_/C1 sky130_fd_sc_hd__buf_4
XFILLER_132_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09947_ _10560_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout932 fanout933/X vssd1 vssd1 vccd1 vccd1 fanout932/X sky130_fd_sc_hd__clkbuf_4
Xfanout943 fanout944/X vssd1 vssd1 vccd1 vccd1 fanout943/X sky130_fd_sc_hd__buf_2
XTAP_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__xnor2_2
XTAP_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08829_ _08828_/B _08829_/B vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__nand2b_2
XFILLER_86_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11840_ _14912_/B _11840_/B vssd1 vssd1 vccd1 vccd1 _11840_/Y sky130_fd_sc_hd__nand2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11771_/A _11771_/B vssd1 vssd1 vccd1 vccd1 _11771_/Y sky130_fd_sc_hd__nand2_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _13267_/X _13511_/B _13509_/Y _13385_/B vssd1 vssd1 vccd1 vccd1 _13510_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ _10722_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__xnor2_4
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14490_ _14557_/B _14490_/B vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__nor2_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ _13441_/A vssd1 vssd1 vccd1 vccd1 _13600_/A sky130_fd_sc_hd__inv_2
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10653_ _10653_/A _10653_/B _10653_/C vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__nand3_2
XFILLER_186_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16160_ _16161_/A _16161_/B vssd1 vssd1 vccd1 vccd1 _16160_/X sky130_fd_sc_hd__or2_1
XFILLER_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13372_ _13496_/A _13370_/Y _13240_/Y _13244_/B vssd1 vssd1 vccd1 vccd1 _13373_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_166_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10584_ _10579_/A _10577_/X _10325_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10584_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15111_ _11469_/X _15804_/A2 _15713_/B1 _15116_/B vssd1 vssd1 vccd1 vccd1 _15111_/X
+ sky130_fd_sc_hd__a22o_1
X_12323_ _12323_/A _12492_/A _12323_/C vssd1 vssd1 vccd1 vccd1 _12492_/B sky130_fd_sc_hd__nor3_2
X_16091_ _16092_/A _16092_/B vssd1 vssd1 vccd1 vccd1 _16200_/A sky130_fd_sc_hd__nand2b_2
XFILLER_5_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15042_ _15130_/S _15401_/A _15796_/B vssd1 vssd1 vccd1 vccd1 _15042_/X sky130_fd_sc_hd__or3_4
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12254_ _12078_/A _12080_/B _12078_/B vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__o21ba_4
XFILLER_141_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ _11739_/A _11205_/B vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__nand2_4
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _11988_/A _11988_/B _11987_/A vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__a21oi_4
X_11136_ _11137_/B _11137_/C _11137_/A vssd1 vssd1 vccd1 vccd1 _11293_/A sky130_fd_sc_hd__o21ai_2
XFILLER_150_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16993_ _17046_/B _16993_/B vssd1 vssd1 vccd1 vccd1 _16996_/B sky130_fd_sc_hd__and2b_1
XFILLER_77_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15944_ _15944_/A _15944_/B vssd1 vssd1 vccd1 vccd1 _15972_/A sky130_fd_sc_hd__xnor2_2
X_11067_ _11069_/B vssd1 vssd1 vccd1 vccd1 _11067_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10018_ _10018_/A _10018_/B _10019_/B vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__or3_1
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15875_ _15875_/A _15875_/B vssd1 vssd1 vccd1 vccd1 _15875_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17614_ fanout946/X _17614_/D vssd1 vssd1 vccd1 vccd1 _17614_/Q sky130_fd_sc_hd__dfxtp_4
X_14826_ _17023_/A _14825_/Y _14764_/Y _14434_/Y vssd1 vssd1 vccd1 vccd1 _14826_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_52_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ fanout946/X _17545_/D vssd1 vssd1 vccd1 vccd1 _17545_/Q sky130_fd_sc_hd__dfxtp_4
X_14757_ _13832_/B _13834_/A _14840_/A vssd1 vssd1 vccd1 vccd1 _14758_/B sky130_fd_sc_hd__mux2_1
X_11969_ _11970_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__or2_4
X_13708_ _13594_/X _13598_/A _13706_/Y _13707_/X vssd1 vssd1 vccd1 vccd1 _13817_/A
+ sky130_fd_sc_hd__o211a_4
X_17476_ fanout929/X _17476_/D vssd1 vssd1 vccd1 vccd1 _17476_/Q sky130_fd_sc_hd__dfxtp_4
X_14688_ _14688_/A _14688_/B vssd1 vssd1 vccd1 vccd1 _14689_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13639_ _13638_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13645_/B sky130_fd_sc_hd__a21o_1
X_16427_ _16333_/X _16337_/B _16335_/B vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__o21ai_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16358_ _16358_/A _16358_/B _16358_/C vssd1 vssd1 vccd1 vccd1 _16359_/B sky130_fd_sc_hd__or3_1
XFILLER_118_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15309_ _15309_/A _15309_/B _15307_/X vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__or3b_1
XFILLER_121_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16289_ _16290_/A _16290_/B _16290_/C vssd1 vssd1 vccd1 vccd1 _16382_/B sky130_fd_sc_hd__o21a_1
XFILLER_173_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout206 _16583_/A1 vssd1 vssd1 vccd1 vccd1 _16735_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_141_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09801_ _09801_/A _09801_/B _09941_/A vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__nor3_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout228 _16008_/B1 vssd1 vssd1 vccd1 vccd1 _15713_/B1 sky130_fd_sc_hd__buf_4
Xfanout239 _16218_/C1 vssd1 vssd1 vccd1 vccd1 _16008_/C1 sky130_fd_sc_hd__buf_6
XFILLER_80_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09732_ _09733_/B _09733_/A vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__and2b_2
XFILLER_189_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _09499_/Y _09500_/X _09789_/A _09774_/B _09774_/A vssd1 vssd1 vccd1 vccd1
+ _09665_/B sky130_fd_sc_hd__a32o_1
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09594_ _09588_/X _09723_/A _09580_/X _09581_/Y vssd1 vssd1 vccd1 vccd1 _09597_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09028_ _12245_/A _12637_/C vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__nand2_8
XFILLER_151_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout740 _17494_/Q vssd1 vssd1 vccd1 vccd1 _13229_/B sky130_fd_sc_hd__buf_8
XFILLER_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout751 _09428_/B vssd1 vssd1 vccd1 vccd1 _10899_/D sky130_fd_sc_hd__buf_6
XFILLER_172_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout762 _10897_/B vssd1 vssd1 vccd1 vccd1 _10791_/C sky130_fd_sc_hd__buf_12
X_13990_ _13990_/A _13990_/B vssd1 vssd1 vccd1 vccd1 _14011_/A sky130_fd_sc_hd__xor2_4
Xfanout773 _13196_/B vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__buf_12
Xfanout784 _10640_/D vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__buf_6
Xfanout795 _10738_/D vssd1 vssd1 vccd1 vccd1 _10933_/D sky130_fd_sc_hd__buf_6
XFILLER_65_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12941_ _17411_/A _13229_/B _13100_/B _17413_/A vssd1 vssd1 vccd1 vccd1 _12945_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15660_ _15660_/A _15661_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _15660_/X sky130_fd_sc_hd__and3_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12872_/A _12872_/B vssd1 vssd1 vccd1 vccd1 _12875_/A sky130_fd_sc_hd__xnor2_4
XFILLER_2_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14612_/A _14612_/B vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__and2b_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11823_ _17304_/A1 _17302_/A1 _12060_/S vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__mux2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/A _15591_/B vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__or2_4
XFILLER_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _13764_/D _17360_/A2 _17329_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17494_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _15457_/B _13015_/B _14210_/B _13012_/X vssd1 vssd1 vccd1 vccd1 _14543_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11754_ _11753_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11755_/B sky130_fd_sc_hd__a21o_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _17596_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17261_/X sky130_fd_sc_hd__a21o_1
X_10705_ _10705_/A _10705_/B vssd1 vssd1 vccd1 vccd1 _11030_/B sky130_fd_sc_hd__nor2_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14473_/A _14473_/B _14473_/C vssd1 vssd1 vccd1 vccd1 _14533_/B sky130_fd_sc_hd__nand3_2
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11685_ _15235_/A _15235_/B vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16212_ _16107_/Y _16111_/B _16210_/Y vssd1 vssd1 vccd1 vccd1 _16212_/Y sky130_fd_sc_hd__o21ai_1
X_13424_ _13308_/A _13309_/B _13421_/Y _13422_/X vssd1 vssd1 vccd1 vccd1 _13428_/A
+ sky130_fd_sc_hd__a211oi_4
X_17192_ input18/X input17/X input19/X input23/X vssd1 vssd1 vccd1 vccd1 _17195_/A
+ sky130_fd_sc_hd__or4b_1
X_10636_ _10550_/X _10634_/Y _10632_/B _10614_/X vssd1 vssd1 vccd1 vccd1 _10636_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16143_ _16241_/B _16143_/B vssd1 vssd1 vccd1 vccd1 _16146_/A sky130_fd_sc_hd__nor2_4
XFILLER_155_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13355_ _13355_/A _13355_/B vssd1 vssd1 vccd1 vccd1 _13357_/B sky130_fd_sc_hd__xnor2_2
XFILLER_154_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__or2_2
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12306_ _12306_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__nor2_4
X_16074_ _16075_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _16188_/B sky130_fd_sc_hd__and2b_1
XFILLER_154_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13286_ _13745_/B _14002_/B _13523_/B _13852_/A vssd1 vssd1 vccd1 vccd1 _13286_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10499_/A sky130_fd_sc_hd__or2_2
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15025_ _15305_/C _15025_/B vssd1 vssd1 vccd1 vccd1 _15025_/Y sky130_fd_sc_hd__nor2_2
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _12237_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12238_/B sky130_fd_sc_hd__nand2_2
XFILLER_151_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12168_ _12169_/A _12169_/B _12169_/C vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__a21oi_1
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11119_ _11124_/C _10971_/B _10878_/A _10876_/Y vssd1 vssd1 vccd1 vccd1 _11121_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12099_ _11891_/A _11891_/Y _12097_/X _12268_/B vssd1 vssd1 vccd1 vccd1 _12122_/A
+ sky130_fd_sc_hd__o211ai_4
X_16976_ _16653_/A _14590_/B _16582_/A _15628_/B vssd1 vssd1 vccd1 vccd1 _16977_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15927_ _15925_/Y _15927_/B vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__and2b_2
Xinput6 i_wb_addr[12] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15858_ _15858_/A _15858_/B vssd1 vssd1 vccd1 vccd1 _15859_/B sky130_fd_sc_hd__xnor2_4
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14809_ _15707_/B _15707_/C _10145_/B vssd1 vssd1 vccd1 vccd1 _15802_/A sky130_fd_sc_hd__a21o_1
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15789_ _15610_/A _15698_/A _15698_/B vssd1 vssd1 vccd1 vccd1 _15789_/X sky130_fd_sc_hd__o21ba_1
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17528_ fanout930/X _17528_/D vssd1 vssd1 vccd1 vccd1 _17528_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17459_ fanout941/X _17459_/D vssd1 vssd1 vccd1 vccd1 _17459_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09715_ _09711_/X _09713_/X _16982_/B _09710_/Y vssd1 vssd1 vccd1 vccd1 _09717_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _09969_/A _09646_/B vssd1 vssd1 vccd1 vccd1 _09647_/C sky130_fd_sc_hd__nor2_1
XFILLER_83_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A _09577_/B _09596_/B vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__and3_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11470_ _14791_/A _11629_/C vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10421_ _10422_/A _10420_/Y _10647_/C _10755_/D vssd1 vssd1 vccd1 vccd1 _10531_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13140_ _13268_/B _13140_/B vssd1 vssd1 vccd1 vccd1 _13140_/Y sky130_fd_sc_hd__nand2_1
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10465_/A sky130_fd_sc_hd__xor2_2
XFILLER_174_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13071_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13244_/A sky130_fd_sc_hd__o21a_2
X_10283_ _10283_/A _10283_/B _10283_/C _10283_/D vssd1 vssd1 vccd1 vccd1 _10283_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_982 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12022_ _10180_/C _14952_/B _12053_/A vssd1 vssd1 vccd1 vccd1 _12022_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16830_ _16830_/A _16830_/B vssd1 vssd1 vccd1 vccd1 _16832_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout570 _11268_/A vssd1 vssd1 vccd1 vccd1 _11553_/B sky130_fd_sc_hd__buf_6
Xfanout581 _14792_/A vssd1 vssd1 vccd1 vccd1 _14922_/S sky130_fd_sc_hd__buf_4
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout592 _12214_/A vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13973_ _13864_/B _13870_/B _13862_/X vssd1 vssd1 vccd1 vccd1 _13974_/B sky130_fd_sc_hd__a21oi_4
X_16761_ _16761_/A _16761_/B vssd1 vssd1 vccd1 vccd1 _16762_/B sky130_fd_sc_hd__xnor2_2
XFILLER_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15712_ _16011_/A _15103_/X _15711_/Y _17164_/C vssd1 vssd1 vccd1 vccd1 _15712_/X
+ sky130_fd_sc_hd__a211o_1
X_12924_ _12924_/A _12924_/B vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__nor2_1
XFILLER_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16692_ _16693_/B _16692_/B vssd1 vssd1 vccd1 vccd1 _16777_/A sky130_fd_sc_hd__nand2b_2
XFILLER_47_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15643_ _15732_/A _15643_/B vssd1 vssd1 vccd1 vccd1 _15742_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _12847_/A _12852_/X _12854_/Y _12850_/X vssd1 vssd1 vccd1 vccd1 _12856_/B
+ sky130_fd_sc_hd__o31a_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _17363_/A _09928_/D _09926_/C vssd1 vssd1 vccd1 vccd1 _11807_/B sky130_fd_sc_hd__a21o_1
X_15574_ _16935_/A _15071_/A _17038_/C vssd1 vssd1 vccd1 vccd1 _15658_/B sky130_fd_sc_hd__a21oi_4
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _14770_/A _13100_/B _13551_/D _14769_/A vssd1 vssd1 vccd1 vccd1 _12790_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14526_/B sky130_fd_sc_hd__o21ai_1
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ input66/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17313_/X sky130_fd_sc_hd__or3_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11739_/B vssd1 vssd1 vccd1 vccd1 _11737_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14456_ _14456_/A _14456_/B _14456_/C vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__nand3_1
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17244_ _17558_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__and2_1
X_11668_ _11646_/A _11646_/B _11646_/C vssd1 vssd1 vccd1 vccd1 _11670_/C sky130_fd_sc_hd__a21o_1
XFILLER_168_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13407_ _13643_/A _13948_/D vssd1 vssd1 vccd1 vccd1 _13408_/B sky130_fd_sc_hd__nand2_2
X_10619_ _10962_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10716_/A sky130_fd_sc_hd__nand2_8
X_17175_ input15/X input18/X input17/X input20/X vssd1 vssd1 vccd1 vccd1 _17181_/C
+ sky130_fd_sc_hd__or4_1
X_14387_ _14387_/A _14554_/B vssd1 vssd1 vccd1 vccd1 _14388_/B sky130_fd_sc_hd__nand2_2
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11599_ _11555_/A _11555_/B _11637_/A vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__o21bai_1
X_16126_ _16315_/B _16681_/D _16409_/B _16025_/A vssd1 vssd1 vccd1 vccd1 _16126_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13338_ _13338_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13339_/C sky130_fd_sc_hd__nor2_1
XFILLER_182_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16057_ _16055_/A _15658_/Y _16827_/D _15081_/A vssd1 vssd1 vccd1 vccd1 _16058_/B
+ sky130_fd_sc_hd__o22a_1
X_13269_ _13010_/B _13511_/A _13267_/X vssd1 vssd1 vccd1 vccd1 _13271_/B sky130_fd_sc_hd__a21oi_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _15008_/A _15008_/B vssd1 vssd1 vccd1 vccd1 _15008_/X sky130_fd_sc_hd__or2_1
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16959_ _17008_/A _17012_/A vssd1 vssd1 vccd1 vccd1 _16960_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09500_ _09620_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09500_/X sky130_fd_sc_hd__or2_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _10255_/A _09428_/B _09430_/B _09427_/Y vssd1 vssd1 vccd1 vccd1 _09433_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09362_ _09497_/A _09361_/Y _12176_/A _09944_/D vssd1 vssd1 vccd1 vccd1 _09504_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_40_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__nor2_1
XANTENNA_11 _17609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _17447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1027 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_33 _17429_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 _15373_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_55 _17306_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_66 _17497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_77 _17542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_88 _14829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10970_ _10970_/A _10970_/B vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__nand2_4
XFILLER_44_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__nand2_2
XFILLER_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12640_ _12640_/A _12792_/A _12640_/C vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__nor3_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12571_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__o21ai_2
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14310_ _14230_/B _14232_/B _14230_/A vssd1 vssd1 vccd1 vccd1 _14312_/B sky130_fd_sc_hd__o21ba_1
XFILLER_15_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11522_ _11522_/A _11522_/B _11523_/B vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__or3_1
XFILLER_169_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15290_ _15774_/A _16136_/B _15291_/A vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__and3_1
XFILLER_183_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14241_ _14450_/A _14318_/B _14641_/D _14545_/C vssd1 vssd1 vccd1 vccd1 _14242_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11453_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__nand2_1
XFILLER_183_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ _10262_/X _10357_/Y _10385_/A _10385_/Y vssd1 vssd1 vccd1 vccd1 _10405_/D
+ sky130_fd_sc_hd__o211a_2
X_14172_ _14173_/A _14173_/B _14173_/C vssd1 vssd1 vccd1 vccd1 _14252_/A sky130_fd_sc_hd__o21ai_4
XFILLER_152_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11384_ _11395_/B _11435_/A _11395_/A vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_178_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ _13123_/A _13123_/B vssd1 vssd1 vccd1 vccd1 _13125_/C sky130_fd_sc_hd__or2_2
X_10335_ _10193_/B _10229_/X _10319_/A _10319_/Y vssd1 vssd1 vccd1 vccd1 _10336_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13054_ _13055_/A _13055_/B vssd1 vssd1 vccd1 vccd1 _13186_/A sky130_fd_sc_hd__or2_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10266_ _10267_/A _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__a21o_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12005_ _12005_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12007_/B sky130_fd_sc_hd__nand2_2
XFILLER_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ _10198_/A _10198_/C vssd1 vssd1 vccd1 vccd1 _10322_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16813_ _16938_/B _16813_/B vssd1 vssd1 vccd1 vccd1 _16813_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16744_ _16744_/A _16744_/B vssd1 vssd1 vccd1 vccd1 _16746_/A sky130_fd_sc_hd__nor2_2
X_13956_ _13958_/A _13958_/B vssd1 vssd1 vccd1 vccd1 _14130_/A sky130_fd_sc_hd__nor2_1
XFILLER_185_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ _12907_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _12908_/B sky130_fd_sc_hd__nand2_2
X_13887_ _13888_/A _13888_/B vssd1 vssd1 vccd1 vccd1 _13990_/A sky130_fd_sc_hd__nor2_4
X_16675_ _16503_/Y _16670_/B _16597_/B _16597_/A vssd1 vssd1 vccd1 vccd1 _16676_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_185_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12838_ _13001_/B _12837_/Y _12689_/A _12691_/A vssd1 vssd1 vccd1 vccd1 _12838_/Y
+ sky130_fd_sc_hd__a211oi_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15626_ _15622_/B _15899_/A2 _15625_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15626_/Y
+ sky130_fd_sc_hd__a211oi_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15557_ _15557_/A _15557_/B vssd1 vssd1 vccd1 vccd1 _15559_/B sky130_fd_sc_hd__xnor2_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12770_/B _12923_/D _12770_/D _12770_/A vssd1 vssd1 vccd1 vccd1 _12771_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14508_ _14508_/A _14508_/B vssd1 vssd1 vccd1 vccd1 _14514_/A sky130_fd_sc_hd__xnor2_1
XFILLER_159_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15488_ _15489_/A _15489_/B vssd1 vssd1 vccd1 vccd1 _15488_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 i_wb_addr[25] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_2
X_17227_ _17443_/Q _17233_/A2 _17225_/X _17226_/X _17372_/C1 vssd1 vssd1 vccd1 vccd1
+ _17443_/D sky130_fd_sc_hd__o221a_1
X_14439_ _14440_/A _14440_/B _14440_/C vssd1 vssd1 vccd1 vccd1 _14441_/A sky130_fd_sc_hd__o21a_1
Xinput31 i_wb_addr[6] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
Xinput42 i_wb_data[15] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 i_wb_data[25] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
Xinput64 i_wb_data[6] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17158_ _11778_/Y _17157_/Y _17070_/B vssd1 vssd1 vccd1 vccd1 _17158_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_116_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _16001_/A _16003_/X _16107_/Y _16108_/X vssd1 vssd1 vccd1 vccd1 _16111_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_171_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17089_ _17089_/A _17089_/B vssd1 vssd1 vccd1 vccd1 _17118_/A sky130_fd_sc_hd__nor2_2
X_09980_ _10236_/B _10479_/B _17468_/D _10236_/A vssd1 vssd1 vccd1 vccd1 _09980_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_115_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08931_ _08929_/A _08929_/Y _08872_/X _08874_/X vssd1 vssd1 vccd1 vccd1 _09016_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_103_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08862_ _08862_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08793_ _12258_/A _12088_/D _08790_/Y _11878_/A vssd1 vssd1 vccd1 vccd1 _08794_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ _12243_/A _12243_/B _09414_/C _09555_/C vssd1 vssd1 vccd1 vccd1 _09415_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_164_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09345_ _09358_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__nor2_1
XFILLER_178_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09276_ _09404_/A _09404_/B vssd1 vssd1 vccd1 vccd1 _09290_/C sky130_fd_sc_hd__nand2_1
XFILLER_193_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10133_/C sky130_fd_sc_hd__nand2_2
XFILLER_164_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10051_ _09930_/A _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__o21ai_1
XFILLER_76_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13810_ _13923_/A _13810_/B vssd1 vssd1 vccd1 vccd1 _13812_/B sky130_fd_sc_hd__or2_2
X_14790_ _14790_/A _14848_/B vssd1 vssd1 vccd1 vccd1 _14790_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13741_ _13741_/A _13741_/B _13741_/C vssd1 vssd1 vccd1 vccd1 _13742_/B sky130_fd_sc_hd__nor3_2
X_10953_ _10953_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _11069_/A sky130_fd_sc_hd__xnor2_4
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16460_ _16550_/B _16460_/B vssd1 vssd1 vccd1 vccd1 _16460_/Y sky130_fd_sc_hd__nand2_1
X_13672_ _13558_/A _13559_/Y _13670_/Y _13770_/B vssd1 vssd1 vccd1 vccd1 _13814_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10884_ _10884_/A _10884_/B vssd1 vssd1 vccd1 vccd1 _10891_/A sky130_fd_sc_hd__xnor2_2
X_15411_ _15140_/Y _15206_/B _15450_/A vssd1 vssd1 vccd1 vccd1 _15956_/B sky130_fd_sc_hd__o21ai_4
X_12623_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__or2_1
X_16391_ _16399_/A _16391_/B vssd1 vssd1 vccd1 vccd1 _16391_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15342_ _15342_/A _15661_/A vssd1 vssd1 vccd1 vccd1 _15342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12554_ _11849_/A _12550_/X _12553_/X _17165_/A1 vssd1 vssd1 vccd1 vccd1 _12555_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1066 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11487_/A _11487_/B _11485_/X vssd1 vssd1 vccd1 vccd1 _11527_/B sky130_fd_sc_hd__o21ba_2
XFILLER_185_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15273_ _15948_/A _15752_/A vssd1 vssd1 vccd1 vccd1 _15578_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12485_ _12311_/A _12311_/B _12310_/A vssd1 vssd1 vccd1 vccd1 _12519_/A sky130_fd_sc_hd__a21oi_4
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14224_ _14680_/A _14599_/B _14485_/D _14360_/C vssd1 vssd1 vccd1 vccd1 _14225_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_184_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17012_ _17012_/A _17012_/B vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11436_ _11436_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__xnor2_4
XFILLER_125_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14155_ _14226_/A _14155_/B vssd1 vssd1 vccd1 vccd1 _14156_/B sky130_fd_sc_hd__nand2_2
XFILLER_153_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11367_ _11367_/A _11448_/A _11367_/C vssd1 vssd1 vccd1 vccd1 _11403_/A sky130_fd_sc_hd__or3_4
XFILLER_99_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__xor2_1
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _10157_/Y _10230_/X _10263_/X _10283_/X vssd1 vssd1 vccd1 vccd1 _10319_/D
+ sky130_fd_sc_hd__a211o_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14086_ _14087_/B _14086_/B vssd1 vssd1 vccd1 vccd1 _14088_/A sky130_fd_sc_hd__nand2b_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11153_/C _11235_/X _11290_/Y _11296_/Y vssd1 vssd1 vccd1 vccd1 _11299_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _17387_/A _13300_/D vssd1 vssd1 vccd1 vccd1 _13038_/B sky130_fd_sc_hd__nand2_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _10262_/A vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14988_ _15100_/A _14988_/B vssd1 vssd1 vccd1 vccd1 _14988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16727_ _16728_/B _16727_/B vssd1 vssd1 vccd1 vccd1 _16794_/B sky130_fd_sc_hd__nand2b_2
X_13939_ _13939_/A vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16658_ _15794_/A _16641_/Y _16648_/X _16657_/X vssd1 vssd1 vccd1 vccd1 _16658_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_179_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15609_ _15609_/A _15609_/B _15609_/C vssd1 vssd1 vccd1 vccd1 _15610_/B sky130_fd_sc_hd__nor3_2
X_16589_ _16812_/A _16589_/B _16743_/C _17043_/B vssd1 vssd1 vccd1 vccd1 _16686_/A
+ sky130_fd_sc_hd__and4_2
X_09130_ _09139_/B _09130_/B vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__nor2_4
XFILLER_188_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_944 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09061_ _09061_/A _09298_/A vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09963_ _09923_/A _09957_/A _09964_/A _09962_/X vssd1 vssd1 vccd1 vccd1 _10091_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08914_ _12107_/B _13094_/B _13088_/B _12275_/A vssd1 vssd1 vccd1 vccd1 _08914_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_58_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09895_/A _09893_/Y _10970_/A _10659_/D vssd1 vssd1 vccd1 vccd1 _10021_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_100_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08845_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__xnor2_1
XFILLER_44_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _09030_/A _12638_/B _08776_/C vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__and3_2
XFILLER_100_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09328_ _09328_/A _09451_/A _09328_/C vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__or3_1
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09259_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09338_/A sky130_fd_sc_hd__or2_2
XFILLER_182_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ _17379_/A _12270_/B _12270_/C _12270_/D vssd1 vssd1 vccd1 vccd1 _12271_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__xor2_4
XFILLER_134_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _11153_/B _11153_/C _11153_/A vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__o21a_4
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10103_ _10057_/A _10057_/C _10057_/B vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__a21oi_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15960_ _15960_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15963_/A sky130_fd_sc_hd__xnor2_4
X_11083_ _11064_/X _11071_/Y _11080_/B _11145_/A vssd1 vssd1 vccd1 vccd1 _11084_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10034_ _10034_/A _10042_/A _10034_/C vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__or3_1
X_14911_ _14788_/A _14911_/B vssd1 vssd1 vccd1 vccd1 _15059_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15891_ _15898_/A _15891_/B _16809_/A vssd1 vssd1 vccd1 vccd1 _15891_/X sky130_fd_sc_hd__or3b_2
XFILLER_76_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14842_ _14667_/A _14839_/Y _14840_/Y _14841_/Y _11848_/Y vssd1 vssd1 vccd1 vccd1
+ _14842_/X sky130_fd_sc_hd__o32a_1
XFILLER_124_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17561_ fanout938/X _17561_/D vssd1 vssd1 vccd1 vccd1 _17561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _11986_/B _11985_/B vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__and2b_2
X_14773_ _16644_/C _16651_/A vssd1 vssd1 vccd1 vccd1 _16649_/B sky130_fd_sc_hd__or2_2
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16512_ _16604_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16514_/C sky130_fd_sc_hd__nand2_1
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13724_ _13614_/A _13614_/B _13612_/A vssd1 vssd1 vccd1 vccd1 _13726_/B sky130_fd_sc_hd__a21oi_1
X_10936_ _10936_/A _10936_/B vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__xnor2_4
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17492_ fanout930/X _17492_/D vssd1 vssd1 vccd1 vccd1 _17492_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_182_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16443_ _16443_/A _16443_/B vssd1 vssd1 vccd1 vccd1 _16457_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13655_ _13654_/B _13655_/B vssd1 vssd1 vccd1 vccd1 _13656_/B sky130_fd_sc_hd__nand2b_1
X_10867_ _14788_/A _14906_/A vssd1 vssd1 vccd1 vccd1 _14801_/A sky130_fd_sc_hd__and2_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12606_ _12607_/A _12607_/B _12607_/C vssd1 vssd1 vccd1 vccd1 _12778_/A sky130_fd_sc_hd__o21ai_2
X_16374_ _16375_/B _16375_/A vssd1 vssd1 vccd1 vccd1 _16470_/A sky130_fd_sc_hd__nand2b_1
X_13586_ _13586_/A _13586_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__nor3_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10798_ _14787_/A _15381_/A vssd1 vssd1 vccd1 vccd1 _10800_/C sky130_fd_sc_hd__and2_4
XFILLER_185_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15325_ _15069_/A _17613_/Q _15071_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15325_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_129_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12537_ _12366_/A _12366_/B _12368_/B _12370_/A _12370_/B vssd1 vssd1 vccd1 vccd1
+ _12540_/B sky130_fd_sc_hd__o32ai_4
XFILLER_118_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12662_/B _12468_/B vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__nor2_4
X_15256_ _14356_/S _16735_/A _12553_/B _15808_/A _15255_/X vssd1 vssd1 vccd1 vccd1
+ _15256_/X sky130_fd_sc_hd__o32a_1
XFILLER_32_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14207_ _14278_/B _14207_/B vssd1 vssd1 vccd1 vccd1 _14207_/X sky130_fd_sc_hd__or2_1
X_11419_ _11419_/A _11419_/B vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__xnor2_4
X_15187_ _11321_/X _15804_/A2 _15184_/X _15186_/X _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15188_/B sky130_fd_sc_hd__a2111o_1
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12399_ _13837_/C _12398_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _12400_/B sky130_fd_sc_hd__mux2_1
XFILLER_67_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14138_ _14138_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14139_/B sky130_fd_sc_hd__and2_1
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14069_ _13978_/A _13980_/B _13978_/B vssd1 vssd1 vccd1 vccd1 _14071_/B sky130_fd_sc_hd__o21ba_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09113_ _09115_/A _09115_/B _09115_/C vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__o21ai_4
XFILLER_149_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ _09041_/Y _09044_/B vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__and2b_2
XFILLER_164_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout900 _10559_/B vssd1 vssd1 vccd1 vccd1 _11553_/D sky130_fd_sc_hd__buf_2
Xfanout911 _17266_/A2 vssd1 vssd1 vccd1 vccd1 _17290_/A2 sky130_fd_sc_hd__buf_6
Xfanout922 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17293_/C1 sky130_fd_sc_hd__buf_4
XFILLER_104_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09946_ _09948_/B _09948_/A vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__and2b_1
Xfanout933 fanout937/X vssd1 vssd1 vccd1 vccd1 fanout933/X sky130_fd_sc_hd__clkbuf_4
Xfanout944 input2/X vssd1 vssd1 vccd1 vccd1 fanout944/X sky130_fd_sc_hd__buf_6
XTAP_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09878_/B _09878_/A vssd1 vssd1 vccd1 vccd1 _09877_/X sky130_fd_sc_hd__and2b_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08829_/B _08828_/B vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__nand2b_1
XFILLER_100_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _12243_/B _11859_/C vssd1 vssd1 vccd1 vccd1 _08776_/C sky130_fd_sc_hd__and2_4
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _10583_/A _11771_/B _11771_/A vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_26_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10722_/B _10722_/A vssd1 vssd1 vccd1 vccd1 _10721_/X sky130_fd_sc_hd__and2b_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _13442_/A _13442_/B vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__and2b_1
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10652_ _10653_/B _10653_/C _10653_/A vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__a21o_1
XFILLER_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _13240_/Y _13244_/B _13496_/A _13370_/Y vssd1 vssd1 vccd1 vccd1 _13496_/B
+ sky130_fd_sc_hd__a211oi_4
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _16972_/A sky130_fd_sc_hd__and2_4
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12322_ _12323_/A _12492_/A _12323_/C vssd1 vssd1 vccd1 vccd1 _12324_/A sky130_fd_sc_hd__o21a_1
X_15110_ _15116_/B _15110_/B vssd1 vssd1 vccd1 vccd1 _15110_/Y sky130_fd_sc_hd__nor2_1
X_16090_ _15984_/A _15984_/B _15975_/Y vssd1 vssd1 vccd1 vccd1 _16092_/B sky130_fd_sc_hd__a21bo_4
XFILLER_155_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15041_ _14792_/A _15373_/B _15274_/A vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _12089_/A _12091_/B _12089_/B vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__o21ba_4
XFILLER_5_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11205_/B sky130_fd_sc_hd__nand2_1
X_12184_ _12351_/A _12351_/B vssd1 vssd1 vccd1 vccd1 _12186_/A sky130_fd_sc_hd__xnor2_4
X_11135_ _11520_/C _11135_/B _11135_/C vssd1 vssd1 vccd1 vccd1 _11137_/C sky130_fd_sc_hd__and3_1
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16992_ _16991_/A _16991_/C _16991_/D _16991_/B vssd1 vssd1 vccd1 vccd1 _16993_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_110_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15943_ _15944_/A _15944_/B vssd1 vssd1 vccd1 vccd1 _16080_/A sky130_fd_sc_hd__nor2_2
X_11066_ _11065_/B _11065_/Y _11055_/X _11056_/Y vssd1 vssd1 vccd1 vccd1 _11069_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10017_ _10017_/A _10140_/A vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__nor2_4
XFILLER_37_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15874_ _15989_/B _15874_/B vssd1 vssd1 vccd1 vccd1 _15875_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17613_ fanout946/X _17613_/D vssd1 vssd1 vccd1 vccd1 _17613_/Q sky130_fd_sc_hd__dfxtp_2
X_14825_ _17023_/B _17024_/A vssd1 vssd1 vccd1 vccd1 _14825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ fanout929/X _17544_/D vssd1 vssd1 vccd1 vccd1 _17544_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756_ _14756_/A1 _14754_/Y _14755_/X _14734_/Y _14735_/X vssd1 vssd1 vccd1 vccd1
+ _17605_/D sky130_fd_sc_hd__a32o_1
X_11968_ _12800_/A _12166_/B vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _13707_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13707_/X sky130_fd_sc_hd__or2_2
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17475_ fanout928/X _17608_/Q vssd1 vssd1 vccd1 vccd1 _17475_/Q sky130_fd_sc_hd__dfxtp_4
X_10919_ _14788_/A _15541_/A vssd1 vssd1 vccd1 vccd1 _10924_/A sky130_fd_sc_hd__nand2_2
X_14687_ _14688_/A _14688_/B vssd1 vssd1 vccd1 vccd1 _14717_/A sky130_fd_sc_hd__or2_1
X_11899_ _11900_/B _12258_/B _12090_/B _12107_/A vssd1 vssd1 vccd1 vccd1 _11901_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16426_ _16527_/A _16426_/B vssd1 vssd1 vccd1 vccd1 _16439_/A sky130_fd_sc_hd__nand2b_2
X_13638_ _13638_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__nand3_2
XFILLER_160_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16357_ _16358_/A _16358_/B _16358_/C vssd1 vssd1 vccd1 vccd1 _16443_/A sky130_fd_sc_hd__o21ai_1
XFILLER_146_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13569_ _13569_/A _13569_/B _13569_/C vssd1 vssd1 vccd1 vccd1 _13571_/A sky130_fd_sc_hd__or3_1
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15308_ _15307_/A _15307_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _15309_/A sky130_fd_sc_hd__o21a_1
X_16288_ _16288_/A _16288_/B vssd1 vssd1 vccd1 vccd1 _16290_/C sky130_fd_sc_hd__xnor2_1
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15239_ _15175_/X _15176_/Y _15174_/Y vssd1 vssd1 vccd1 vccd1 _15241_/C sky130_fd_sc_hd__a21bo_1
XFILLER_161_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09800_ _09801_/B _09941_/A _09801_/A vssd1 vssd1 vccd1 vccd1 _09805_/B sky130_fd_sc_hd__o21a_2
Xfanout207 _11849_/Y vssd1 vssd1 vccd1 vccd1 _16583_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout218 _16745_/B vssd1 vssd1 vccd1 vccd1 _16935_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout229 _14933_/Y vssd1 vssd1 vccd1 vccd1 _16008_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_101_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09731_ _09731_/A _09872_/A vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09662_ _09662_/A _09662_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__nor2_4
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09593_ _09580_/X _09581_/Y _09588_/X _09723_/A vssd1 vssd1 vccd1 vccd1 _09597_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1071 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09027_ _09027_/A _09027_/B _09033_/B vssd1 vssd1 vccd1 vccd1 _09048_/B sky130_fd_sc_hd__or3_2
XFILLER_163_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout730 _09892_/C vssd1 vssd1 vccd1 vccd1 _10755_/D sky130_fd_sc_hd__clkbuf_8
Xfanout741 _10993_/D vssd1 vssd1 vccd1 vccd1 _09892_/D sky130_fd_sc_hd__buf_8
X_09929_ _09929_/A _10184_/A vssd1 vssd1 vccd1 vccd1 _09930_/C sky130_fd_sc_hd__nor2_1
Xfanout752 fanout757/X vssd1 vssd1 vccd1 vccd1 _09428_/B sky130_fd_sc_hd__buf_8
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout763 _17492_/Q vssd1 vssd1 vccd1 vccd1 _10897_/B sky130_fd_sc_hd__buf_6
XFILLER_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout774 _13196_/B vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__clkbuf_4
Xfanout785 _10791_/D vssd1 vssd1 vccd1 vccd1 _10640_/D sky130_fd_sc_hd__buf_8
Xfanout796 _11135_/B vssd1 vssd1 vccd1 vccd1 _10738_/D sky130_fd_sc_hd__buf_8
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _12780_/A _12779_/B _12779_/A vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__o21ba_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _17401_/A _13564_/C vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__nand2_2
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14610_ _14683_/A _14610_/B vssd1 vssd1 vccd1 vccd1 _14612_/B sky130_fd_sc_hd__nor2_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11820_/Y _11821_/X _15538_/A vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__mux2_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15590_/A _15590_/B _15590_/C vssd1 vssd1 vccd1 vccd1 _15591_/B sky130_fd_sc_hd__and3_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11753_ _11753_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11759_/A sky130_fd_sc_hd__and3_4
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14421_/S _14637_/A1 _11820_/A _08718_/A vssd1 vssd1 vccd1 vccd1 _14541_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _10905_/B _11005_/B _10805_/D _10905_/A vssd1 vssd1 vccd1 vccd1 _10705_/B
+ sky130_fd_sc_hd__a22oi_4
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17260_ _17454_/Q _17293_/A2 _17258_/X _17259_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17454_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14472_ _14531_/B _14472_/B vssd1 vssd1 vccd1 vccd1 _14473_/C sky130_fd_sc_hd__or2_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _15235_/A _15235_/C vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16211_ _16107_/Y _16111_/B _16210_/B vssd1 vssd1 vccd1 vccd1 _16300_/B sky130_fd_sc_hd__o21ba_1
X_13423_ _13545_/A _13423_/B _13423_/C vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__nand3_2
X_10635_ _10614_/X _10632_/B _10634_/Y _10550_/X vssd1 vssd1 vccd1 vccd1 _10670_/A
+ sky130_fd_sc_hd__a211o_4
X_17191_ _17191_/A _17191_/B _17191_/C _17191_/D vssd1 vssd1 vccd1 vccd1 _17196_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _16142_/A _16142_/B vssd1 vssd1 vccd1 vccd1 _16143_/B sky130_fd_sc_hd__and2_1
X_13354_ _17415_/A _13866_/D vssd1 vssd1 vccd1 vccd1 _13355_/B sky130_fd_sc_hd__nand2_2
XFILLER_182_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10566_ _10566_/A _10566_/B _10566_/C vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__and3_1
XFILLER_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _12305_/A _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__and3_1
XFILLER_170_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16073_ _16188_/A _16073_/B vssd1 vssd1 vccd1 vccd1 _16075_/B sky130_fd_sc_hd__nor2_1
X_13285_ _13285_/A _13285_/B vssd1 vssd1 vccd1 vccd1 _13292_/A sky130_fd_sc_hd__xnor2_1
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__xnor2_1
X_15024_ _14874_/X _14878_/X _15071_/A vssd1 vssd1 vccd1 vccd1 _15024_/Y sky130_fd_sc_hd__a21oi_4
X_12236_ _12236_/A _12236_/B vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__nor2_4
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12167_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12169_/C sky130_fd_sc_hd__xor2_1
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11118_ _11118_/A _11246_/A vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__nor2_4
X_12098_ _12268_/A _12098_/B _12098_/C vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__nand3_4
X_16975_ _14767_/Y _14929_/X _17163_/A2 _16970_/A _16974_/Y vssd1 vssd1 vccd1 vccd1
+ _16977_/B sky130_fd_sc_hd__o221a_1
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15926_ _15926_/A _15926_/B vssd1 vssd1 vccd1 vccd1 _15927_/B sky130_fd_sc_hd__nand2_1
X_11049_ _11049_/A _11049_/B _11049_/C vssd1 vssd1 vccd1 vccd1 _11051_/C sky130_fd_sc_hd__or3_2
Xinput7 i_wb_addr[13] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ _15858_/A _15858_/B vssd1 vssd1 vccd1 vccd1 _15857_/X sky130_fd_sc_hd__or2_1
XTAP_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14808_ _15622_/B _15623_/A _10269_/X vssd1 vssd1 vccd1 vccd1 _15707_/C sky130_fd_sc_hd__a21o_1
XFILLER_149_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _15788_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _15788_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17527_ fanout930/X _17527_/D vssd1 vssd1 vccd1 vccd1 _17527_/Q sky130_fd_sc_hd__dfxtp_4
X_14739_ _17167_/A _14739_/B vssd1 vssd1 vccd1 vccd1 _14739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17458_ fanout942/X _17458_/D vssd1 vssd1 vccd1 vccd1 _17458_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ _16410_/A _16409_/B vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__nor2_1
X_17389_ _17389_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17389_/X sky130_fd_sc_hd__or2_1
XFILLER_9_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09714_ _16982_/B _09710_/Y _09713_/X vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__o21a_2
XFILLER_142_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _09645_/A _09645_/B _09793_/A vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__nor3_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A _09721_/A vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__nand2_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_24 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _10532_/B _10534_/D _10647_/D _10419_/A vssd1 vssd1 vccd1 vccd1 _10420_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _10345_/A _10343_/Y _10070_/A _10072_/Y vssd1 vssd1 vccd1 vccd1 _10581_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_152_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13070_ _13070_/A _13070_/B vssd1 vssd1 vccd1 vccd1 _13072_/C sky130_fd_sc_hd__xnor2_1
X_10282_ _10134_/Y _10231_/X _10249_/Y _10262_/X vssd1 vssd1 vccd1 vccd1 _10283_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _14952_/B sky130_fd_sc_hd__and2_1
XFILLER_133_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout560 _13390_/S vssd1 vssd1 vccd1 vccd1 _17164_/A sky130_fd_sc_hd__buf_4
Xfanout571 _17513_/Q vssd1 vssd1 vccd1 vccd1 _11268_/A sky130_fd_sc_hd__clkbuf_16
X_16760_ _17119_/A _16760_/B vssd1 vssd1 vccd1 vccd1 _16761_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout582 _11480_/A vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__buf_6
XFILLER_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _14058_/B _13972_/B vssd1 vssd1 vccd1 vccd1 _13974_/A sky130_fd_sc_hd__nand2_4
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout593 _11630_/A vssd1 vssd1 vccd1 vccd1 _11520_/C sky130_fd_sc_hd__buf_4
XFILLER_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15711_ _15711_/A _15711_/B vssd1 vssd1 vccd1 vccd1 _15711_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12923_ _17425_/A _17423_/A _13067_/D _12923_/D vssd1 vssd1 vccd1 vccd1 _12924_/B
+ sky130_fd_sc_hd__and4_1
X_16691_ _16601_/A _16614_/B _16601_/B vssd1 vssd1 vccd1 vccd1 _16693_/B sky130_fd_sc_hd__a21boi_1
XFILLER_111_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15642_ _16226_/C _16812_/A _16745_/B _15726_/A vssd1 vssd1 vccd1 vccd1 _15643_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _14734_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _12854_/Y sky130_fd_sc_hd__nand2_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11802_/Y _11804_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15573_ _15573_/A _15573_/B vssd1 vssd1 vccd1 vccd1 _15584_/A sky130_fd_sc_hd__xnor2_4
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12655_/A _12655_/B _12671_/B _12670_/B _12670_/A vssd1 vssd1 vccd1 vccd1
+ _12822_/B sky130_fd_sc_hd__a32o_2
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _17485_/Q _17328_/A2 _17311_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17485_/D
+ sky130_fd_sc_hd__o211a_1
X_14524_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14583_/A sky130_fd_sc_hd__or3_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _11736_/A _11736_/B _11735_/Y vssd1 vssd1 vccd1 vccd1 _11739_/B sky130_fd_sc_hd__nor3b_2
XFILLER_30_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17243_ _17590_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__a21o_1
X_14455_ _14509_/C _14455_/B vssd1 vssd1 vccd1 vccd1 _14456_/C sky130_fd_sc_hd__and2_1
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11667_ _11686_/B _11686_/A vssd1 vssd1 vccd1 vccd1 _11690_/A sky130_fd_sc_hd__and2b_1
XFILLER_179_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13406_ _13406_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13408_/A sky130_fd_sc_hd__nor2_4
X_10618_ _10963_/A _10963_/B _10920_/B _10962_/B vssd1 vssd1 vccd1 vccd1 _10621_/A
+ sky130_fd_sc_hd__and4_1
X_17174_ input19/X input22/X input21/X input23/X vssd1 vssd1 vccd1 vccd1 _17181_/B
+ sky130_fd_sc_hd__or4b_1
X_14386_ _14386_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__nor2_4
X_11598_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__xor2_4
X_16125_ _16125_/A vssd1 vssd1 vccd1 vccd1 _17558_/D sky130_fd_sc_hd__inv_2
XFILLER_6_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13337_ _13337_/A _13455_/A _13337_/C vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__nor3_2
XFILLER_127_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10549_ _10671_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10550_/C sky130_fd_sc_hd__and2_2
XFILLER_170_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16056_ _16056_/A _16352_/B _16454_/A vssd1 vssd1 vccd1 vccd1 _16058_/A sky130_fd_sc_hd__and3_1
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13268_ _13268_/A _13268_/B vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15007_ _11675_/C _11655_/A _14793_/Y _15108_/A _15006_/Y vssd1 vssd1 vccd1 vccd1
+ _15007_/X sky130_fd_sc_hd__o311a_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ _12213_/X _12218_/Y _17369_/A vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13199_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13200_/B sky130_fd_sc_hd__nor3_1
XFILLER_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16958_ _16958_/A _16958_/B vssd1 vssd1 vccd1 vccd1 _17012_/B sky130_fd_sc_hd__xor2_4
X_15909_ _15884_/Y _15885_/Y _15884_/A vssd1 vssd1 vccd1 vccd1 _15994_/A sky130_fd_sc_hd__o21ai_4
XFILLER_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16889_ _16888_/A _16888_/B _16888_/C vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__a21o_2
X_09430_ _09427_/Y _09430_/B vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__and2b_2
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09361_ _09360_/A _17466_/D _09502_/C vssd1 vssd1 vccd1 vccd1 _09361_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_75_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _09292_/A _09437_/A vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__nand2_2
XFILLER_21_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_12 _17609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_23 _17453_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _15116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_1039 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_45 _09470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_56 _17304_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 _17497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_78 _17452_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_89 _09654_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _09628_/A _09628_/B _09628_/C vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__or3_4
XFILLER_189_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09559_ _09559_/A _09559_/B vssd1 vssd1 vccd1 vccd1 _09689_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12570_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12572_/C sky130_fd_sc_hd__xor2_2
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _11521_/A _11565_/A vssd1 vssd1 vccd1 vccd1 _11523_/B sky130_fd_sc_hd__nor2_4
XFILLER_157_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14240_ _14318_/B _14641_/D _14545_/C _14450_/A vssd1 vssd1 vccd1 vccd1 _14242_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11452_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__or2_4
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10403_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10405_/C sky130_fd_sc_hd__a21oi_4
X_14171_ _14171_/A _14245_/B vssd1 vssd1 vccd1 vccd1 _14173_/C sky130_fd_sc_hd__nor2_2
X_11383_ _11395_/B _11383_/B _11383_/C vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__nand3_4
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10334_ _10451_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__xnor2_4
X_13122_ _13121_/A _13121_/B _13121_/C vssd1 vssd1 vccd1 vccd1 _13123_/B sky130_fd_sc_hd__o21a_1
XFILLER_152_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13053_ _12907_/A _13947_/B _12908_/A _12905_/X vssd1 vssd1 vccd1 vccd1 _13055_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_127_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10267_/C sky130_fd_sc_hd__xnor2_2
XFILLER_105_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _12200_/B _12004_/B vssd1 vssd1 vccd1 vccd1 _12007_/A sky130_fd_sc_hd__nor2_4
XFILLER_87_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10196_ _10321_/A _09172_/B _10062_/B _12487_/B vssd1 vssd1 vccd1 vccd1 _10198_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16812_ _16812_/A _16938_/B _16938_/D _16883_/C vssd1 vssd1 vccd1 vccd1 _16816_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_121_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout390 _12500_/A vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__buf_4
X_16743_ _16814_/B _16809_/C _16743_/C _17043_/B vssd1 vssd1 vccd1 vccd1 _16744_/B
+ sky130_fd_sc_hd__and4_1
X_13955_ _14134_/A _13955_/B vssd1 vssd1 vccd1 vccd1 _13958_/C sky130_fd_sc_hd__and2_1
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ _12749_/Y _13182_/C _12905_/X vssd1 vssd1 vccd1 vccd1 _12908_/A sky130_fd_sc_hd__a21oi_4
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16674_ _16751_/B _16674_/B vssd1 vssd1 vccd1 vccd1 _16677_/B sky130_fd_sc_hd__nand2_1
X_13886_ _13779_/B _13781_/B _13779_/A vssd1 vssd1 vccd1 vccd1 _13888_/B sky130_fd_sc_hd__o21ba_2
XFILLER_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _10269_/X _15804_/A2 _15713_/B1 _15624_/A vssd1 vssd1 vccd1 vccd1 _15625_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12837_ _12833_/Y _12835_/X _12651_/A _12655_/A vssd1 vssd1 vccd1 vccd1 _12837_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_62_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15556_ _16226_/B _16246_/A vssd1 vssd1 vccd1 vccd1 _15557_/B sky130_fd_sc_hd__nand2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12765_/Y _12920_/B _12612_/A _12612_/Y vssd1 vssd1 vccd1 vccd1 _12782_/B
+ sky130_fd_sc_hd__a211o_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14508_/A _14508_/B vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__nand2b_1
XFILLER_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11719_ _11719_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__and2_1
X_15487_ _15406_/A _15406_/B _15403_/X vssd1 vssd1 vccd1 vccd1 _15489_/B sky130_fd_sc_hd__a21o_4
X_12699_ _13003_/A _12698_/B _17070_/B vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17226_ _17552_/Q _17229_/B vssd1 vssd1 vccd1 vccd1 _17226_/X sky130_fd_sc_hd__and2_1
X_14438_ _14438_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14440_/C sky130_fd_sc_hd__nor2_1
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 i_wb_addr[16] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 i_wb_addr[26] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 i_wb_addr[7] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 i_wb_data[16] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput54 i_wb_data[26] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
X_17157_ _17138_/A _17138_/B _10098_/A vssd1 vssd1 vccd1 vccd1 _17157_/Y sky130_fd_sc_hd__a21boi_4
X_14369_ _16965_/C _14641_/D _14368_/C vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__a21oi_1
Xinput65 i_wb_data[7] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_2
XFILLER_157_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16108_ _16114_/A _16108_/B _16108_/C vssd1 vssd1 vccd1 vccd1 _16108_/X sky130_fd_sc_hd__and3b_2
XFILLER_143_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17088_ _17088_/A _17088_/B _17088_/C vssd1 vssd1 vccd1 vccd1 _17089_/B sky130_fd_sc_hd__nor3_1
XFILLER_131_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16039_ _16595_/A _16039_/B vssd1 vssd1 vccd1 vccd1 _16040_/B sky130_fd_sc_hd__nor2_4
X_08930_ _08930_/A _08930_/B _08930_/C vssd1 vssd1 vccd1 vccd1 _08930_/X sky130_fd_sc_hd__or3_4
XFILLER_131_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08861_ _08861_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__xnor2_2
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08792_ _11878_/A _12088_/D _12258_/A _08792_/D vssd1 vssd1 vccd1 vccd1 _11878_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09413_ _12243_/B _09414_/C _09555_/C _12243_/A vssd1 vssd1 vccd1 vccd1 _09415_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_164_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09344_ _09344_/A _09344_/B _09344_/C vssd1 vssd1 vccd1 vccd1 _09344_/Y sky130_fd_sc_hd__nor3_4
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _09275_/A _09275_/B vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__xnor2_2
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ _10050_/A _10050_/B _10163_/A vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__nand3_2
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13740_ _13741_/A _13741_/B _13741_/C vssd1 vssd1 vccd1 vccd1 _13742_/A sky130_fd_sc_hd__o21a_2
X_10952_ _10953_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__or2_4
XFILLER_113_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _13671_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__and3_4
X_10883_ _10883_/A _10883_/B _10883_/C vssd1 vssd1 vccd1 vccd1 _10893_/B sky130_fd_sc_hd__nand3_2
XFILLER_188_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _15140_/Y _15206_/B _15450_/A vssd1 vssd1 vccd1 vccd1 _15497_/B sky130_fd_sc_hd__o21a_4
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _12623_/A _12623_/B vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__nand2_4
X_16390_ _14776_/A _16644_/B _16399_/A vssd1 vssd1 vccd1 vccd1 _16390_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_58_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15341_ _15948_/A _16041_/A vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__nor2_8
XFILLER_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _15457_/B _12553_/B vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__or2_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ _11499_/A _11499_/C _11499_/B vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__o21a_2
X_15272_ _15207_/X _15270_/X _14906_/A vssd1 vssd1 vccd1 vccd1 _15752_/A sky130_fd_sc_hd__a21bo_4
XFILLER_106_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12484_ _12354_/A _12353_/B _12353_/A vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__a21bo_2
XFILLER_185_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17011_ _17014_/A _17014_/B vssd1 vssd1 vccd1 vccd1 _17060_/A sky130_fd_sc_hd__nor2_1
X_14223_ _14599_/B _14485_/D _14360_/C _14680_/A vssd1 vssd1 vccd1 vccd1 _14225_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11435_ _11435_/A _11435_/B _11435_/C vssd1 vssd1 vccd1 vccd1 _11444_/A sky130_fd_sc_hd__nand3_4
XFILLER_172_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14154_ _14154_/A _14154_/B vssd1 vssd1 vccd1 vccd1 _14156_/A sky130_fd_sc_hd__nor2_1
X_11366_ _11341_/A _11341_/B _11341_/C vssd1 vssd1 vccd1 vccd1 _11367_/C sky130_fd_sc_hd__a21oi_2
XFILLER_152_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10317_ _10330_/A _10287_/Y _10303_/Y _10315_/X vssd1 vssd1 vccd1 vccd1 _10319_/C
+ sky130_fd_sc_hd__a211o_2
X_13105_ _13106_/B _13106_/A vssd1 vssd1 vccd1 vccd1 _13236_/B sky130_fd_sc_hd__and2b_1
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14085_ _16864_/A _16918_/A _13998_/B vssd1 vssd1 vccd1 vccd1 _14086_/B sky130_fd_sc_hd__o21ba_1
XFILLER_140_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _11290_/Y _11296_/Y _11153_/C _11235_/X vssd1 vssd1 vccd1 vccd1 _11299_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _13036_/A _13036_/B vssd1 vssd1 vccd1 vccd1 _13038_/A sky130_fd_sc_hd__nor2_1
X_10248_ _10261_/B _10261_/C _10261_/A vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__a21o_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10179_ _10430_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10180_/C sky130_fd_sc_hd__and2_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14987_ _11841_/B _12054_/B _12077_/C _10543_/B _09779_/A _14982_/A vssd1 vssd1 vccd1
+ vccd1 _14988_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16726_ _16568_/A _16568_/B _16641_/A _11762_/X vssd1 vssd1 vccd1 vccd1 _16728_/B
+ sky130_fd_sc_hd__a31oi_2
X_13938_ _13010_/B _13511_/X _13934_/Y _13935_/Y _13937_/X vssd1 vssd1 vccd1 vccd1
+ _13941_/B sky130_fd_sc_hd__a311oi_4
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16657_ _17169_/A1 _16649_/X _16650_/Y _16652_/X _16656_/X vssd1 vssd1 vccd1 vccd1
+ _16657_/X sky130_fd_sc_hd__o311a_1
X_13869_ _13869_/A _13869_/B vssd1 vssd1 vccd1 vccd1 _13870_/B sky130_fd_sc_hd__xnor2_4
XFILLER_179_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _15609_/A _15609_/B _15609_/C vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__o21a_2
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16588_ _16747_/A _16662_/C _16662_/D _16814_/A vssd1 vssd1 vccd1 vccd1 _16590_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15539_ _15901_/S _14989_/X _15538_/X _15806_/B1 vssd1 vssd1 vccd1 vccd1 _15539_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_176_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _09061_/A _09059_/Y _12907_/A _11881_/D vssd1 vssd1 vccd1 vccd1 _09298_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_124_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17437_/Q _17233_/A2 _17207_/X _17208_/X _17428_/B vssd1 vssd1 vccd1 vccd1
+ _17437_/D sky130_fd_sc_hd__o221a_1
XFILLER_162_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ _09813_/X _09829_/Y _09960_/A _09960_/Y vssd1 vssd1 vccd1 vccd1 _09962_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08913_ _12275_/A _12107_/B _13094_/B _13088_/B vssd1 vssd1 vccd1 vccd1 _08916_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _10036_/B _09892_/C _09892_/D _10525_/A vssd1 vssd1 vccd1 vccd1 _09893_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_98_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08845_/B _08845_/A vssd1 vssd1 vccd1 vccd1 _08844_/X sky130_fd_sc_hd__and2b_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08775_ _09030_/A _12638_/B _08776_/C vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__a21oi_2
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09327_ _09462_/A _09326_/Y _15538_/A _11808_/B vssd1 vssd1 vccd1 vccd1 _09468_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_159_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09258_ _09071_/A _09071_/C _09071_/B vssd1 vssd1 vccd1 vccd1 _09259_/B sky130_fd_sc_hd__o21a_1
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09189_ _09189_/A _09221_/A _09189_/C vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__nor3_2
XFILLER_147_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__xnor2_4
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11151_ _11153_/B _11151_/B _11151_/C vssd1 vssd1 vccd1 vccd1 _11153_/C sky130_fd_sc_hd__nor3_4
XFILLER_175_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10102_ _10086_/A _10086_/C _10086_/B vssd1 vssd1 vccd1 vccd1 _10216_/B sky130_fd_sc_hd__o21ai_2
XFILLER_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__xnor2_4
XFILLER_103_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10033_ _10033_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14910_ _17131_/A _15660_/A _15726_/A vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__and3_1
X_15890_ _16809_/A _16108_/B _15898_/A vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__a21bo_1
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14841_ _15457_/B _14841_/B vssd1 vssd1 vccd1 vccd1 _14841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17560_ fanout938/X _17560_/D vssd1 vssd1 vccd1 vccd1 _17560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14772_ _16723_/A _14863_/B vssd1 vssd1 vccd1 vccd1 _16729_/B sky130_fd_sc_hd__or2_1
X_11984_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16511_ _16511_/A _16511_/B vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__or2_1
XFILLER_147_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13723_ _13723_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13726_/A sky130_fd_sc_hd__xnor2_1
X_10935_ _10935_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10936_/B sky130_fd_sc_hd__nor2_4
X_17491_ fanout930/X _17491_/D vssd1 vssd1 vccd1 vccd1 _17491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16442_ _16442_/A _16442_/B vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__xor2_1
X_13654_ _13655_/B _13654_/B vssd1 vssd1 vccd1 vccd1 _13654_/X sky130_fd_sc_hd__and2b_1
XFILLER_140_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10866_ _14786_/A _14787_/A _14848_/A _15175_/B vssd1 vssd1 vccd1 vccd1 _10870_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12607_/C sky130_fd_sc_hd__xnor2_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _16283_/A _16283_/B _16277_/A vssd1 vssd1 vccd1 vccd1 _16375_/B sky130_fd_sc_hd__o21a_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13586_/A _13586_/B _13586_/C vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__o21a_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10797_ _11260_/C _10920_/B vssd1 vssd1 vccd1 vccd1 _10803_/A sky130_fd_sc_hd__nand2_2
XFILLER_158_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15324_ _16226_/C _16136_/B vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__nand2_4
XFILLER_185_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _12536_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__xnor2_4
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15255_ _15245_/X _15252_/X _15254_/X _15253_/X _15537_/A _15806_/B1 vssd1 vssd1
+ vccd1 vccd1 _15255_/X sky130_fd_sc_hd__mux4_1
XFILLER_184_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ _12467_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__and2_1
XFILLER_144_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14206_ _14278_/B _14207_/B vssd1 vssd1 vccd1 vccd1 _14206_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11418_ _11418_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11708_/B sky130_fd_sc_hd__xnor2_4
XFILLER_193_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15186_ _14848_/B _14848_/C _15185_/Y vssd1 vssd1 vccd1 vccd1 _15186_/X sky130_fd_sc_hd__o21a_1
X_12398_ _12040_/Y _12061_/Y _12398_/S vssd1 vssd1 vccd1 vccd1 _12398_/X sky130_fd_sc_hd__mux2_1
X_14137_ _14138_/A _14138_/B vssd1 vssd1 vccd1 vccd1 _14221_/A sky130_fd_sc_hd__nor2_2
XFILLER_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11349_ _11349_/A _11349_/B _11349_/C vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__and3_4
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14068_ _14068_/A _14068_/B vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__xnor2_1
XFILLER_140_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13019_ _13019_/A _13019_/B vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__nor2_2
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16709_ _16709_/A _16709_/B vssd1 vssd1 vccd1 vccd1 _16711_/C sky130_fd_sc_hd__xnor2_2
XFILLER_23_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09112_ _09092_/A _09314_/B _09093_/A vssd1 vssd1 vccd1 vccd1 _09115_/C sky130_fd_sc_hd__o21a_4
XFILLER_148_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09043_/A _17081_/B vssd1 vssd1 vccd1 vccd1 _09044_/B sky130_fd_sc_hd__nand2_2
XFILLER_11_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout901 _10559_/B vssd1 vssd1 vccd1 vccd1 _11605_/B sky130_fd_sc_hd__buf_6
XFILLER_132_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _09945_/A _10064_/A vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__nor2_2
Xfanout912 _17171_/X vssd1 vssd1 vccd1 vccd1 _17266_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout923 _17358_/C1 vssd1 vssd1 vccd1 vccd1 _17290_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout934 fanout936/X vssd1 vssd1 vccd1 vccd1 fanout934/X sky130_fd_sc_hd__clkbuf_4
Xfanout945 fanout946/X vssd1 vssd1 vccd1 vccd1 fanout945/X sky130_fd_sc_hd__buf_4
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09876_/A _10018_/A vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__nor2_2
XTAP_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08893_/A _08826_/B _08826_/A vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__o21ba_1
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08758_ _11027_/A _09892_/C _10993_/D _11867_/A vssd1 vssd1 vccd1 vccd1 _08758_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _10720_/A _11013_/A vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__nor2_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10651_ _10653_/B _10653_/C _10653_/A vssd1 vssd1 vccd1 vccd1 _10651_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ _13369_/B _13369_/C _13369_/A vssd1 vssd1 vccd1 vccd1 _13370_/Y sky130_fd_sc_hd__a21oi_4
X_10582_ _10582_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _12488_/A _12637_/D vssd1 vssd1 vccd1 vccd1 _12323_/C sky130_fd_sc_hd__nand2_1
XFILLER_166_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15040_ _16011_/C _15034_/Y _15037_/X _15039_/X _15035_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15040_/X sky130_fd_sc_hd__mux4_2
XFILLER_181_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12252_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12265_/B sky130_fd_sc_hd__or3_4
XFILLER_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__or2_2
X_12183_ _12183_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12351_/B sky130_fd_sc_hd__nor2_4
XFILLER_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11134_ _11137_/B _11134_/B vssd1 vssd1 vccd1 vccd1 _11135_/C sky130_fd_sc_hd__nor2_1
X_16991_ _16991_/A _16991_/B _16991_/C _16991_/D vssd1 vssd1 vccd1 vccd1 _17046_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15942_ _15837_/A _15837_/B _15826_/Y vssd1 vssd1 vccd1 vccd1 _15944_/B sky130_fd_sc_hd__a21oi_4
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11065_ _11065_/A _11065_/B _11065_/C _11065_/D vssd1 vssd1 vccd1 vccd1 _11065_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10016_ _10017_/A _10015_/Y _10508_/C _10745_/D vssd1 vssd1 vccd1 vccd1 _10140_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_49_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15873_ _16281_/A _16352_/B _15872_/C vssd1 vssd1 vccd1 vccd1 _15874_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17612_ fanout945/X _17612_/D vssd1 vssd1 vccd1 vccd1 _17612_/Q sky130_fd_sc_hd__dfxtp_2
X_14824_ _14767_/Y _16971_/A _16970_/A vssd1 vssd1 vccd1 vccd1 _17024_/A sky130_fd_sc_hd__o21ai_2
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17543_ fanout929/X _17543_/D vssd1 vssd1 vccd1 vccd1 _17543_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _14755_/A _14755_/B vssd1 vssd1 vccd1 vccd1 _14755_/X sky130_fd_sc_hd__or2_1
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _11967_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__nand2_1
XFILLER_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13706_ _13707_/A _13707_/B vssd1 vssd1 vccd1 vccd1 _13706_/Y sky130_fd_sc_hd__nand2_2
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10918_ _10918_/A _10918_/B vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__xnor2_4
X_17474_ fanout928/X _17607_/Q vssd1 vssd1 vccd1 vccd1 _17474_/Q sky130_fd_sc_hd__dfxtp_4
X_14686_ _14719_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14688_/B sky130_fd_sc_hd__xnor2_1
X_11898_ _12138_/B _11898_/B vssd1 vssd1 vccd1 vccd1 _11908_/A sky130_fd_sc_hd__nor2_1
X_16425_ _16425_/A _16425_/B _16423_/Y vssd1 vssd1 vccd1 vccd1 _16426_/B sky130_fd_sc_hd__or3b_2
X_13637_ _13637_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13638_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _10850_/A _10850_/C vssd1 vssd1 vccd1 vccd1 _10855_/B sky130_fd_sc_hd__nor2_2
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16356_ _16356_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16358_/C sky130_fd_sc_hd__xnor2_1
XFILLER_158_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13568_ _13568_/A _13568_/B vssd1 vssd1 vccd1 vccd1 _13569_/C sky130_fd_sc_hd__xnor2_2
XFILLER_185_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15307_ _15307_/A _15307_/B _15307_/C vssd1 vssd1 vccd1 vccd1 _15307_/X sky130_fd_sc_hd__or3_1
XFILLER_146_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12519_ _12519_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__xnor2_2
X_16287_ _16288_/B _16288_/A vssd1 vssd1 vccd1 vccd1 _16287_/Y sky130_fd_sc_hd__nand2b_1
X_13499_ _13500_/A _13500_/B _13500_/C vssd1 vssd1 vccd1 vccd1 _13501_/A sky130_fd_sc_hd__o21a_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15238_ _15238_/A _15796_/B _10419_/A vssd1 vssd1 vccd1 vccd1 _15241_/B sky130_fd_sc_hd__or3b_2
XFILLER_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15169_ _15169_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__xnor2_2
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout208 _12053_/A vssd1 vssd1 vccd1 vccd1 _14912_/B sky130_fd_sc_hd__buf_4
XFILLER_119_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout219 _15638_/Y vssd1 vssd1 vccd1 vccd1 _16745_/B sky130_fd_sc_hd__buf_6
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09730_ _09731_/A _09729_/Y _11902_/A _09892_/D vssd1 vssd1 vccd1 vccd1 _09872_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_86_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _09658_/A _09789_/A _09499_/Y _09500_/X vssd1 vssd1 vccd1 vccd1 _09662_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09592_ _09722_/A _09722_/B vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__and2_2
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_1042 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09026_ _09026_/A _09269_/A vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__nor2_2
XFILLER_156_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout720 _12950_/B vssd1 vssd1 vccd1 vccd1 _11867_/C sky130_fd_sc_hd__buf_6
XFILLER_120_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout731 _11841_/B vssd1 vssd1 vccd1 vccd1 _09892_/C sky130_fd_sc_hd__buf_6
Xfanout742 _10993_/D vssd1 vssd1 vccd1 vccd1 _10534_/D sky130_fd_sc_hd__buf_4
X_09928_ _09929_/A _09927_/Y _09928_/C _09928_/D vssd1 vssd1 vccd1 vccd1 _10184_/A
+ sky130_fd_sc_hd__and4bb_1
Xfanout753 _16114_/A vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__buf_8
Xfanout764 _13434_/C vssd1 vssd1 vccd1 vccd1 _13551_/D sky130_fd_sc_hd__buf_8
Xfanout775 _13196_/B vssd1 vssd1 vccd1 vccd1 _13434_/D sky130_fd_sc_hd__buf_6
Xfanout786 _17490_/Q vssd1 vssd1 vccd1 vccd1 _10791_/D sky130_fd_sc_hd__buf_8
X_09859_ _10255_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__nand2_4
Xfanout797 _15703_/A vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__buf_4
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12870_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__nor2_4
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11821_ _11802_/Y _11804_/Y _11807_/Y _11809_/Y _17365_/A _17367_/A vssd1 vssd1 vccd1
+ vccd1 _11821_/X sky130_fd_sc_hd__mux4_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14763_/S _14538_/X _14585_/B _14483_/Y vssd1 vssd1 vccd1 vccd1 _17599_/D
+ sky130_fd_sc_hd__a31o_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11223_/A _11223_/B _11224_/X vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__a21o_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _11005_/A _10912_/C vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__nand2_4
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14471_/A _14471_/B vssd1 vssd1 vccd1 vccd1 _14472_/B sky130_fd_sc_hd__and2_1
XFILLER_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _15106_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _15235_/C sky130_fd_sc_hd__or2_2
XFILLER_186_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16210_ _16300_/A _16210_/B vssd1 vssd1 vccd1 vccd1 _16210_/Y sky130_fd_sc_hd__nor2_1
X_13422_ _13545_/A _13423_/B _13423_/C vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__and3_2
X_17190_ input9/X input8/X input10/X input16/X vssd1 vssd1 vccd1 vccd1 _17191_/D sky130_fd_sc_hd__or4_1
X_10634_ _10550_/A _10550_/B _10550_/C vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16141_ _16142_/A _16142_/B vssd1 vssd1 vccd1 vccd1 _16241_/B sky130_fd_sc_hd__nor2_2
X_13353_ _13353_/A _13353_/B vssd1 vssd1 vccd1 vccd1 _13355_/A sky130_fd_sc_hd__nor2_1
XFILLER_139_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10565_ _10566_/A _10566_/B _10566_/C vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__a21oi_4
X_12304_ _12305_/A _12305_/B _12305_/C vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__a21oi_4
X_16072_ _16072_/A _16072_/B _16072_/C vssd1 vssd1 vccd1 vccd1 _16073_/B sky130_fd_sc_hd__nor3_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ _13285_/B _13285_/A vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__nand2b_2
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__xor2_1
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15023_ _15081_/A _16025_/A _15415_/A _15734_/A vssd1 vssd1 vccd1 vccd1 _15089_/S
+ sky130_fd_sc_hd__or4_4
X_12235_ _17403_/A _13229_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__and3_2
XFILLER_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12166_ _12166_/A _12166_/B vssd1 vssd1 vccd1 vccd1 _12167_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11118_/A _11116_/Y _11260_/C _14906_/B vssd1 vssd1 vccd1 vccd1 _11246_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12097_ _12268_/A _12098_/B _12098_/C vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__a21o_2
X_16974_ _16974_/A _16974_/B vssd1 vssd1 vccd1 vccd1 _16974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15925_ _15926_/A _15926_/B vssd1 vssd1 vccd1 vccd1 _15925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11051_/B sky130_fd_sc_hd__xor2_2
Xinput8 i_wb_addr[14] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _15666_/B _15853_/A _15756_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _15858_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14807_ _14785_/X _14806_/X _10716_/A vssd1 vssd1 vccd1 vccd1 _15623_/A sky130_fd_sc_hd__a21bo_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15787_ _15883_/B _15787_/B _15788_/B vssd1 vssd1 vccd1 vccd1 _15787_/X sky130_fd_sc_hd__or3b_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ _12999_/A _12999_/B vssd1 vssd1 vccd1 vccd1 _13001_/C sky130_fd_sc_hd__nand2_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14738_ _14738_/A _17153_/A vssd1 vssd1 vccd1 vccd1 _17151_/A sky130_fd_sc_hd__nand2_2
X_17526_ fanout930/X _17526_/D vssd1 vssd1 vccd1 vccd1 _17526_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ fanout942/X _17457_/D vssd1 vssd1 vccd1 vccd1 _17457_/Q sky130_fd_sc_hd__dfxtp_4
X_14669_ _14638_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__and2b_1
XFILLER_20_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16408_ _16108_/C _16317_/B _15209_/Y _16129_/B vssd1 vssd1 vccd1 vccd1 _16411_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17388_ input39/X _17396_/A2 _17387_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17522_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ _16339_/A _16339_/B _16339_/C vssd1 vssd1 vccd1 vccd1 _16340_/B sky130_fd_sc_hd__and3_1
XFILLER_146_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09713_ _10254_/B _10013_/B _10738_/D _09566_/A vssd1 vssd1 vccd1 vccd1 _09713_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09644_ _09645_/B _09793_/A _09645_/A vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__o21a_1
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09575_ _09576_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09721_/A sky130_fd_sc_hd__nand3_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10350_ _17105_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__nor2_1
XFILLER_191_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09009_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10281_ _10275_/X _10388_/A _10266_/X _10267_/Y vssd1 vssd1 vccd1 vccd1 _10283_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_151_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12020_ _12053_/A _12020_/B vssd1 vssd1 vccd1 vccd1 _12020_/Y sky130_fd_sc_hd__nand2_1
XFILLER_183_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout550 _11122_/B vssd1 vssd1 vccd1 vccd1 _10933_/B sky130_fd_sc_hd__buf_6
Xfanout561 _14637_/A1 vssd1 vssd1 vccd1 vccd1 _13390_/S sky130_fd_sc_hd__buf_4
Xfanout572 _09780_/A vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__clkbuf_4
X_13971_ _13971_/A _13971_/B vssd1 vssd1 vccd1 vccd1 _13972_/B sky130_fd_sc_hd__or2_2
XFILLER_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout583 _14792_/A vssd1 vssd1 vccd1 vccd1 _11480_/A sky130_fd_sc_hd__buf_6
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout594 _10899_/C vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__buf_6
XFILLER_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15710_ _16115_/A _15811_/B _15710_/C vssd1 vssd1 vccd1 vccd1 _15710_/X sky130_fd_sc_hd__or3_1
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ _17423_/A _13067_/D _12923_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _12924_/A
+ sky130_fd_sc_hd__a22oi_2
X_16690_ _16690_/A _16690_/B vssd1 vssd1 vccd1 vccd1 _16692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15641_ _15913_/A _16419_/A vssd1 vssd1 vccd1 vccd1 _15732_/A sky130_fd_sc_hd__or2_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _14734_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__and2_2
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _14912_/B _11804_/B vssd1 vssd1 vccd1 vccd1 _11804_/Y sky130_fd_sc_hd__nand2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15572_ _15573_/B _15573_/A vssd1 vssd1 vccd1 vccd1 _15572_/Y sky130_fd_sc_hd__nand2b_2
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12784_ _12781_/X _12938_/B _12784_/B1 _12631_/Y vssd1 vssd1 vccd1 vccd1 _12825_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ input65/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17311_/X sky130_fd_sc_hd__or3_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14577_/A _14523_/B vssd1 vssd1 vccd1 vccd1 _14524_/C sky130_fd_sc_hd__nand2_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11221_/A _11221_/B _11219_/Y vssd1 vssd1 vccd1 vccd1 _11735_/Y sky130_fd_sc_hd__o21ai_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17448_/Q _17290_/A2 _17240_/X _17241_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17448_/D sky130_fd_sc_hd__o221a_1
X_14454_ _14454_/A _14454_/B vssd1 vssd1 vccd1 vccd1 _14455_/B sky130_fd_sc_hd__or2_1
XFILLER_30_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11666_ _11666_/A _11674_/A vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__nor2_2
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13405_ _13852_/A _13405_/B _13844_/D _14002_/B vssd1 vssd1 vccd1 vccd1 _13406_/B
+ sky130_fd_sc_hd__and4_2
X_10617_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__nor2_2
X_17173_ input27/X input26/X input24/X vssd1 vssd1 vccd1 vccd1 _17191_/A sky130_fd_sc_hd__or3b_4
X_14385_ _14450_/A _14641_/C _14509_/A vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__and3_2
X_11597_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__and2_4
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16124_ _16103_/Y _16106_/Y _16123_/X _14871_/Y _16935_/A vssd1 vssd1 vccd1 vccd1
+ _16125_/A sky130_fd_sc_hd__a32o_1
X_13336_ _13337_/A _13455_/A _13337_/C vssd1 vssd1 vccd1 vccd1 _13338_/A sky130_fd_sc_hd__o21a_1
XFILLER_182_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _10547_/A _10547_/B _10547_/C vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__o21ai_1
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16055_ _16055_/A _16827_/D vssd1 vssd1 vccd1 vccd1 _16454_/A sky130_fd_sc_hd__nor2_4
X_13267_ _13002_/A _13134_/Y _13137_/B vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__o21a_1
X_10479_ _11027_/B _10479_/B vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__nand2_2
XFILLER_68_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15006_ _11655_/A _14793_/Y _11675_/C vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12218_ _12218_/A vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13198_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13369_/A sky130_fd_sc_hd__o21a_2
XFILLER_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12149_ _12149_/A _12149_/B vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16957_ _16958_/A _16958_/B vssd1 vssd1 vccd1 vccd1 _17037_/A sky130_fd_sc_hd__nand2b_1
XFILLER_96_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15908_ _15908_/A vssd1 vssd1 vccd1 vccd1 _17556_/D sky130_fd_sc_hd__inv_2
X_16888_ _16888_/A _16888_/B _16888_/C vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__nand3_1
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15839_ _15841_/A _15841_/B vssd1 vssd1 vccd1 vccd1 _15839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09360_ _09360_/A _17466_/D _09502_/C vssd1 vssd1 vccd1 vccd1 _09497_/A sky130_fd_sc_hd__and3_2
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17509_ fanout944/X _17509_/D vssd1 vssd1 vccd1 vccd1 _17509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09291_ _09292_/A _09291_/B _09291_/C vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__nand3_2
XFILLER_178_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_13 _17610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_24 _17435_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 _14213_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 _10559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_68 _17505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _17458_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09627_ _09627_/A _09773_/A vssd1 vssd1 vccd1 vccd1 _09628_/C sky130_fd_sc_hd__nor2_2
XFILLER_46_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09558_ _09558_/A _09558_/B vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__xnor2_4
XFILLER_102_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09489_ _09498_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__xnor2_4
XFILLER_169_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11520_ _11521_/A _11519_/Y _11520_/C _11561_/C vssd1 vssd1 vccd1 vccd1 _11565_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_180_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _11451_/A _11451_/B _11495_/A vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__nor3b_4
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10402_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10402_/Y sky130_fd_sc_hd__nand3_4
XFILLER_183_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14170_ _14170_/A _14245_/A _14170_/C vssd1 vssd1 vccd1 vccd1 _14245_/B sky130_fd_sc_hd__nor3_4
X_11382_ _11376_/A _11376_/C _11376_/B vssd1 vssd1 vccd1 vccd1 _11383_/C sky130_fd_sc_hd__a21o_1
XFILLER_180_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13121_/A _13121_/B _13121_/C vssd1 vssd1 vccd1 vccd1 _13123_/A sky130_fd_sc_hd__nor3_2
X_10333_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__xnor2_4
XFILLER_178_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _13052_/A _13314_/A vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__or2_2
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10264_ _10249_/Y _10262_/X _10134_/Y _10231_/X vssd1 vssd1 vccd1 vccd1 _10283_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_133_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ _12200_/A _12001_/Y _09250_/Y _09255_/B vssd1 vssd1 vccd1 vccd1 _12004_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10195_ _10560_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10322_/A sky130_fd_sc_hd__nand2_2
XFILLER_132_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16811_ _16811_/A _16811_/B vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout380 _17532_/Q vssd1 vssd1 vccd1 vccd1 _12166_/A sky130_fd_sc_hd__buf_6
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout391 _17531_/Q vssd1 vssd1 vccd1 vccd1 _12500_/A sky130_fd_sc_hd__buf_8
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13954_ _13954_/A _13954_/B _13954_/C vssd1 vssd1 vccd1 vccd1 _13955_/B sky130_fd_sc_hd__or3_1
X_16742_ _15658_/Y _16662_/C _16662_/D _16938_/B vssd1 vssd1 vccd1 vccd1 _16744_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _17385_/A _17383_/A _13300_/C _13300_/D vssd1 vssd1 vccd1 vccd1 _12905_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16673_ _16673_/A _16673_/B vssd1 vssd1 vccd1 vccd1 _16674_/B sky130_fd_sc_hd__or2_1
XFILLER_62_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13885_ _13885_/A _13885_/B vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__xor2_4
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12836_ _12651_/A _12655_/A _12833_/Y _12835_/X vssd1 vssd1 vccd1 vccd1 _13001_/B
+ sky130_fd_sc_hd__a211o_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ _15624_/A _15624_/B vssd1 vssd1 vccd1 vccd1 _15624_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _15645_/B _15555_/B vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__xor2_4
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12612_/A _12612_/Y _12765_/Y _12920_/B vssd1 vssd1 vccd1 vccd1 _12938_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14565_/A _14506_/B vssd1 vssd1 vccd1 vccd1 _14508_/B sky130_fd_sc_hd__nor2_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11718_ _11717_/A _16387_/C _11717_/X _16206_/A _11231_/X vssd1 vssd1 vccd1 vccd1
+ _16568_/A sky130_fd_sc_hd__a221o_4
X_15486_ _15486_/A _15486_/B vssd1 vssd1 vccd1 vccd1 _15489_/A sky130_fd_sc_hd__xnor2_4
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12698_ _13003_/A _12698_/B vssd1 vssd1 vccd1 vccd1 _12698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _16965_/C _14641_/C _14437_/C vssd1 vssd1 vccd1 vccd1 _14438_/B sky130_fd_sc_hd__and3_1
X_17225_ _17584_/Q _17270_/A2 _17270_/B1 vssd1 vssd1 vccd1 vccd1 _17225_/X sky130_fd_sc_hd__a21o_1
Xinput11 i_wb_addr[17] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_2
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__xor2_4
XFILLER_174_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput22 i_wb_addr[27] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
Xinput33 i_wb_addr[8] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17156_ _17156_/A _17156_/B _17154_/X vssd1 vssd1 vccd1 vccd1 _17156_/X sky130_fd_sc_hd__or3b_2
Xinput44 i_wb_data[17] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_2
X_14368_ _16965_/C _14641_/D _14368_/C vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__and3_1
Xinput55 i_wb_data[27] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput66 i_wb_data[8] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16107_ _16108_/C _16209_/B _16114_/A vssd1 vssd1 vccd1 vccd1 _16107_/Y sky130_fd_sc_hd__a21boi_4
X_13319_ _13316_/Y _13431_/B _13189_/A _13189_/Y vssd1 vssd1 vccd1 vccd1 _13329_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_192_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17087_ _17088_/A _17088_/B _17088_/C vssd1 vssd1 vccd1 vccd1 _17089_/A sky130_fd_sc_hd__o21a_1
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _14599_/B _14545_/D _14485_/D _14680_/A vssd1 vssd1 vccd1 vccd1 _14302_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_170_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16038_ _15647_/A _16745_/B _15916_/X _15918_/X vssd1 vssd1 vccd1 vccd1 _16044_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_131_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _17381_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__nand2_2
XFILLER_96_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08791_ _12088_/A _12088_/B _11881_/D _11870_/B vssd1 vssd1 vccd1 vccd1 _11878_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09412_ _12245_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _16983_/A sky130_fd_sc_hd__nand2_8
XFILLER_164_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09343_ _09344_/A _09344_/B _09344_/C vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__o21a_4
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09274_ _16982_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09404_/A sky130_fd_sc_hd__xnor2_4
XFILLER_138_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _10951_/A _11065_/A vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__and2_4
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _13671_/A _13671_/B _13671_/C vssd1 vssd1 vccd1 vccd1 _13670_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10882_ _10883_/B _10883_/C _10883_/A vssd1 vssd1 vccd1 vccd1 _10893_/A sky130_fd_sc_hd__a21o_1
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _12621_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__xnor2_4
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15340_ _16315_/C _15948_/A _16041_/A _15081_/A vssd1 vssd1 vccd1 vccd1 _15340_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12552_ _13516_/S _12552_/B vssd1 vssd1 vccd1 vccd1 _12553_/B sky130_fd_sc_hd__or2_2
XFILLER_157_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ _11502_/B _11502_/C _11502_/A vssd1 vssd1 vccd1 vccd1 _11543_/B sky130_fd_sc_hd__o21a_1
X_15271_ _15207_/X _15270_/X _14906_/A vssd1 vssd1 vccd1 vccd1 _16505_/A sky130_fd_sc_hd__a21boi_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12483_ _12479_/Y _12480_/X _12312_/A _12314_/A vssd1 vssd1 vccd1 vccd1 _12522_/B
+ sky130_fd_sc_hd__o211a_1
X_17010_ _17037_/B _17010_/B vssd1 vssd1 vccd1 vccd1 _17014_/B sky130_fd_sc_hd__xor2_4
X_14222_ _14222_/A _14222_/B vssd1 vssd1 vccd1 vccd1 _14262_/A sky130_fd_sc_hd__nand2_1
XFILLER_138_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11434_ _11433_/B _11433_/C _11433_/A vssd1 vssd1 vccd1 vccd1 _11435_/C sky130_fd_sc_hd__a21bo_2
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14153_ _14153_/A _14153_/B _14153_/C _14215_/B vssd1 vssd1 vccd1 vccd1 _14154_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_138_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ _11447_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__or2_2
XFILLER_153_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13104_ _12964_/A _12966_/B _12964_/B vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__o21ba_2
X_10316_ _10303_/Y _10315_/X _10330_/A _10287_/Y vssd1 vssd1 vccd1 vccd1 _10330_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14084_ _14084_/A _14084_/B vssd1 vssd1 vccd1 vccd1 _14087_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11296_ _11345_/A _11345_/B vssd1 vssd1 vccd1 vccd1 _11296_/Y sky130_fd_sc_hd__nand2b_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13658_/A _13298_/A _13169_/D _13908_/B vssd1 vssd1 vccd1 vccd1 _13036_/B
+ sky130_fd_sc_hd__and4_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ _10358_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10261_/C sky130_fd_sc_hd__nand2_2
XFILLER_152_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10178_ _09928_/C _09928_/D _09929_/A _09927_/Y vssd1 vssd1 vccd1 vccd1 _10184_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14986_ _15100_/A _14986_/B vssd1 vssd1 vccd1 vccd1 _14986_/Y sky130_fd_sc_hd__nand2_1
X_16725_ _16791_/A _16723_/Y _16643_/A _16648_/C vssd1 vssd1 vccd1 vccd1 _16725_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13937_ _13727_/A _13825_/Y _13826_/Y _13936_/Y vssd1 vssd1 vccd1 vccd1 _13937_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13868_ _14215_/A _14050_/D vssd1 vssd1 vccd1 vccd1 _13869_/B sky130_fd_sc_hd__nand2_4
X_16656_ _16582_/A _15246_/X _16653_/X _16655_/X vssd1 vssd1 vccd1 vccd1 _16656_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15607_ _15607_/A _15607_/B vssd1 vssd1 vccd1 vccd1 _15609_/C sky130_fd_sc_hd__xor2_2
XFILLER_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12819_ _12820_/A _12820_/B _12820_/C vssd1 vssd1 vccd1 vccd1 _12819_/X sky130_fd_sc_hd__a21o_2
X_16587_ _16566_/A _16566_/B _16560_/A vssd1 vssd1 vccd1 vccd1 _16639_/A sky130_fd_sc_hd__o21ai_2
X_13799_ _13800_/A _13800_/B _13800_/C vssd1 vssd1 vccd1 vccd1 _13801_/A sky130_fd_sc_hd__a21oi_2
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15538_ _15538_/A _15538_/B vssd1 vssd1 vccd1 vccd1 _15538_/X sky130_fd_sc_hd__or2_1
XFILLER_187_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15469_ _15450_/A _16008_/C1 _15468_/X vssd1 vssd1 vccd1 vccd1 _17551_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17208_ _17546_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17208_/X sky130_fd_sc_hd__and2_1
X_17139_ _17139_/A _17139_/B vssd1 vssd1 vccd1 vccd1 _17140_/C sky130_fd_sc_hd__nor2_1
XFILLER_116_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09961_ _09960_/A _09960_/Y _09813_/X _09829_/Y vssd1 vssd1 vccd1 vccd1 _09964_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_170_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08918_/A sky130_fd_sc_hd__nor2_2
XFILLER_98_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _10525_/A _10036_/B _09892_/C _09892_/D vssd1 vssd1 vccd1 vccd1 _09895_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08843_/A _08912_/A vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08774_ _08780_/B _08780_/A vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__and2b_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ _12135_/B _09926_/B _10180_/B _12135_/A vssd1 vssd1 vccd1 vccd1 _09326_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_90_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09257_ _09257_/A _09257_/B vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__xnor2_4
XFILLER_182_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09188_ _09189_/A _09221_/A _09189_/C vssd1 vssd1 vccd1 vccd1 _09190_/A sky130_fd_sc_hd__o21a_1
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11150_ _11145_/A _11145_/B _11145_/C vssd1 vssd1 vccd1 vccd1 _11151_/C sky130_fd_sc_hd__a21oi_4
XFILLER_190_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10101_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__nor2_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11081_ _11080_/B _11145_/A _11064_/X _11071_/Y vssd1 vssd1 vccd1 vccd1 _11084_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_191_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10032_ _09910_/B _10030_/Y _10027_/C _10010_/A vssd1 vssd1 vccd1 vccd1 _10033_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14840_ _14840_/A _14840_/B vssd1 vssd1 vccd1 vccd1 _14840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14771_ _14771_/A _14863_/A vssd1 vssd1 vccd1 vccd1 _16796_/B sky130_fd_sc_hd__or2_1
XFILLER_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11983_ _11984_/A _11984_/B vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__and2b_1
XFILLER_84_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16510_ _16616_/A _16510_/B vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__or2_1
X_13722_ _13723_/A _13723_/B vssd1 vssd1 vccd1 vccd1 _13824_/B sky130_fd_sc_hd__or2_1
XFILLER_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10934_ _10933_/B _11132_/C _10933_/D _10933_/A vssd1 vssd1 vccd1 vccd1 _10935_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_17_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17490_ fanout931/X _17490_/D vssd1 vssd1 vccd1 vccd1 _17490_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16441_ _16442_/A _16442_/B vssd1 vssd1 vccd1 vccd1 _16550_/A sky130_fd_sc_hd__nand2_1
X_13653_ _13543_/A _13543_/B _13537_/Y vssd1 vssd1 vccd1 vccd1 _13654_/B sky130_fd_sc_hd__o21bai_1
XFILLER_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10865_ _10865_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__xnor2_4
X_12604_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12764_/B sky130_fd_sc_hd__nand2b_2
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _16372_/A _16372_/B vssd1 vssd1 vccd1 vccd1 _16375_/A sky130_fd_sc_hd__xnor2_4
XFILLER_176_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _13584_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13586_/C sky130_fd_sc_hd__xnor2_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10901_/B _10796_/B _10860_/B vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__or3_4
XFILLER_185_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _14906_/A _16008_/C1 _15322_/X vssd1 vssd1 vccd1 vccd1 _17549_/D sky130_fd_sc_hd__a21oi_4
XFILLER_169_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12535_ _12331_/Y _12333_/B _12336_/A vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__a21oi_4
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15254_ _14992_/Y _14998_/Y _15254_/S vssd1 vssd1 vccd1 vccd1 _15254_/X sky130_fd_sc_hd__mux2_1
X_12466_ _12467_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__nor2_2
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ _14279_/A _14205_/B vssd1 vssd1 vccd1 vccd1 _14207_/B sky130_fd_sc_hd__and2b_1
X_11417_ _11418_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__and2b_2
X_15185_ _14848_/B _14848_/C _16115_/A vssd1 vssd1 vccd1 vccd1 _15185_/Y sky130_fd_sc_hd__a21oi_1
X_12397_ _15095_/B _12397_/B vssd1 vssd1 vccd1 vccd1 _13837_/C sky130_fd_sc_hd__or2_1
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14136_ _14218_/B _14136_/B vssd1 vssd1 vccd1 vccd1 _14138_/B sky130_fd_sc_hd__or2_1
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11348_ _11348_/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11349_/C sky130_fd_sc_hd__and2_2
XFILLER_98_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _14068_/A _14068_/B vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__and2b_1
XFILLER_152_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11279_ _11561_/B _15703_/A _15530_/A _11561_/A vssd1 vssd1 vccd1 vccd1 _11280_/B
+ sky130_fd_sc_hd__a22oi_1
X_13018_ _17403_/A _17399_/A _14215_/B _13564_/C vssd1 vssd1 vccd1 vccd1 _13019_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14969_ _14899_/X _14968_/X _08727_/Y vssd1 vssd1 vccd1 vccd1 _14969_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16708_ _16709_/B _16709_/A vssd1 vssd1 vccd1 vccd1 _16784_/B sky130_fd_sc_hd__nand2b_1
XFILLER_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16639_ _16639_/A _16854_/C vssd1 vssd1 vccd1 vccd1 _16639_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09111_ _09153_/B _09111_/B vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__or2_4
XFILLER_148_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09042_ _17387_/A _11867_/D vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__nand2_2
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09944_ _09945_/A _09943_/Y _10062_/A _09944_/D vssd1 vssd1 vccd1 vccd1 _10064_/A
+ sky130_fd_sc_hd__and4bb_1
Xfanout902 _10559_/B vssd1 vssd1 vccd1 vccd1 _11370_/D sky130_fd_sc_hd__buf_4
Xfanout913 _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17392_/C1 sky130_fd_sc_hd__buf_4
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout924 _08730_/Y vssd1 vssd1 vccd1 vccd1 _17358_/C1 sky130_fd_sc_hd__buf_6
XFILLER_48_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout935 fanout937/X vssd1 vssd1 vccd1 vccd1 fanout935/X sky130_fd_sc_hd__clkbuf_2
Xfanout946 input2/X vssd1 vssd1 vccd1 vccd1 fanout946/X sky130_fd_sc_hd__buf_6
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _09876_/A _09874_/Y _10508_/C _10036_/D vssd1 vssd1 vccd1 vccd1 _10018_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08826_/A _08826_/B vssd1 vssd1 vccd1 vccd1 _08893_/B sky130_fd_sc_hd__nor2_2
XFILLER_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__xor2_4
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ _10735_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _10653_/C sky130_fd_sc_hd__nand2_2
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ _09303_/X _09439_/A _09316_/A _09296_/Y vssd1 vssd1 vccd1 vccd1 _09316_/B
+ sky130_fd_sc_hd__o211ai_4
X_10581_ _10581_/A _10581_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _11771_/B sky130_fd_sc_hd__or3_2
XFILLER_167_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12320_ _12487_/A _12487_/B _12659_/B _13194_/D vssd1 vssd1 vccd1 vccd1 _12492_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_182_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12251_ _12252_/A _12252_/B _12252_/C vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__o21ai_4
XFILLER_181_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__and2_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__xor2_4
X_11133_ _11561_/B _11132_/C _11334_/C _14922_/S vssd1 vssd1 vccd1 vccd1 _11134_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_122_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16990_ _16990_/A _16990_/B vssd1 vssd1 vccd1 vccd1 _16991_/D sky130_fd_sc_hd__nand2_2
XFILLER_123_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15941_ _15941_/A _15941_/B vssd1 vssd1 vccd1 vccd1 _15944_/A sky130_fd_sc_hd__xnor2_4
XFILLER_150_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11064_ _11065_/A _11065_/B _11065_/C _11065_/D vssd1 vssd1 vccd1 vccd1 _11064_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10015_ _14784_/A _10743_/C _10640_/D _10392_/A vssd1 vssd1 vccd1 vccd1 _10015_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15872_ _15872_/A _16352_/B _15872_/C vssd1 vssd1 vccd1 vccd1 _15989_/B sky130_fd_sc_hd__and3_1
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17611_ fanout945/X _17611_/D vssd1 vssd1 vccd1 vccd1 _17611_/Q sky130_fd_sc_hd__dfxtp_1
X_14823_ _16918_/B _16918_/C _14080_/C vssd1 vssd1 vccd1 vccd1 _16971_/A sky130_fd_sc_hd__a21oi_2
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ fanout926/X _17542_/D vssd1 vssd1 vccd1 vccd1 _17542_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14754_ _14755_/A _14755_/B vssd1 vssd1 vccd1 vccd1 _14754_/Y sky130_fd_sc_hd__nand2_1
X_11966_ _11965_/B _11966_/B vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__nand2b_1
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13705_ _13705_/A _13705_/B vssd1 vssd1 vccd1 vccd1 _13707_/B sky130_fd_sc_hd__xnor2_2
X_10917_ _10918_/B _10918_/A vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__and2b_2
X_14685_ _14710_/C _14710_/B _14684_/A vssd1 vssd1 vccd1 vccd1 _14686_/B sky130_fd_sc_hd__a21oi_1
X_17473_ fanout928/X _17546_/Q vssd1 vssd1 vccd1 vccd1 _17473_/Q sky130_fd_sc_hd__dfxtp_2
X_11897_ _12104_/A _12270_/D _11894_/Y _12138_/A vssd1 vssd1 vccd1 vccd1 _11898_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13636_ _13635_/A _13741_/A _13635_/C vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__o21ai_2
X_16424_ _16425_/A _16425_/B _16423_/A _16509_/B vssd1 vssd1 vccd1 vccd1 _16527_/A
+ sky130_fd_sc_hd__o211a_2
X_10848_ _15116_/A _15206_/A _10836_/A _10834_/Y vssd1 vssd1 vccd1 vccd1 _10850_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_158_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16355_ _16536_/A _16355_/B vssd1 vssd1 vccd1 vccd1 _16356_/B sky130_fd_sc_hd__nand2_1
X_13567_ _14387_/A _14213_/C _13568_/A vssd1 vssd1 vccd1 vccd1 _13695_/B sky130_fd_sc_hd__and3_1
XFILLER_185_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10779_ _10779_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__xnor2_4
XFILLER_157_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12518_ _12518_/A _12518_/B vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__xnor2_4
X_15306_ _15241_/B _15241_/C _15241_/A vssd1 vssd1 vccd1 vccd1 _15307_/C sky130_fd_sc_hd__a21boi_2
X_16286_ _16189_/B _16191_/B _16187_/Y vssd1 vssd1 vccd1 vccd1 _16288_/B sky130_fd_sc_hd__o21a_1
X_13498_ _13498_/A _13498_/B vssd1 vssd1 vccd1 vccd1 _13500_/C sky130_fd_sc_hd__xnor2_1
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12449_ _12276_/A _12278_/B _12276_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__o21ba_2
X_15237_ _10419_/A _15373_/B _15238_/A vssd1 vssd1 vccd1 vccd1 _15241_/A sky130_fd_sc_hd__a21bo_1
XFILLER_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15168_ _15169_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15168_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_158_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14119_ _14119_/A _14119_/B _14117_/X vssd1 vssd1 vccd1 vccd1 _14120_/B sky130_fd_sc_hd__or3b_1
XFILLER_140_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15099_ _14863_/A _14864_/A _11808_/B _09652_/B _10430_/A _14958_/A vssd1 vssd1 vccd1
+ vccd1 _15100_/B sky130_fd_sc_hd__mux4_1
Xfanout209 _12053_/A vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _09499_/Y _09500_/X _09658_/A _09789_/A vssd1 vssd1 vccd1 vccd1 _09662_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09591_ _09591_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09722_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09025_ _09026_/A _09024_/Y _09025_/C _09509_/B vssd1 vssd1 vccd1 vccd1 _09269_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_152_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout710 _16571_/A vssd1 vssd1 vccd1 vccd1 _13564_/D sky130_fd_sc_hd__buf_8
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout721 _12054_/B vssd1 vssd1 vccd1 vccd1 _12950_/B sky130_fd_sc_hd__clkbuf_16
Xfanout732 _12068_/C vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__buf_6
XFILLER_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _09926_/A _10309_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09927_/Y sky130_fd_sc_hd__a21oi_1
Xfanout743 _14859_/B vssd1 vssd1 vccd1 vccd1 _10993_/D sky130_fd_sc_hd__buf_6
Xfanout754 _16114_/A vssd1 vssd1 vccd1 vccd1 _15204_/A sky130_fd_sc_hd__buf_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout765 _16683_/A vssd1 vssd1 vccd1 vccd1 _16880_/A sky130_fd_sc_hd__clkbuf_8
Xfanout776 _16758_/A vssd1 vssd1 vccd1 vccd1 _16807_/A sky130_fd_sc_hd__clkbuf_8
Xfanout787 _14901_/B vssd1 vssd1 vccd1 vccd1 _16938_/A sky130_fd_sc_hd__buf_8
X_09858_ _10255_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _16809_/B sky130_fd_sc_hd__and2_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout798 _11135_/B vssd1 vssd1 vccd1 vccd1 _15703_/A sky130_fd_sc_hd__buf_12
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _08815_/B _08815_/A vssd1 vssd1 vccd1 vccd1 _08831_/B sky130_fd_sc_hd__and2b_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09790_/B sky130_fd_sc_hd__nor2_1
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11820_/A vssd1 vssd1 vccd1 vccd1 _11820_/Y sky130_fd_sc_hd__inv_2
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11739_/B _11739_/C _11739_/A vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__o21ai_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10702_ _10905_/A _10905_/B _11005_/B _10805_/D vssd1 vssd1 vccd1 vccd1 _10705_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14470_ _14471_/A _14471_/B vssd1 vssd1 vccd1 vccd1 _14531_/B sky130_fd_sc_hd__nor2_1
XFILLER_159_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11681_/A _11678_/A _11681_/B _11662_/B _11680_/Y vssd1 vssd1 vccd1 vccd1
+ _11683_/B sky130_fd_sc_hd__a311o_1
XFILLER_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13421_ _13545_/A _13423_/B _13423_/C vssd1 vssd1 vccd1 vccd1 _13421_/Y sky130_fd_sc_hd__a21oi_4
X_10633_ _10632_/A _10632_/Y _10519_/Y _10588_/X vssd1 vssd1 vccd1 vccd1 wire120/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_128_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16140_ _16140_/A _16140_/B vssd1 vssd1 vccd1 vccd1 _16142_/B sky130_fd_sc_hd__xor2_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13352_ _14765_/A _14766_/A _13764_/D _13664_/D vssd1 vssd1 vccd1 vccd1 _13353_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10564_ _10564_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10566_/C sky130_fd_sc_hd__nand2_2
XFILLER_127_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12303_ _12303_/A _12303_/B vssd1 vssd1 vccd1 vccd1 _12305_/C sky130_fd_sc_hd__xnor2_4
X_16071_ _16072_/A _16072_/B _16072_/C vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__o21a_1
X_13283_ _13149_/A _13151_/B _13149_/B vssd1 vssd1 vccd1 vccd1 _13285_/B sky130_fd_sc_hd__o21ba_1
X_10495_ _10496_/B _10496_/A vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__nand2b_2
X_15022_ _15918_/A _15278_/A _15821_/A _15660_/A vssd1 vssd1 vccd1 vccd1 _15030_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ _17403_/A _13229_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _12236_/A sky130_fd_sc_hd__a21oi_2
XFILLER_107_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12165_ _12165_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11116_ _11258_/B _11563_/D _11561_/D _11115_/A vssd1 vssd1 vccd1 vccd1 _11116_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_123_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12096_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12098_/C sky130_fd_sc_hd__xnor2_4
X_16973_ _14865_/B _16868_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _16973_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_122_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15924_ _16036_/A _15924_/B vssd1 vssd1 vccd1 vccd1 _15926_/B sky130_fd_sc_hd__or2_1
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11047_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11047_/Y sky130_fd_sc_hd__nor2_2
XFILLER_65_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput9 i_wb_addr[15] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15855_ _15855_/A _15855_/B vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__xnor2_4
XFILLER_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14806_ _14806_/A _15456_/A vssd1 vssd1 vccd1 vccd1 _14806_/X sky130_fd_sc_hd__or2_2
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _15786_/A _15786_/B vssd1 vssd1 vccd1 vccd1 _15788_/B sky130_fd_sc_hd__or2_4
XFILLER_33_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12998_ _12997_/A _12997_/B _12997_/C vssd1 vssd1 vccd1 vccd1 _12999_/B sky130_fd_sc_hd__o21ai_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17525_ fanout930/X _17525_/D vssd1 vssd1 vccd1 vccd1 _17525_/Q sky130_fd_sc_hd__dfxtp_1
X_14737_ _17167_/A _14739_/B vssd1 vssd1 vccd1 vccd1 _14737_/X sky130_fd_sc_hd__or2_1
XFILLER_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11949_ _09016_/A _09016_/Y _11947_/X _11948_/Y vssd1 vssd1 vccd1 vccd1 _11949_/Y
+ sky130_fd_sc_hd__a211oi_4
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17456_ fanout942/X _17456_/D vssd1 vssd1 vccd1 vccd1 _17456_/Q sky130_fd_sc_hd__dfxtp_2
X_14668_ _17164_/A _12394_/A _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14668_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_177_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16407_ _16407_/A vssd1 vssd1 vccd1 vccd1 _17561_/D sky130_fd_sc_hd__inv_2
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13619_ _13619_/A _13619_/B vssd1 vssd1 vccd1 vccd1 _13621_/B sky130_fd_sc_hd__nand2_1
X_17387_ _17387_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17387_/X sky130_fd_sc_hd__or2_1
X_14599_ _14599_/A _14599_/B _14708_/C _14599_/D vssd1 vssd1 vccd1 vccd1 _14600_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_125_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16338_ _16339_/A _16339_/B _16339_/C vssd1 vssd1 vccd1 vccd1 _16444_/A sky130_fd_sc_hd__a21oi_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16269_ _16270_/A _16270_/B _16270_/C vssd1 vssd1 vccd1 vccd1 _16271_/A sky130_fd_sc_hd__o21a_1
XFILLER_145_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09712_ _10255_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__nand2_4
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _10067_/A _09937_/B _09643_/C vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__and3_1
XFILLER_95_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09574_ _09574_/A _09574_/B _09574_/C vssd1 vssd1 vccd1 vccd1 _09575_/C sky130_fd_sc_hd__or3_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__or2_4
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10280_ _10266_/X _10267_/Y _10275_/X _10388_/A vssd1 vssd1 vccd1 vccd1 _10283_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout540 _09470_/B vssd1 vssd1 vccd1 vccd1 _12135_/B sky130_fd_sc_hd__buf_6
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout551 fanout554/X vssd1 vssd1 vccd1 vccd1 _11122_/B sky130_fd_sc_hd__buf_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout562 _11268_/A vssd1 vssd1 vccd1 vccd1 _14637_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13970_ _13971_/A _13971_/B vssd1 vssd1 vccd1 vccd1 _14058_/B sky130_fd_sc_hd__nand2_2
Xfanout573 _10431_/A vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__clkbuf_4
Xfanout584 _17512_/Q vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout595 _12214_/A vssd1 vssd1 vccd1 vccd1 _10899_/C sky130_fd_sc_hd__buf_2
XFILLER_24_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12921_ _12920_/A _12920_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12933_/B sky130_fd_sc_hd__a21oi_4
XFILLER_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15640_ _16812_/A _16745_/B vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__nand2_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _17164_/A _12852_/B vssd1 vssd1 vccd1 vccd1 _12852_/X sky130_fd_sc_hd__or2_4
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11803_ _17363_/A _10431_/B _10309_/C vssd1 vssd1 vccd1 vccd1 _11804_/B sky130_fd_sc_hd__a21o_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _15486_/A _15486_/B _15483_/Y vssd1 vssd1 vccd1 vccd1 _15573_/B sky130_fd_sc_hd__o21a_2
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12784_/B1 _12631_/Y _12781_/X _12938_/B vssd1 vssd1 vccd1 vccd1 _12825_/A
+ sky130_fd_sc_hd__o211a_4
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _12463_/D _17328_/A2 _17309_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17484_/D
+ sky130_fd_sc_hd__o211a_1
X_14522_ _14519_/X _14520_/Y _14463_/B _14465_/A vssd1 vssd1 vccd1 vccd1 _14523_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11731_/B _11729_/C _11729_/B vssd1 vssd1 vccd1 vccd1 _11736_/B sky130_fd_sc_hd__o21a_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17557_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__and2_1
XFILLER_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14453_ _14454_/A _14454_/B vssd1 vssd1 vccd1 vccd1 _14509_/C sky130_fd_sc_hd__nand2_1
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11665_ _11673_/A _11673_/B vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__and2_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13404_ _13405_/B _13844_/D _14002_/B _13852_/A vssd1 vssd1 vccd1 vccd1 _13406_/A
+ sky130_fd_sc_hd__a22oi_4
X_10616_ _10508_/C _10970_/B _10509_/A _10507_/Y vssd1 vssd1 vccd1 vccd1 _10617_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14384_ _14450_/A _14641_/C _14509_/A vssd1 vssd1 vccd1 vccd1 _14386_/A sky130_fd_sc_hd__a21oi_2
X_17172_ input69/X input68/X input35/X vssd1 vssd1 vccd1 vccd1 _17172_/Y sky130_fd_sc_hd__nand3b_1
X_11596_ _11630_/A _15116_/B _11628_/B _11593_/Y vssd1 vssd1 vccd1 vccd1 _11598_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_167_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ _14387_/A _13564_/D vssd1 vssd1 vccd1 vccd1 _13337_/C sky130_fd_sc_hd__nand2_1
X_16123_ _17169_/A1 _16112_/X _16113_/Y _16122_/X _16111_/X vssd1 vssd1 vccd1 vccd1
+ _16123_/X sky130_fd_sc_hd__o311a_1
X_10547_ _10547_/A _10547_/B _10547_/C vssd1 vssd1 vccd1 vccd1 _10671_/A sky130_fd_sc_hd__or3_1
XFILLER_170_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16054_ _16935_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16827_/D sky130_fd_sc_hd__nand2_4
XFILLER_157_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ _13266_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _13271_/A sky130_fd_sc_hd__xnor2_1
X_10478_ _10478_/A _10478_/B vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__nor2_2
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12217_ _17367_/A _12217_/B vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__nor2_4
X_15005_ _14941_/X _15002_/X _15003_/X _15004_/Y _15309_/B vssd1 vssd1 vccd1 vccd1
+ _15005_/X sky130_fd_sc_hd__a311o_1
XFILLER_68_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13197_ _13197_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13199_/C sky130_fd_sc_hd__xnor2_1
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/B sky130_fd_sc_hd__and3_1
XFILLER_29_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16956_ _16900_/A _16900_/C _16900_/B vssd1 vssd1 vccd1 vccd1 _16958_/B sky130_fd_sc_hd__a21bo_2
XFILLER_38_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12079_ _12079_/A _13094_/B vssd1 vssd1 vccd1 vccd1 _12080_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15907_ _16807_/A _16806_/A2 _15887_/Y _15906_/X vssd1 vssd1 vccd1 vccd1 _15908_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16887_ _16887_/A _16887_/B vssd1 vssd1 vccd1 vccd1 _16888_/C sky130_fd_sc_hd__or2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15838_ _15741_/A _15741_/B _15731_/X vssd1 vssd1 vccd1 vccd1 _15841_/B sky130_fd_sc_hd__o21a_1
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15769_ _15769_/A _15769_/B _15769_/C vssd1 vssd1 vccd1 vccd1 _15776_/B sky130_fd_sc_hd__nor3_1
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17508_ fanout944/X _17508_/D vssd1 vssd1 vccd1 vccd1 _17508_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09290_ _09290_/A _09290_/B _09290_/C vssd1 vssd1 vccd1 vccd1 _09291_/C sky130_fd_sc_hd__nand3_1
XFILLER_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_14 _17544_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ fanout937/X _17439_/D vssd1 vssd1 vccd1 vccd1 _17439_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_25 _17454_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_36 _17411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_58 fanout944/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 _17528_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_554 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput110 _17438_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ _09626_/A _09629_/B _09626_/C vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__and3_2
XFILLER_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09557_ _12245_/A _12158_/C vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__nand2_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09488_ _09388_/A _09486_/Y _09484_/B _09460_/X vssd1 vssd1 vccd1 vccd1 _09488_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_93_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ _11403_/B _11400_/B _11400_/C vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__a21oi_4
XFILLER_165_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10401_ _10402_/A _10402_/B _10402_/C vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__and3_2
XFILLER_109_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11381_ _11380_/A _11426_/A vssd1 vssd1 vccd1 vccd1 _11383_/B sky130_fd_sc_hd__nand2b_2
XFILLER_125_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13121_/C sky130_fd_sc_hd__xor2_2
XFILLER_125_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ _10333_/B _10333_/A vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__and2b_1
XFILLER_192_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13051_ _17385_/A _17383_/A _13947_/B _13300_/C vssd1 vssd1 vccd1 vccd1 _13314_/A
+ sky130_fd_sc_hd__and4_2
X_10263_ _10249_/Y _10262_/X _10134_/Y _10231_/X vssd1 vssd1 vccd1 vccd1 _10263_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_87_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12002_ _09250_/Y _09255_/B _12200_/A _12001_/Y vssd1 vssd1 vccd1 vccd1 _12200_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10194_ _10194_/A _10194_/B _10194_/C vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__nor3_2
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16810_ _15801_/A _15658_/Y _16662_/D _16808_/X vssd1 vssd1 vccd1 vccd1 _16811_/B
+ sky130_fd_sc_hd__o31a_1
Xfanout370 _14383_/A vssd1 vssd1 vccd1 vccd1 _14318_/B sky130_fd_sc_hd__buf_6
XFILLER_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout381 _17532_/Q vssd1 vssd1 vccd1 vccd1 _12795_/A sky130_fd_sc_hd__buf_6
X_16741_ _16715_/Y _16717_/Y _16853_/A vssd1 vssd1 vccd1 vccd1 _16787_/A sky130_fd_sc_hd__o21ai_2
Xfanout392 _14008_/A vssd1 vssd1 vccd1 vccd1 _14254_/A sky130_fd_sc_hd__buf_6
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13953_ _14044_/A vssd1 vssd1 vccd1 vccd1 _14134_/A sky130_fd_sc_hd__clkinv_2
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _17383_/A _13300_/C vssd1 vssd1 vccd1 vccd1 _13182_/C sky130_fd_sc_hd__nand2_2
XFILLER_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ _16673_/A _16673_/B vssd1 vssd1 vccd1 vccd1 _16751_/B sky130_fd_sc_hd__nand2_1
X_13884_ _13885_/B _13885_/A vssd1 vssd1 vccd1 vccd1 _13986_/B sky130_fd_sc_hd__and2b_1
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ _15623_/A _15623_/B vssd1 vssd1 vccd1 vccd1 _15623_/X sky130_fd_sc_hd__xor2_2
XFILLER_185_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12835_ _12991_/B _12834_/B _12834_/C vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__o21a_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ _15645_/B _15555_/B vssd1 vssd1 vccd1 vccd1 _15554_/Y sky130_fd_sc_hd__nor2_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ _12766_/A _12928_/B _12766_/C vssd1 vssd1 vccd1 vccd1 _12920_/B sky130_fd_sc_hd__or3_4
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14505_ _14505_/A _14505_/B vssd1 vssd1 vccd1 vccd1 _14506_/B sky130_fd_sc_hd__and2_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11717_/A _16295_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__and3_1
X_15485_ _16136_/B _16536_/A vssd1 vssd1 vccd1 vccd1 _15486_/B sky130_fd_sc_hd__nand2_4
X_12697_ _12379_/B _13004_/A _12695_/X vssd1 vssd1 vccd1 vccd1 _12698_/B sky130_fd_sc_hd__o21a_1
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ _17442_/Q _17233_/A2 _17222_/X _17223_/X _17372_/C1 vssd1 vssd1 vccd1 vccd1
+ _17442_/D sky130_fd_sc_hd__o221a_1
X_14436_ _16965_/C _14318_/C _14437_/C vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__a21oi_1
X_11648_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__xnor2_4
Xinput12 i_wb_addr[18] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 i_wb_addr[28] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput34 i_wb_addr[9] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17155_ _17152_/Y _17153_/X _17133_/A _17136_/X vssd1 vssd1 vccd1 vccd1 _17156_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput45 i_wb_data[18] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_2
X_14367_ _14367_/A _17023_/A vssd1 vssd1 vccd1 vccd1 _14368_/C sky130_fd_sc_hd__xor2_1
X_11579_ _11579_/A _11579_/B _11579_/C vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__nand3_4
Xinput56 i_wb_data[28] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput67 i_wb_data[9] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16106_ _16389_/A _16106_/B vssd1 vssd1 vccd1 vccd1 _16106_/Y sky130_fd_sc_hd__nand2_4
X_13318_ _13189_/A _13189_/Y _13316_/Y _13431_/B vssd1 vssd1 vccd1 vccd1 _13329_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14298_ _14214_/A _14216_/B _14214_/B vssd1 vssd1 vccd1 vccd1 _14306_/A sky130_fd_sc_hd__o21ba_2
XFILLER_143_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17086_ _17086_/A _17086_/B vssd1 vssd1 vccd1 vccd1 _17088_/C sky130_fd_sc_hd__and2_1
XFILLER_182_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _16595_/A _16041_/B _15935_/A _15933_/B vssd1 vssd1 vccd1 vccd1 _16046_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13249_ _13249_/A _13249_/B _13249_/C _13249_/D vssd1 vssd1 vccd1 vccd1 _13249_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_69_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08790_ _08792_/D vssd1 vssd1 vccd1 vccd1 _08790_/Y sky130_fd_sc_hd__inv_2
X_16939_ _16983_/A _16939_/B vssd1 vssd1 vccd1 vccd1 _16986_/A sky130_fd_sc_hd__or2_2
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09411_ _09411_/A _09411_/B _09417_/B vssd1 vssd1 vccd1 vccd1 _09434_/B sky130_fd_sc_hd__or3_2
XFILLER_92_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09344_/C sky130_fd_sc_hd__nor2_2
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09273_ _09273_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__nor2_2
XFILLER_166_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08988_ _12770_/A _11920_/B _11920_/D _10446_/B vssd1 vssd1 vccd1 vccd1 _08989_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ _10857_/Y _10863_/B _10951_/A _10949_/Y vssd1 vssd1 vccd1 vccd1 _11065_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_44_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09609_ _09610_/A _09610_/C vssd1 vssd1 vccd1 vccd1 _09614_/B sky130_fd_sc_hd__nor2_2
X_10881_ _10883_/B _10883_/C _10883_/A vssd1 vssd1 vccd1 vccd1 _10881_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12620_ _12620_/A _12923_/D vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__nand2_4
XFILLER_189_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12551_ _11827_/X _11854_/C _17164_/B vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__mux2_1
XFILLER_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _11502_/A _11502_/B _11502_/C vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__nor3_4
X_15270_ _15270_/A _15270_/B _15270_/C vssd1 vssd1 vccd1 vccd1 _15270_/X sky130_fd_sc_hd__or3_4
X_12482_ _12312_/A _12314_/A _12479_/Y _12480_/X vssd1 vssd1 vccd1 vccd1 _12522_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14221_ _14221_/A _14221_/B _14221_/C vssd1 vssd1 vccd1 vccd1 _14222_/B sky130_fd_sc_hd__or3_1
X_11433_ _11433_/A _11433_/B _11433_/C vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__nand3_2
XFILLER_153_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _14153_/B _14153_/C _14215_/B _14153_/A vssd1 vssd1 vccd1 vccd1 _14154_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_98_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11364_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _10315_/A _10315_/B _10315_/C vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__and3_4
X_13103_ _13103_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__xnor2_1
X_14083_ _14168_/A _14545_/C _14084_/A vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__and3_2
XFILLER_153_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11295_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11345_/B sky130_fd_sc_hd__xnor2_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13298_/A _13169_/D _13908_/B _13658_/A vssd1 vssd1 vccd1 vccd1 _13036_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10246_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10358_/B sky130_fd_sc_hd__xor2_4
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10177_ _10177_/A _10177_/B _10289_/A vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__nand3_4
XFILLER_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14985_ _12245_/B _12021_/B _09928_/D _09926_/B _10542_/A _14982_/A vssd1 vssd1 vccd1
+ vccd1 _14986_/B sky130_fd_sc_hd__mux4_1
XFILLER_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16724_ _16643_/Y _16647_/A _16723_/B _16723_/A _16721_/Y vssd1 vssd1 vccd1 vccd1
+ _16791_/B sky130_fd_sc_hd__a221o_1
X_13936_ _13936_/A _13936_/B _13728_/Y vssd1 vssd1 vccd1 vccd1 _13936_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16655_ _16649_/A _17163_/A2 _16654_/X vssd1 vssd1 vccd1 vccd1 _16655_/X sky130_fd_sc_hd__o21ba_1
X_13867_ _13867_/A _13867_/B vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__nor2_2
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15606_ _15607_/A _15607_/B vssd1 vssd1 vccd1 vccd1 _15606_/Y sky130_fd_sc_hd__nand2_2
X_12818_ _12820_/A _12820_/B _12820_/C vssd1 vssd1 vccd1 vccd1 _12821_/A sky130_fd_sc_hd__a21oi_1
X_16586_ _16571_/A _16806_/A2 _16575_/X _16585_/X vssd1 vssd1 vccd1 vccd1 _17563_/D
+ sky130_fd_sc_hd__a22oi_4
X_13798_ _13906_/B _13798_/B vssd1 vssd1 vccd1 vccd1 _13800_/C sky130_fd_sc_hd__nand2_1
XFILLER_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15537_ _15537_/A _15537_/B vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__or2_2
X_12749_ _17385_/A _13300_/D vssd1 vssd1 vccd1 vccd1 _12749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15468_ _15446_/Y _15447_/X _15467_/X _15445_/X vssd1 vssd1 vccd1 vccd1 _15468_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17207_ _17578_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17207_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14419_ _14533_/A _14419_/B vssd1 vssd1 vccd1 vccd1 _14419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15399_ _15816_/A _15932_/B _16041_/B _15820_/A vssd1 vssd1 vccd1 vccd1 _15400_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17138_ _17138_/A _17138_/B vssd1 vssd1 vccd1 vccd1 _17138_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17069_ _14434_/Y _14764_/Y _14825_/Y _17023_/A vssd1 vssd1 vccd1 vccd1 _17069_/Y
+ sky130_fd_sc_hd__o211ai_1
X_09960_ _09960_/A _09960_/B _09960_/C vssd1 vssd1 vccd1 vccd1 _09960_/Y sky130_fd_sc_hd__nand3_2
XFILLER_171_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08911_ _17381_/A _12088_/C _08843_/A _08841_/Y vssd1 vssd1 vccd1 vccd1 _08912_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__nand2_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08843_/A _08841_/Y _17381_/A _12088_/C vssd1 vssd1 vccd1 vccd1 _08912_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_97_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A _08804_/A vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__nor2_2
XFILLER_111_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _12135_/A _12135_/B _09926_/B _10180_/B vssd1 vssd1 vccd1 vccd1 _09462_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _09256_/A _09256_/B vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__xnor2_4
XFILLER_193_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09187_ _12488_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _09189_/C sky130_fd_sc_hd__nand2_1
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _10090_/A _10088_/X _10081_/A _10084_/A vssd1 vssd1 vccd1 vccd1 _10101_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11080_ _11080_/A _11080_/B _11080_/C _11080_/D vssd1 vssd1 vccd1 vccd1 _11145_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_68_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _10010_/A _10027_/C _10030_/Y _09910_/B vssd1 vssd1 vccd1 vccd1 _10033_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _14770_/A _14864_/A vssd1 vssd1 vccd1 vccd1 _16864_/B sky130_fd_sc_hd__or2_2
X_11982_ _11982_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _11984_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13721_ _13577_/B _13579_/B _13577_/A vssd1 vssd1 vccd1 vccd1 _13723_/B sky130_fd_sc_hd__o21ba_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10933_ _10933_/A _10933_/B _11132_/C _10933_/D vssd1 vssd1 vccd1 vccd1 _10935_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _16331_/A _16331_/B _16345_/A vssd1 vssd1 vccd1 vccd1 _16442_/B sky130_fd_sc_hd__a21o_1
X_13652_ _13652_/A _13652_/B vssd1 vssd1 vccd1 vccd1 _13655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10864_ _10863_/B _10863_/C _10863_/A vssd1 vssd1 vccd1 vccd1 _10864_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12603_ _12603_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__xnor2_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _16372_/B _16372_/A vssd1 vssd1 vccd1 vccd1 _16371_/Y sky130_fd_sc_hd__nand2b_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _14226_/A _16480_/A vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10795_ _10884_/A _10794_/B _10794_/A vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__o21ba_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15322_ _15794_/A _15303_/Y _15321_/X _15301_/Y vssd1 vssd1 vccd1 vccd1 _15322_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__xnor2_4
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15253_ _14988_/Y _14999_/Y _15384_/S vssd1 vssd1 vccd1 vccd1 _15253_/X sky130_fd_sc_hd__mux2_1
X_12465_ _12772_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__nand2_1
XFILLER_184_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14204_ _14204_/A _14279_/B vssd1 vssd1 vccd1 vccd1 _14278_/B sky130_fd_sc_hd__or2_1
XFILLER_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11416_ _11416_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__or2_4
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15184_ _14790_/Y _14929_/X _15713_/B1 _14848_/B vssd1 vssd1 vccd1 vccd1 _15184_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12396_ _12388_/X _14210_/A _14840_/A vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__mux2_1
XFILLER_137_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14135_ _14134_/A _14134_/B _14134_/C vssd1 vssd1 vccd1 vccd1 _14136_/B sky130_fd_sc_hd__o21a_1
X_11347_ _11347_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__nand2_1
XFILLER_193_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14066_ _14066_/A _14066_/B vssd1 vssd1 vccd1 vccd1 _14068_/B sky130_fd_sc_hd__xnor2_2
X_11278_ _11561_/A _15703_/A _11387_/C vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__and3_2
X_13017_ _17399_/A _14215_/B _13564_/C _17403_/A vssd1 vssd1 vccd1 vccd1 _13019_/A
+ sky130_fd_sc_hd__a22oi_4
X_10229_ _10192_/B _10207_/B _10192_/D _10193_/A vssd1 vssd1 vccd1 vccd1 _10229_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_79_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14968_ _14966_/X _14967_/X _15143_/A vssd1 vssd1 vccd1 vccd1 _14968_/X sky130_fd_sc_hd__a21o_4
X_16707_ _16542_/A _16626_/B _16624_/X vssd1 vssd1 vccd1 vccd1 _16709_/B sky130_fd_sc_hd__a21oi_4
X_13919_ _14018_/B _13919_/B vssd1 vssd1 vccd1 vccd1 _13921_/C sky130_fd_sc_hd__nand2_1
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14899_ _14899_/A _14906_/B _14899_/C vssd1 vssd1 vccd1 vccd1 _14899_/X sky130_fd_sc_hd__or3_4
X_16638_ _16638_/A _16638_/B vssd1 vssd1 vccd1 vccd1 _16854_/C sky130_fd_sc_hd__xnor2_4
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16569_ _16568_/A _16568_/B _16207_/B _16568_/Y vssd1 vssd1 vccd1 vccd1 _16569_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09110_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09041_ _09043_/A _17081_/B vssd1 vssd1 vccd1 vccd1 _09041_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09943_ _09942_/A _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _09943_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout903 _10559_/B vssd1 vssd1 vccd1 vccd1 _11027_/D sky130_fd_sc_hd__buf_8
Xfanout914 _17322_/C1 vssd1 vssd1 vccd1 vccd1 _17380_/C1 sky130_fd_sc_hd__buf_4
Xfanout925 fanout926/X vssd1 vssd1 vccd1 vccd1 fanout925/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout936 fanout937/X vssd1 vssd1 vccd1 vccd1 fanout936/X sky130_fd_sc_hd__buf_4
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _14784_/A _10645_/C _10412_/C _10392_/A vssd1 vssd1 vccd1 vccd1 _09874_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08825_ _12088_/B _11867_/C _11867_/D _12088_/A vssd1 vssd1 vccd1 vccd1 _08826_/B
+ sky130_fd_sc_hd__a22oi_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08756_ _08757_/B _08757_/A vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__nand2b_2
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09308_ _09316_/A _09296_/Y _09303_/X _09439_/A vssd1 vssd1 vccd1 vccd1 _09311_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_167_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _10582_/A _10582_/B vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__or2_1
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09239_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09240_/B sky130_fd_sc_hd__nor2_1
XFILLER_182_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12250_ _12250_/A _12250_/B vssd1 vssd1 vccd1 vccd1 _12252_/C sky130_fd_sc_hd__xnor2_4
XFILLER_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _16387_/A sky130_fd_sc_hd__xnor2_4
XFILLER_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _11978_/A _11980_/B _11978_/B vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__o21ba_4
XFILLER_123_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _11561_/A _11561_/B _11132_/C _11334_/C vssd1 vssd1 vccd1 vccd1 _11137_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15940_ _16072_/B _15940_/B vssd1 vssd1 vccd1 vccd1 _15941_/B sky130_fd_sc_hd__nor2_4
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11063_ _11061_/A _11061_/C _11077_/A vssd1 vssd1 vccd1 vccd1 _11065_/D sky130_fd_sc_hd__a21o_2
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _10392_/A _14784_/A _10412_/C _10640_/D vssd1 vssd1 vccd1 vccd1 _10017_/A
+ sky130_fd_sc_hd__and4_2
X_15871_ _15871_/A _15871_/B vssd1 vssd1 vccd1 vccd1 _15872_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17610_ fanout926/X _17610_/D vssd1 vssd1 vccd1 vccd1 _17610_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14822_ _16864_/B _16865_/A _16864_/A vssd1 vssd1 vccd1 vccd1 _16918_/C sky130_fd_sc_hd__a21bo_1
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17541_ fanout944/X _17541_/D vssd1 vssd1 vccd1 vccd1 _17541_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14701_/A _14701_/B _14725_/Y _14752_/Y vssd1 vssd1 vccd1 vccd1 _14755_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11965_ _11966_/B _11965_/B vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__nand2b_4
XFILLER_45_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13704_ _14254_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _13705_/B sky130_fd_sc_hd__nand2_1
XFILLER_189_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17472_ fanout928/X _17545_/Q vssd1 vssd1 vccd1 vccd1 _17472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10916_ _10808_/A _10807_/B _10807_/A vssd1 vssd1 vccd1 vccd1 _10918_/B sky130_fd_sc_hd__o21ba_2
X_14684_ _14684_/A vssd1 vssd1 vccd1 vccd1 _14719_/B sky130_fd_sc_hd__inv_2
XFILLER_44_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11896_ _11894_/Y _12138_/A _12104_/A _12270_/D vssd1 vssd1 vccd1 vccd1 _12138_/B
+ sky130_fd_sc_hd__and4bb_2
X_16423_ _16423_/A _16509_/B vssd1 vssd1 vccd1 vccd1 _16423_/Y sky130_fd_sc_hd__nand2_1
X_13635_ _13635_/A _13741_/A _13635_/C vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__or3_2
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _10828_/A _10827_/B _10827_/A vssd1 vssd1 vccd1 vccd1 _10855_/A sky130_fd_sc_hd__o21ba_4
X_16354_ _16354_/A _16354_/B vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13566_ _14387_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13568_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _10778_/A _11742_/A vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__nor2_4
XFILLER_185_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15305_ _15314_/A _15373_/B _15305_/C vssd1 vssd1 vccd1 vccd1 _15307_/B sky130_fd_sc_hd__and3b_1
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12517_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12518_/B sky130_fd_sc_hd__xnor2_4
XFILLER_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16285_ _16285_/A _16285_/B vssd1 vssd1 vccd1 vccd1 _16288_/A sky130_fd_sc_hd__xor2_2
XFILLER_173_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13497_ _13498_/B _13498_/A vssd1 vssd1 vccd1 vccd1 _13497_/X sky130_fd_sc_hd__and2b_2
XFILLER_173_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15236_ _15235_/B _15235_/C _15235_/A vssd1 vssd1 vccd1 vccd1 _15236_/X sky130_fd_sc_hd__a21o_1
XFILLER_172_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12448_ _12448_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12451_/A sky130_fd_sc_hd__xnor2_4
X_15167_ _15089_/S _15687_/A _15170_/B vssd1 vssd1 vccd1 vccd1 _15169_/B sky130_fd_sc_hd__o21ai_4
X_12379_ _12696_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__or2_4
XFILLER_158_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14118_ _14119_/A _14119_/B _14117_/X vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__o21ba_1
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15098_ _17164_/D _15097_/X _15130_/S vssd1 vssd1 vccd1 vccd1 _15715_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14049_ _14050_/B _14141_/D _14050_/D _14050_/A vssd1 vssd1 vccd1 vccd1 _14051_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_79_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09590_ _09750_/C _10311_/D _09473_/A _09465_/Y vssd1 vssd1 vccd1 vccd1 _09591_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09024_ _09023_/B _09555_/C _09647_/B _09023_/A vssd1 vssd1 vccd1 vccd1 _09024_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_117_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout700 _14052_/B vssd1 vssd1 vccd1 vccd1 _13564_/C sky130_fd_sc_hd__buf_8
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout711 _17498_/Q vssd1 vssd1 vccd1 vccd1 _16571_/A sky130_fd_sc_hd__buf_8
X_09926_ _09926_/A _09926_/B _09926_/C vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__and3_1
Xfanout722 _10753_/B vssd1 vssd1 vccd1 vccd1 _10659_/D sky130_fd_sc_hd__buf_4
XFILLER_104_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout733 _16298_/A vssd1 vssd1 vccd1 vccd1 _13866_/D sky130_fd_sc_hd__clkbuf_16
Xfanout744 _17494_/Q vssd1 vssd1 vccd1 vccd1 _14859_/B sky130_fd_sc_hd__buf_6
Xfanout755 _17119_/A vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__clkbuf_4
Xfanout766 _16014_/A vssd1 vssd1 vccd1 vccd1 _16683_/A sky130_fd_sc_hd__buf_4
Xfanout777 _15898_/A vssd1 vssd1 vccd1 vccd1 _16758_/A sky130_fd_sc_hd__clkbuf_8
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09710_/Y _09856_/Y _09855_/X vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__a21o_2
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout788 _17490_/Q vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__buf_4
Xfanout799 _17489_/Q vssd1 vssd1 vccd1 vccd1 _11135_/B sky130_fd_sc_hd__buf_6
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _08808_/A _08883_/A vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__nor2_2
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__and2_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _17607_/Q _17608_/Q vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__nand2b_4
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__xor2_4
XFILLER_92_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__xor2_4
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _15235_/B sky130_fd_sc_hd__or2_1
X_13420_ _13420_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13423_/C sky130_fd_sc_hd__xnor2_4
X_10632_ _10632_/A _10632_/B _10632_/C _10632_/D vssd1 vssd1 vccd1 vccd1 _10632_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_179_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13351_ _14766_/A _13764_/D _13664_/D _14765_/A vssd1 vssd1 vccd1 vccd1 _13353_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10563_ _10563_/A _10563_/B vssd1 vssd1 vccd1 vccd1 _10564_/B sky130_fd_sc_hd__or2_1
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _17373_/A _12592_/C _12470_/B vssd1 vssd1 vccd1 vccd1 _12303_/B sky130_fd_sc_hd__and3_2
X_16070_ _16070_/A _16070_/B vssd1 vssd1 vccd1 vccd1 _16072_/C sky130_fd_sc_hd__xnor2_1
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13282_ _13282_/A _13282_/B vssd1 vssd1 vccd1 vccd1 _13285_/A sky130_fd_sc_hd__xnor2_2
XFILLER_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10601_/A _10493_/B _10493_/A vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__o21ba_1
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15021_ _15401_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15734_/A sky130_fd_sc_hd__nand2_4
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12233_ _17399_/A _13966_/D vssd1 vssd1 vccd1 vccd1 _12235_/C sky130_fd_sc_hd__and2_4
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12164_ _12163_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__o21a_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11115_ _11115_/A _11258_/B _11377_/C _11561_/D vssd1 vssd1 vccd1 vccd1 _11118_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12095_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12286_/B sky130_fd_sc_hd__nand2b_2
X_16972_ _16972_/A _16972_/B vssd1 vssd1 vccd1 vccd1 _16972_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15923_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _15924_/B sky130_fd_sc_hd__and2_1
X_11046_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__nand2_2
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15854_ _16171_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _15855_/B sky130_fd_sc_hd__nand2_4
XFILLER_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14805_ _14805_/A _14805_/B _14805_/C vssd1 vssd1 vccd1 vccd1 _15456_/A sky130_fd_sc_hd__and3_1
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _15883_/B _15787_/B vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__or2_4
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ _12997_/A _12997_/B _12997_/C vssd1 vssd1 vccd1 vccd1 _12999_/A sky130_fd_sc_hd__or3_2
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17524_ fanout931/X _17524_/D vssd1 vssd1 vccd1 vccd1 _17524_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _14736_/A _14744_/A vssd1 vssd1 vccd1 vccd1 _14739_/B sky130_fd_sc_hd__nand2_1
X_11948_ _11917_/X _11918_/Y _12156_/B _11947_/D vssd1 vssd1 vccd1 vccd1 _11948_/Y
+ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ fanout942/X _17455_/D vssd1 vssd1 vccd1 vccd1 _17455_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14667_ _14667_/A _14667_/B vssd1 vssd1 vccd1 vccd1 _14667_/Y sky130_fd_sc_hd__nand2_1
X_11879_ _08760_/Y _16302_/A _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _11886_/A
+ sky130_fd_sc_hd__o22ai_4
X_16406_ _16386_/Y _16389_/Y _16405_/X _16806_/A2 _16399_/A vssd1 vssd1 vccd1 vccd1
+ _16407_/A sky130_fd_sc_hd__a32o_1
XFILLER_177_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13618_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13729_/B sky130_fd_sc_hd__xnor2_2
XFILLER_193_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17386_ input38/X _17396_/A2 _17385_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17521_/D
+ sky130_fd_sc_hd__o211a_1
X_14598_ _14599_/B _14708_/C _14599_/D _14680_/A vssd1 vssd1 vccd1 vccd1 _14600_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16337_ _16337_/A _16337_/B vssd1 vssd1 vccd1 vccd1 _16339_/C sky130_fd_sc_hd__xnor2_1
X_13549_ _13662_/B _13547_/X _13425_/Y _13430_/A vssd1 vssd1 vccd1 vccd1 _13558_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _16268_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16270_/C sky130_fd_sc_hd__xnor2_1
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15219_ _15220_/A _15220_/B vssd1 vssd1 vccd1 vccd1 _15287_/A sky130_fd_sc_hd__nand2b_4
X_16199_ _16200_/A _16200_/B _16200_/C vssd1 vssd1 vccd1 vccd1 _16382_/A sky130_fd_sc_hd__a21oi_4
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09711_ _10255_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__and2_1
XFILLER_101_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09643_/C sky130_fd_sc_hd__xnor2_1
XFILLER_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09573_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__xnor2_2
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09007_ _09007_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__xnor2_1
XFILLER_152_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout530 _09470_/A vssd1 vssd1 vccd1 vccd1 _08718_/A sky130_fd_sc_hd__buf_8
Xfanout541 _12847_/A vssd1 vssd1 vccd1 vccd1 _14421_/S sky130_fd_sc_hd__buf_6
X_09909_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__and3_2
Xfanout552 fanout554/X vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__buf_6
Xfanout563 _11268_/A vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__buf_6
Xfanout574 _15254_/S vssd1 vssd1 vccd1 vccd1 _10431_/A sky130_fd_sc_hd__buf_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout585 _12214_/A vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__buf_6
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout596 _17511_/Q vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__clkbuf_8
X_12920_ _12920_/A _12920_/B _12920_/C vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__and3_2
XFILLER_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12851_ _12220_/X _12229_/C _16011_/B vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11802_ _14912_/B _11802_/B vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__nand2_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15570_/A _15570_/B vssd1 vssd1 vccd1 vccd1 _15573_/A sky130_fd_sc_hd__xor2_4
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12938_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12938_/B sky130_fd_sc_hd__nand3_4
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14463_/B _14465_/A _14519_/X _14520_/Y vssd1 vssd1 vccd1 vccd1 _14577_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11732_/B _11732_/C _11732_/A vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__o21a_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17589_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17240_/X sky130_fd_sc_hd__a21o_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14387_/A _14708_/C _14388_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14454_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11673_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13403_ _13403_/A _13403_/B vssd1 vssd1 vccd1 vccd1 _13409_/A sky130_fd_sc_hd__nand2_2
X_10615_ _10615_/A _10615_/B _10615_/C vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__nand3_2
X_17171_ input69/X input68/X input35/X vssd1 vssd1 vccd1 vccd1 _17171_/X sky130_fd_sc_hd__and3b_1
X_14383_ _14383_/A _14708_/D vssd1 vssd1 vccd1 vccd1 _14509_/A sky130_fd_sc_hd__and2_2
X_11595_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__xnor2_4
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16122_ _16122_/A _16122_/B _16122_/C vssd1 vssd1 vccd1 vccd1 _16122_/X sky130_fd_sc_hd__and3_1
XFILLER_183_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13334_ _16913_/C _14383_/A _13450_/D _13966_/D vssd1 vssd1 vccd1 vccd1 _13455_/A
+ sky130_fd_sc_hd__and4_2
X_10546_ _10546_/A _10655_/A vssd1 vssd1 vccd1 vccd1 _10547_/C sky130_fd_sc_hd__nor2_1
XFILLER_155_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16053_ _16935_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16695_/B sky130_fd_sc_hd__and2_4
XFILLER_143_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265_ _13266_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__or2_1
X_10477_ _10694_/A _10694_/B _17469_/D _17468_/D vssd1 vssd1 vccd1 vccd1 _10478_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15004_ _15002_/X _15003_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _15004_/Y sky130_fd_sc_hd__a21oi_1
X_12216_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__inv_2
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13196_ _17421_/A _13196_/B vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12147_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__a21oi_2
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16955_ _16955_/A _16955_/B vssd1 vssd1 vccd1 vccd1 _16958_/A sky130_fd_sc_hd__xnor2_4
X_12078_ _12078_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11029_ _11032_/A _11029_/B _11025_/Y vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__or3b_4
X_15906_ _16207_/B _15889_/Y _15894_/X _15905_/X vssd1 vssd1 vccd1 vccd1 _15906_/X
+ sky130_fd_sc_hd__o211a_1
X_16886_ _16886_/A _16886_/B vssd1 vssd1 vccd1 vccd1 _16887_/B sky130_fd_sc_hd__and2_1
X_15837_ _15837_/A _15837_/B vssd1 vssd1 vccd1 vccd1 _15841_/A sky130_fd_sc_hd__xnor2_2
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15768_ _15769_/A _15769_/B _15769_/C vssd1 vssd1 vccd1 vccd1 _15877_/A sky130_fd_sc_hd__o21a_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14719_ _14719_/A _14719_/B _14719_/C vssd1 vssd1 vccd1 vccd1 _14747_/B sky130_fd_sc_hd__or3_1
XFILLER_75_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17507_ fanout944/X _17507_/D vssd1 vssd1 vccd1 vccd1 _17507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15699_ _15610_/Y _15611_/X _15610_/A vssd1 vssd1 vccd1 vccd1 _15700_/B sky130_fd_sc_hd__a21oi_2
XFILLER_177_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17438_ fanout934/X _17438_/D vssd1 vssd1 vccd1 vccd1 _17438_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _17546_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _17456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 _17411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ _17369_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17369_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_59 _17515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput100 _17458_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput111 _17439_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_161_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09625_ _09627_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09626_/C sky130_fd_sc_hd__nor2_1
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _09556_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _09460_/X _09484_/B _09486_/Y _09388_/A vssd1 vssd1 vccd1 vccd1 _09487_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_54_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ _10501_/A _10501_/B _10396_/X vssd1 vssd1 vccd1 vccd1 _10402_/C sky130_fd_sc_hd__a21o_2
XFILLER_164_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11380_ _11380_/A _11380_/B _11380_/C vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__or3_2
XFILLER_176_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10331_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__xor2_4
XFILLER_191_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13050_ _17383_/A _13947_/B _13300_/C _17385_/A vssd1 vssd1 vccd1 vccd1 _13052_/A
+ sky130_fd_sc_hd__a22oi_1
X_10262_ _10262_/A _10262_/B _10262_/C vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__and3_4
XFILLER_140_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _11998_/X _11999_/Y _09122_/A _09255_/X vssd1 vssd1 vccd1 vccd1 _12001_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10193_ _10193_/A _10193_/B vssd1 vssd1 vccd1 vccd1 _10194_/C sky130_fd_sc_hd__nor2_1
XFILLER_160_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout360 _17413_/A vssd1 vssd1 vccd1 vccd1 _14769_/A sky130_fd_sc_hd__buf_8
Xfanout371 _13895_/B vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__buf_12
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16740_ _16722_/A _17170_/B1 _16719_/Y _16739_/X vssd1 vssd1 vccd1 vccd1 _17565_/D
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout382 _10560_/A vssd1 vssd1 vccd1 vccd1 _10067_/A sky130_fd_sc_hd__clkbuf_4
X_13952_ _13954_/A _13954_/B _13954_/C vssd1 vssd1 vccd1 vccd1 _14044_/A sky130_fd_sc_hd__o21a_1
Xfanout393 _17405_/A vssd1 vssd1 vccd1 vccd1 _14008_/A sky130_fd_sc_hd__buf_4
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _12903_/A _12903_/B vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__or2_1
X_16671_ _16671_/A _16671_/B vssd1 vssd1 vccd1 vccd1 _16673_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13883_ _13774_/A _13776_/B _13774_/B vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__o21ba_2
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15622_ _15622_/A _15622_/B vssd1 vssd1 vccd1 vccd1 _15623_/B sky130_fd_sc_hd__nand2_1
X_12834_ _12991_/B _12834_/B _12834_/C vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__or3_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15553_ _15553_/A _15553_/B _16827_/B vssd1 vssd1 vccd1 vccd1 _15555_/B sky130_fd_sc_hd__or3_4
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12928_/B _12766_/C _12766_/A vssd1 vssd1 vccd1 vccd1 _12765_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14505_/A _14505_/B vssd1 vssd1 vccd1 vccd1 _14565_/A sky130_fd_sc_hd__nor2_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11302_/B _16294_/A _11302_/A vssd1 vssd1 vccd1 vccd1 _16387_/C sky130_fd_sc_hd__o21a_2
X_15484_ _15484_/A _15567_/A vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__xnor2_4
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__or2_1
XFILLER_187_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17223_ _17551_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17223_/X sky130_fd_sc_hd__and2_1
X_14435_ _17023_/A _14492_/A _14432_/X vssd1 vssd1 vccd1 vccd1 _14437_/C sky130_fd_sc_hd__o21a_1
X_11647_ _11624_/A _11624_/B _15524_/B _15524_/C vssd1 vssd1 vccd1 vccd1 _15525_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 i_wb_addr[19] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17154_ _17133_/A _17136_/X _17152_/Y _17153_/X vssd1 vssd1 vccd1 vccd1 _17154_/X
+ sky130_fd_sc_hd__a211o_1
Xinput24 i_wb_addr[29] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_2
X_14366_ _14599_/B _17028_/A vssd1 vssd1 vccd1 vccd1 _17023_/A sky130_fd_sc_hd__nand2_8
XFILLER_168_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 i_wb_cyc vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_8
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11578_ _11574_/A _11574_/C _11607_/A vssd1 vssd1 vccd1 vccd1 _11579_/C sky130_fd_sc_hd__o21ai_4
Xinput46 i_wb_data[19] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
Xinput57 i_wb_data[29] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
Xinput68 i_wb_stb vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_6
X_16105_ _16105_/A _16105_/B vssd1 vssd1 vccd1 vccd1 _16106_/B sky130_fd_sc_hd__xor2_4
X_13317_ _13317_/A _13317_/B _13317_/C vssd1 vssd1 vccd1 vccd1 _13431_/B sky130_fd_sc_hd__and3_4
X_17085_ _17085_/A _17085_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17086_/B sky130_fd_sc_hd__or3_1
XFILLER_128_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10529_ _10647_/C _10755_/D _10422_/A _10420_/Y vssd1 vssd1 vccd1 vccd1 _10531_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_14297_ _14297_/A _14297_/B vssd1 vssd1 vccd1 vccd1 _14337_/A sky130_fd_sc_hd__xor2_4
XFILLER_182_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16036_ _16036_/A _16036_/B vssd1 vssd1 vccd1 vccd1 _16048_/A sky130_fd_sc_hd__xnor2_2
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ _13248_/A _13248_/B _13248_/C vssd1 vssd1 vccd1 vccd1 _13249_/D sky130_fd_sc_hd__or3_2
XFILLER_124_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _13046_/A _13047_/B _13177_/Y _13312_/B vssd1 vssd1 vccd1 vccd1 _13189_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_111_411 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16938_ _16938_/A _16938_/B _16939_/B _16938_/D vssd1 vssd1 vccd1 vccd1 _16994_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16869_ _16864_/B _17162_/A2 _16974_/B _14864_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16869_/X sky130_fd_sc_hd__a221o_1
X_09410_ _09410_/A _09548_/A vssd1 vssd1 vccd1 vccd1 _09417_/B sky130_fd_sc_hd__nor2_4
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09341_ _09214_/A _09214_/B _09214_/C vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09272_ _12243_/A _12243_/B _12659_/B _09414_/C vssd1 vssd1 vccd1 vccd1 _09273_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_179_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08987_ _11920_/B _11920_/D _10446_/B _12770_/A vssd1 vssd1 vccd1 vccd1 _08989_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_130_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _15537_/A _14864_/A _09602_/A _09471_/Y vssd1 vssd1 vccd1 vccd1 _09610_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_189_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _11114_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _10883_/C sky130_fd_sc_hd__nand2_2
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09539_ _09531_/X _09532_/Y _09487_/X _09530_/B vssd1 vssd1 vccd1 vccd1 _09540_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12550_ _12545_/X _12549_/X _17371_/A vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ _11456_/X _11490_/Y _11499_/A _11539_/A vssd1 vssd1 vccd1 vccd1 _11502_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_169_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12481_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12481_/Y sky130_fd_sc_hd__nand3_2
X_14220_ _14221_/A _14221_/B _14221_/C vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__o21ai_4
XFILLER_156_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11432_ _11426_/A _11426_/C _11426_/B vssd1 vssd1 vccd1 vccd1 _11433_/C sky130_fd_sc_hd__a21o_1
XFILLER_149_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14151_ _14151_/A _14151_/B vssd1 vssd1 vccd1 vccd1 _14190_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__nand2b_1
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102_ _13103_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__and2b_1
XFILLER_180_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10315_/C sky130_fd_sc_hd__xnor2_4
X_14082_ _14168_/A _14545_/C vssd1 vssd1 vccd1 vccd1 _14084_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11294_ _11299_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__nand2_4
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13033_ _13033_/A _13033_/B _13033_/C vssd1 vssd1 vccd1 vccd1 _13046_/B sky130_fd_sc_hd__nand3_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10245_ _10245_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10358_/A sky130_fd_sc_hd__xnor2_4
XFILLER_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10176_ _10177_/B _10289_/A _10177_/A vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__a21o_4
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14984_ _15252_/B _14983_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _15537_/B sky130_fd_sc_hd__mux2_1
Xfanout190 _15263_/Y vssd1 vssd1 vccd1 vccd1 _16533_/A sky130_fd_sc_hd__buf_6
XFILLER_47_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16723_ _16723_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _16723_/Y sky130_fd_sc_hd__nand2_1
X_13935_ _13935_/A _13935_/B _13510_/X vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__nor3b_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16654_ _16649_/B _17162_/A2 _16974_/B _12245_/B _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16654_/X sky130_fd_sc_hd__a221o_1
XFILLER_170_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13866_ _14213_/A _14213_/B _13866_/C _13866_/D vssd1 vssd1 vccd1 vccd1 _13867_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_35_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15605_ _15507_/A _15507_/B _15509_/Y vssd1 vssd1 vccd1 vccd1 _15607_/B sky130_fd_sc_hd__a21o_2
XFILLER_37_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12817_ _12817_/A _12817_/B vssd1 vssd1 vccd1 vccd1 _12820_/C sky130_fd_sc_hd__xnor2_2
X_16585_ _16566_/Y _16567_/X _16579_/X _16584_/X vssd1 vssd1 vccd1 vccd1 _16585_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13797_ _14326_/A _14485_/D _13796_/C vssd1 vssd1 vccd1 vccd1 _13798_/B sky130_fd_sc_hd__a21o_1
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15536_ _10716_/A _14785_/X _14806_/X _15535_/Y vssd1 vssd1 vccd1 vccd1 _15536_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12595_/B _13300_/D _13169_/D _12595_/A vssd1 vssd1 vccd1 vccd1 _12751_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15467_ _15454_/X _15467_/B _15467_/C _15467_/D vssd1 vssd1 vccd1 vccd1 _15467_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_129_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12679_ _12679_/A _12679_/B vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__nand2_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17206_ _17436_/Q _17233_/A2 _17204_/X _17205_/X _17428_/B vssd1 vssd1 vccd1 vccd1
+ _17436_/D sky130_fd_sc_hd__o221a_1
X_14418_ _14533_/A _14419_/B vssd1 vssd1 vccd1 vccd1 _14418_/X sky130_fd_sc_hd__or2_1
X_15398_ _15913_/A _15832_/A vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__nor2_4
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17137_ _17167_/A _14829_/X _14828_/Y _14597_/B vssd1 vssd1 vccd1 vccd1 _17137_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14349_ _14350_/A _14350_/B _14350_/C vssd1 vssd1 vccd1 vccd1 _14349_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17068_ _17064_/X _17065_/X _17066_/X _17018_/Y vssd1 vssd1 vccd1 vccd1 _17068_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16019_ _16019_/A vssd1 vssd1 vccd1 vccd1 _17557_/D sky130_fd_sc_hd__inv_2
X_08910_ _08910_/A _08910_/B _08910_/C vssd1 vssd1 vccd1 vccd1 _08910_/Y sky130_fd_sc_hd__nand3_2
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09890_/A _09898_/A _09890_/C vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__or3_1
XFILLER_112_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _12107_/B _12088_/D _11881_/D _12275_/A vssd1 vssd1 vccd1 vccd1 _08841_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_97_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08772_ _09025_/C _11961_/B _08772_/C _08772_/D vssd1 vssd1 vccd1 vccd1 _08804_/A
+ sky130_fd_sc_hd__and4_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ _09328_/A _09451_/A _09328_/C vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__o21ai_4
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _09256_/A _09255_/B _09255_/C vssd1 vssd1 vccd1 vccd1 _09255_/X sky130_fd_sc_hd__and3_2
XFILLER_167_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09186_ _11953_/A _11953_/B _12338_/D _12174_/D vssd1 vssd1 vccd1 vccd1 _09221_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10030_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_68_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11981_ _11982_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__and2b_1
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13720_ _13720_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__xnor2_2
X_10932_ _11124_/C _10932_/B vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__nand2_2
XFILLER_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13651_ _13643_/A _13745_/D _13534_/A _13532_/B vssd1 vssd1 vccd1 vccd1 _13652_/B
+ sky130_fd_sc_hd__a31o_1
X_10863_ _10863_/A _10863_/B _10863_/C vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__or3_4
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12602_ _12603_/B _12603_/A vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__nand2b_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16272_/A _16271_/B _16271_/A vssd1 vssd1 vccd1 vccd1 _16372_/B sky130_fd_sc_hd__o21ba_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A _13582_/B vssd1 vssd1 vccd1 vccd1 _13584_/A sky130_fd_sc_hd__nor2_1
X_10794_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15321_ _15321_/A _15321_/B _15321_/C _15321_/D vssd1 vssd1 vccd1 vccd1 _15321_/X
+ sky130_fd_sc_hd__and4_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12533_ _12534_/B _12534_/A vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__and2b_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _15254_/S _15252_/B vssd1 vssd1 vccd1 vccd1 _15252_/X sky130_fd_sc_hd__or2_4
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12464_ _12464_/A _12662_/A vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__or2_1
XFILLER_173_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14203_ _14202_/A _14202_/B _14202_/C vssd1 vssd1 vccd1 vccd1 _14279_/B sky130_fd_sc_hd__a21oi_2
XFILLER_144_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ _11415_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__nand2_4
X_15183_ _11321_/X _14790_/Y _14798_/Y _16485_/A _15182_/Y vssd1 vssd1 vccd1 vccd1
+ _15188_/A sky130_fd_sc_hd__o311a_1
X_12395_ _12391_/X _12394_/Y _13838_/S vssd1 vssd1 vccd1 vccd1 _14210_/A sky130_fd_sc_hd__mux2_1
XFILLER_181_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _14134_/A _14134_/B _14134_/C vssd1 vssd1 vccd1 vccd1 _14218_/B sky130_fd_sc_hd__nor3_4
XFILLER_141_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11346_ _11343_/A _11312_/Y _11329_/Y _11367_/A vssd1 vssd1 vccd1 vccd1 _11349_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14065_ _14226_/A _14153_/C vssd1 vssd1 vccd1 vccd1 _14066_/B sky130_fd_sc_hd__nand2_2
XFILLER_79_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11277_ _11651_/A _15530_/A vssd1 vssd1 vccd1 vccd1 _11387_/C sky130_fd_sc_hd__and2_2
X_13016_ _17371_/A _13516_/S _11820_/A _13015_/Y _08718_/A vssd1 vssd1 vccd1 vccd1
+ _13016_/X sky130_fd_sc_hd__a311o_1
X_10228_ _10214_/A _10214_/C _10214_/B vssd1 vssd1 vccd1 vccd1 _10228_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10159_ _10053_/A _10053_/B _10053_/C vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14967_ _15617_/A _15530_/A _14967_/C _14967_/D vssd1 vssd1 vccd1 vccd1 _14967_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _16784_/A _16706_/B vssd1 vssd1 vccd1 vccd1 _16709_/A sky130_fd_sc_hd__and2_2
X_13918_ _13918_/A _13918_/B vssd1 vssd1 vccd1 vccd1 _13919_/B sky130_fd_sc_hd__or2_1
X_14898_ _14899_/C vssd1 vssd1 vccd1 vccd1 _14898_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13849_ _13849_/A _13849_/B _13849_/C vssd1 vssd1 vccd1 vccd1 _13851_/A sky130_fd_sc_hd__nor3_1
X_16637_ _16714_/A _16637_/B vssd1 vssd1 vccd1 vccd1 _16638_/B sky130_fd_sc_hd__or2_4
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16568_ _16568_/A _16568_/B vssd1 vssd1 vccd1 vccd1 _16568_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15519_ _15520_/A _15520_/B _15520_/C vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__o21a_1
X_16499_ _16747_/A _16499_/B _16499_/C vssd1 vssd1 vccd1 vccd1 _16609_/B sky130_fd_sc_hd__or3_2
XFILLER_175_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09040_ _09566_/A _09428_/B vssd1 vssd1 vccd1 vccd1 _17081_/B sky130_fd_sc_hd__nand2_8
XFILLER_175_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap121 _08929_/A vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__buf_2
XFILLER_117_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09942_ _09942_/A _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__and3_1
XFILLER_89_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout904 _17478_/Q vssd1 vssd1 vccd1 vccd1 _10559_/B sky130_fd_sc_hd__buf_12
Xfanout915 _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17402_/C1 sky130_fd_sc_hd__buf_4
Xfanout926 fanout927/X vssd1 vssd1 vccd1 vccd1 fanout926/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _10392_/A _14784_/A _10645_/C _10412_/C vssd1 vssd1 vccd1 vccd1 _09876_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout937 input2/X vssd1 vssd1 vccd1 vccd1 fanout937/X sky130_fd_sc_hd__buf_6
XFILLER_135_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _12258_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__nand2_4
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08755_ _08755_/A _08768_/A vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__nor2_4
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09307_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__and2_2
XFILLER_70_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09238_ _09238_/A _09238_/B _09238_/C vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__nor3_1
XFILLER_103_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09178_/B sky130_fd_sc_hd__nand2b_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11200_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _12180_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__nor2_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__xnor2_2
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11062_ _10951_/A _10949_/Y _10857_/Y _10863_/B vssd1 vssd1 vccd1 vccd1 _11065_/C
+ sky130_fd_sc_hd__a211o_4
XFILLER_150_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10013_ _15262_/B _10013_/B vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__nand2_4
X_15870_ _15868_/A _15868_/B _15871_/B vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__o21ba_1
XFILLER_130_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14821_ _16796_/B _16797_/A _16796_/A vssd1 vssd1 vccd1 vccd1 _16865_/A sky130_fd_sc_hd__a21bo_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _14729_/A _14726_/X _14728_/B vssd1 vssd1 vccd1 vccd1 _14752_/Y sky130_fd_sc_hd__o21ai_1
X_17540_ fanout944/X _17540_/D vssd1 vssd1 vccd1 vccd1 _17540_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11964_ _12166_/A _12158_/C _09225_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _11965_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13703_/A _13703_/B vssd1 vssd1 vccd1 vccd1 _13705_/A sky130_fd_sc_hd__nor2_2
XTAP_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17471_ fanout928/X _17544_/Q vssd1 vssd1 vccd1 vccd1 _17471_/Q sky130_fd_sc_hd__dfxtp_1
X_10915_ _10915_/A _10915_/B vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__xnor2_4
X_14683_ _14683_/A _14693_/B vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__and2_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11895_ _11895_/A _12270_/B _12102_/D _12734_/C vssd1 vssd1 vccd1 vccd1 _12138_/A
+ sky130_fd_sc_hd__and4_2
X_13634_ _13635_/A _13741_/A _13635_/C vssd1 vssd1 vccd1 vccd1 _13741_/B sky130_fd_sc_hd__nor3_2
X_16422_ _16422_/A _16422_/B vssd1 vssd1 vccd1 vccd1 _16509_/B sky130_fd_sc_hd__nand2_2
X_10846_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__xnor2_4
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16353_ _16619_/A _15658_/Y _16681_/C _16446_/A vssd1 vssd1 vccd1 vccd1 _16354_/B
+ sky130_fd_sc_hd__o22a_1
X_13565_ _13565_/A _13695_/A vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__nor2_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _10777_/A _10778_/A _10777_/C vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__nor3_2
XFILLER_157_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ _15305_/C _15373_/B _15314_/A vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__a21boi_1
X_12516_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12516_/Y sky130_fd_sc_hd__nand2b_1
X_16284_ _16192_/A _16192_/B _16184_/A vssd1 vssd1 vccd1 vccd1 _16285_/B sky130_fd_sc_hd__a21o_1
XFILLER_160_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13496_ _13496_/A _13496_/B vssd1 vssd1 vccd1 vccd1 _13498_/B sky130_fd_sc_hd__nor2_1
XFILLER_172_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15235_ _15235_/A _15235_/B _15235_/C vssd1 vssd1 vccd1 vccd1 _15235_/Y sky130_fd_sc_hd__nand3_1
XFILLER_126_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12447_ _12907_/A _12595_/C vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__nand2_4
XFILLER_160_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15166_ _15166_/A _15166_/B vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__xnor2_4
X_12378_ _11781_/B _12377_/Y _13005_/A vssd1 vssd1 vccd1 vccd1 _12379_/B sky130_fd_sc_hd__a21oi_2
XFILLER_119_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ _14117_/A _14117_/B vssd1 vssd1 vccd1 vccd1 _14117_/X sky130_fd_sc_hd__xor2_1
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11329_ _11331_/B _11331_/C _11331_/A vssd1 vssd1 vccd1 vccd1 _11329_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_158_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15097_ _15097_/A _15097_/B vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__or2_2
X_14048_ _14150_/A _14048_/B vssd1 vssd1 vccd1 vccd1 _14057_/A sky130_fd_sc_hd__or2_2
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15999_ _16317_/A _16108_/B _16014_/A vssd1 vssd1 vccd1 vccd1 _16001_/A sky130_fd_sc_hd__a21bo_2
XFILLER_36_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09023_ _09023_/A _09023_/B _09555_/C _09647_/B vssd1 vssd1 vccd1 vccd1 _09026_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout701 _14052_/B vssd1 vssd1 vccd1 vccd1 _14213_/D sky130_fd_sc_hd__buf_8
XFILLER_160_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout712 _13088_/B vssd1 vssd1 vccd1 vccd1 _11870_/B sky130_fd_sc_hd__buf_6
X_09925_ _10542_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _09926_/C sky130_fd_sc_hd__and2_1
Xfanout723 _12054_/B vssd1 vssd1 vccd1 vccd1 _10753_/B sky130_fd_sc_hd__buf_8
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout734 _16298_/A vssd1 vssd1 vccd1 vccd1 _13764_/C sky130_fd_sc_hd__buf_6
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout745 fanout757/X vssd1 vssd1 vccd1 vccd1 _12638_/B sky130_fd_sc_hd__buf_8
XFILLER_113_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout756 fanout757/X vssd1 vssd1 vccd1 vccd1 _17119_/A sky130_fd_sc_hd__buf_4
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _10254_/A _10736_/C vssd1 vssd1 vccd1 vccd1 _09856_/Y sky130_fd_sc_hd__nand2_1
Xfanout767 _13434_/C vssd1 vssd1 vccd1 vccd1 _16014_/A sky130_fd_sc_hd__buf_4
XFILLER_100_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout778 _13196_/B vssd1 vssd1 vccd1 vccd1 _15898_/A sky130_fd_sc_hd__buf_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout789 _13321_/D vssd1 vssd1 vccd1 vccd1 _14901_/B sky130_fd_sc_hd__clkbuf_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08807_ _08808_/A _08806_/Y _09025_/C _12158_/C vssd1 vssd1 vccd1 vccd1 _08883_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_58_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__or2_4
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _17614_/Q _08737_/Y _17131_/A vssd1 vssd1 vccd1 vccd1 _17614_/D sky130_fd_sc_hd__mux2_1
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10700_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__nand2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_186_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ _10632_/A _10632_/B _10632_/C _10632_/D vssd1 vssd1 vccd1 vccd1 _10631_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13350_ _13195_/A _13197_/B _13195_/B vssd1 vssd1 vccd1 vccd1 _13357_/A sky130_fd_sc_hd__o21ba_2
XFILLER_155_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10562_ _10671_/A _10671_/B vssd1 vssd1 vccd1 vccd1 _10672_/A sky130_fd_sc_hd__or2_2
XFILLER_10_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _17375_/A _12270_/C _12105_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12303_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13281_ _13950_/A _13895_/C vssd1 vssd1 vccd1 vccd1 _13282_/B sky130_fd_sc_hd__nand2_1
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__nor2_2
X_15020_ _15401_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15020_/X sky130_fd_sc_hd__and2_1
XFILLER_108_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12232_ _17070_/B _12210_/Y _12231_/X vssd1 vssd1 vccd1 vccd1 _17578_/D sky130_fd_sc_hd__o21ai_1
XFILLER_182_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12163_ _12163_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__nor3_1
XFILLER_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11114_ _11114_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _11130_/A sky130_fd_sc_hd__xnor2_4
XFILLER_190_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16971_ _16971_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _16971_/Y sky130_fd_sc_hd__xnor2_1
X_12094_ _12286_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__and2_4
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15922_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _16036_/A sky130_fd_sc_hd__nor2_4
X_11045_ _11032_/A _11029_/B _11025_/Y vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__o21bai_1
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15855_/A sky130_fd_sc_hd__xnor2_4
XFILLER_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14804_ _14803_/A _14803_/B _10799_/Y vssd1 vssd1 vccd1 vccd1 _14805_/C sky130_fd_sc_hd__o21ai_1
XTAP_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15784_ _15784_/A _15784_/B vssd1 vssd1 vccd1 vccd1 _15787_/B sky130_fd_sc_hd__nor2_1
X_12996_ _12996_/A vssd1 vssd1 vccd1 vccd1 _12997_/C sky130_fd_sc_hd__inv_2
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ fanout930/X _17523_/D vssd1 vssd1 vccd1 vccd1 _17523_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11947_ _11917_/X _11918_/Y _12156_/B _11947_/D vssd1 vssd1 vccd1 vccd1 _11947_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14735_ _17164_/A _13628_/B _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14735_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ fanout941/X _17454_/D vssd1 vssd1 vccd1 vccd1 _17454_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _13390_/X _13393_/B _14666_/S vssd1 vssd1 vccd1 vccd1 _14667_/B sky130_fd_sc_hd__mux2_1
XFILLER_178_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11878_ _11878_/A _11878_/B vssd1 vssd1 vccd1 vccd1 _11888_/A sky130_fd_sc_hd__or2_2
X_13617_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13617_/X sky130_fd_sc_hd__and2b_1
X_16405_ _14938_/X _16396_/Y _16398_/X _17169_/A1 _16404_/X vssd1 vssd1 vccd1 vccd1
+ _16405_/X sky130_fd_sc_hd__o221a_1
XFILLER_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10829_ _10829_/A _10829_/B vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__xnor2_4
X_14597_ _14597_/A _14597_/B vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17385_ _17385_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17385_/X sky130_fd_sc_hd__or2_1
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16336_ _16760_/B _16814_/B vssd1 vssd1 vccd1 vccd1 _16337_/B sky130_fd_sc_hd__nand2_2
X_13548_ _13425_/Y _13430_/A _13662_/B _13547_/X vssd1 vssd1 vccd1 vccd1 _13558_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_158_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16267_ _16268_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16267_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13479_ _13479_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_962 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15218_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15220_/B sky130_fd_sc_hd__xor2_4
XFILLER_173_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16198_ _16290_/B _16198_/B vssd1 vssd1 vccd1 vccd1 _16200_/C sky130_fd_sc_hd__nand2b_2
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15149_ _15204_/A _16880_/A _16807_/A _14901_/B _15147_/A vssd1 vssd1 vccd1 vccd1
+ _15149_/X sky130_fd_sc_hd__o41a_1
XFILLER_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09710_ _10254_/B _10738_/D vssd1 vssd1 vccd1 vccd1 _09710_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ _09642_/B _09642_/A vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__and2b_1
XFILLER_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09572_ _09573_/B _09573_/A vssd1 vssd1 vccd1 vccd1 _09581_/B sky130_fd_sc_hd__nand2b_2
XFILLER_82_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1012 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _09007_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _09006_/X sky130_fd_sc_hd__or2_2
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout520 _11260_/C vssd1 vssd1 vccd1 vccd1 _14788_/A sky130_fd_sc_hd__buf_8
Xfanout531 _17515_/Q vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__buf_8
Xfanout542 _12847_/A vssd1 vssd1 vccd1 vccd1 _14356_/S sky130_fd_sc_hd__buf_6
XFILLER_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09908_ _09932_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09909_/C sky130_fd_sc_hd__and2_1
Xfanout553 fanout554/X vssd1 vssd1 vccd1 vccd1 _11377_/B sky130_fd_sc_hd__clkbuf_4
Xfanout564 _10647_/C vssd1 vssd1 vccd1 vccd1 _15711_/A sky130_fd_sc_hd__buf_6
XFILLER_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout575 _12845_/S vssd1 vssd1 vccd1 vccd1 _15254_/S sky130_fd_sc_hd__buf_4
XFILLER_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout586 _14982_/A vssd1 vssd1 vccd1 vccd1 _09928_/C sky130_fd_sc_hd__buf_2
XFILLER_86_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09839_ _10235_/A _10490_/D _17469_/D _09838_/A vssd1 vssd1 vccd1 vccd1 _09839_/Y
+ sky130_fd_sc_hd__a22oi_2
Xfanout597 _11839_/S vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12850_ _14840_/A _12849_/X _12847_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _12850_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _17363_/A _12077_/C _10543_/C vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__a21o_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12938_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__a21o_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _14519_/B _14519_/C _14519_/A vssd1 vssd1 vccd1 vccd1 _14520_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11732_/Y sky130_fd_sc_hd__nor3_4
XFILLER_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14451_/A _14567_/A vssd1 vssd1 vccd1 vccd1 _14454_/A sky130_fd_sc_hd__nor2_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11663_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__and2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13526_/B _13401_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13403_/B sky130_fd_sc_hd__a21o_2
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17170_ _17150_/X _17156_/X _17169_/X _17170_/B1 _17153_/A vssd1 vssd1 vccd1 vccd1
+ _17574_/D sky130_fd_sc_hd__a32oi_4
X_10614_ _10615_/A _10615_/B _10615_/C vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__a21o_4
X_14382_ _14382_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__or2_2
XFILLER_167_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11594_ _11630_/A _15116_/B vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__nand2_2
XFILLER_183_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _11848_/Y _13832_/Y _16120_/X vssd1 vssd1 vccd1 vccd1 _16122_/C sky130_fd_sc_hd__a21oi_1
X_13333_ _14383_/A _13450_/D _13966_/D _16913_/C vssd1 vssd1 vccd1 vccd1 _13337_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10545_ _10546_/A _10544_/Y _10993_/C _10545_/D vssd1 vssd1 vccd1 vccd1 _10655_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_182_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _15964_/A _15964_/B _15962_/Y vssd1 vssd1 vccd1 vccd1 _16075_/A sky130_fd_sc_hd__a21oi_2
XFILLER_109_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13264_ _13264_/A _13264_/B vssd1 vssd1 vccd1 vccd1 _13266_/B sky130_fd_sc_hd__nor2_1
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10476_ _10694_/B _10360_/D _10809_/D _10115_/A vssd1 vssd1 vccd1 vccd1 _10478_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15003_ _15056_/A _15008_/A _15891_/B vssd1 vssd1 vccd1 vccd1 _15003_/X sky130_fd_sc_hd__or3_2
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12215_ _12546_/B _11816_/Y _12214_/Y vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__a21oi_1
X_13195_ _13195_/A _13195_/B vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__nor2_1
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__nand2_1
XFILLER_111_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16954_ _16758_/C _16893_/A _16935_/A _16758_/B vssd1 vssd1 vccd1 vccd1 _16955_/B
+ sky130_fd_sc_hd__o211a_4
X_12077_ _12243_/A _12243_/B _12077_/C _12950_/B vssd1 vssd1 vccd1 vccd1 _12078_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11028_ _11027_/B _17467_/D _11027_/D _10694_/B vssd1 vssd1 vccd1 vccd1 _11029_/B
+ sky130_fd_sc_hd__a22oi_2
X_15905_ _16015_/A _16014_/B _15898_/Y _15904_/X _15897_/X vssd1 vssd1 vccd1 vccd1
+ _15905_/X sky130_fd_sc_hd__o311a_1
X_16885_ _16886_/A _16886_/B vssd1 vssd1 vccd1 vccd1 _16887_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15836_ _15836_/A _15836_/B vssd1 vssd1 vccd1 vccd1 _15837_/B sky130_fd_sc_hd__xnor2_4
XFILLER_65_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ _15866_/B _15767_/B vssd1 vssd1 vccd1 vccd1 _15769_/C sky130_fd_sc_hd__nor2_1
XFILLER_18_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12979_ _12979_/A _12979_/B vssd1 vssd1 vccd1 vccd1 _12981_/B sky130_fd_sc_hd__xnor2_2
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17506_ fanout933/X _17506_/D vssd1 vssd1 vccd1 vccd1 _17506_/Q sky130_fd_sc_hd__dfxtp_4
X_14718_ _14747_/A _14718_/B vssd1 vssd1 vccd1 vccd1 _14719_/C sky130_fd_sc_hd__nand2_1
XFILLER_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _15698_/A _15698_/B vssd1 vssd1 vccd1 vccd1 _15700_/A sky130_fd_sc_hd__nor2_2
XFILLER_178_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17437_ fanout936/X _17437_/D vssd1 vssd1 vccd1 vccd1 _17437_/Q sky130_fd_sc_hd__dfxtp_4
X_14649_ _14649_/A _14649_/B vssd1 vssd1 vccd1 vccd1 _14651_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_16 _17477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_27 _17457_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_38 _14776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17368_ input58/X _17377_/B _17367_/Y _17372_/C1 vssd1 vssd1 vccd1 vccd1 _17512_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_49 _12245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16319_ _16229_/A _16229_/B _16227_/B vssd1 vssd1 vccd1 vccd1 _16321_/B sky130_fd_sc_hd__a21o_1
XFILLER_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17299_ input47/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17299_/X sky130_fd_sc_hd__or3_1
XFILLER_118_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput101 _17459_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_12_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput112 _17440_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09624_ _09624_/A _09624_/B _09624_/C vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__nor3_1
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09555_ _12243_/A _12243_/B _09555_/C _12923_/D vssd1 vssd1 vccd1 vccd1 _09556_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_93_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _09387_/A _09387_/B _09387_/C vssd1 vssd1 vccd1 vccd1 _09486_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_93_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire217 wire217/A vssd1 vssd1 vccd1 vccd1 wire217/X sky130_fd_sc_hd__buf_2
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ _10330_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__nand2_4
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ _10261_/A _10261_/B _10261_/C vssd1 vssd1 vccd1 vccd1 _10262_/C sky130_fd_sc_hd__nand3_4
X_12000_ _09122_/A _09255_/X _11998_/X _11999_/Y vssd1 vssd1 vccd1 vccd1 _12200_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10192_ _10193_/A _10192_/B _10207_/B _10192_/D vssd1 vssd1 vccd1 vccd1 _10193_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout350 _17537_/Q vssd1 vssd1 vccd1 vccd1 _13977_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_143_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout361 _16913_/C vssd1 vssd1 vccd1 vccd1 _14450_/A sky130_fd_sc_hd__buf_4
XFILLER_28_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout372 _17534_/Q vssd1 vssd1 vccd1 vccd1 _13895_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13951_ _13951_/A _13951_/B vssd1 vssd1 vccd1 vccd1 _13954_/C sky130_fd_sc_hd__xnor2_1
Xfanout383 _17532_/Q vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__buf_6
XFILLER_115_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout394 _16644_/C vssd1 vssd1 vccd1 vccd1 _17405_/A sky130_fd_sc_hd__buf_6
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12902_ _12902_/A _12902_/B _12902_/C vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__nand3_2
X_13882_ _13882_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__xnor2_4
X_16670_ _16670_/A _16670_/B _16670_/C vssd1 vssd1 vccd1 vccd1 _16751_/A sky130_fd_sc_hd__nand3_2
XFILLER_35_919 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ _12991_/B _12834_/B _12834_/C vssd1 vssd1 vccd1 vccd1 _12833_/Y sky130_fd_sc_hd__nor3_4
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15621_ _15621_/A _15621_/B vssd1 vssd1 vccd1 vccd1 _15621_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _17038_/C _15552_/B vssd1 vssd1 vccd1 vccd1 _15552_/X sky130_fd_sc_hd__or2_2
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12764_/A _12764_/B _12764_/C vssd1 vssd1 vccd1 vccd1 _12766_/C sky130_fd_sc_hd__and3_2
XFILLER_42_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14441_/B _14443_/B _14441_/A vssd1 vssd1 vccd1 vccd1 _14505_/B sky130_fd_sc_hd__o21ba_1
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ _16295_/A _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16387_/B sky130_fd_sc_hd__and3_2
XFILLER_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15483_ _15484_/A _15567_/A vssd1 vssd1 vccd1 vccd1 _15483_/Y sky130_fd_sc_hd__nand2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12372_/X _12538_/Y _12539_/Y vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__a21o_1
XFILLER_188_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17222_ _17583_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17222_/X sky130_fd_sc_hd__a21o_1
X_14434_ _14492_/A vssd1 vssd1 vccd1 vccd1 _14434_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11646_ _11646_/A _11646_/B _11646_/C vssd1 vssd1 vccd1 vccd1 _15524_/C sky130_fd_sc_hd__and3_2
XFILLER_175_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 i_wb_addr[1] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_2
X_14365_ _14440_/B _14365_/B vssd1 vssd1 vccd1 vccd1 _14400_/A sky130_fd_sc_hd__nor2_1
XFILLER_167_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17153_ _17153_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _17153_/X sky130_fd_sc_hd__and2_1
Xinput25 i_wb_addr[2] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_8
Xinput36 i_wb_data[0] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
X_11577_ _11582_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput47 i_wb_data[1] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_4
X_13316_ _13317_/A _13317_/B _13317_/C vssd1 vssd1 vccd1 vccd1 _13316_/Y sky130_fd_sc_hd__a21oi_4
Xinput58 i_wb_data[2] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_2
X_16104_ _11465_/A _11465_/B _11707_/Y vssd1 vssd1 vccd1 vccd1 _16105_/B sky130_fd_sc_hd__o21ai_4
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17084_ _17085_/A _17085_/B _17085_/C vssd1 vssd1 vccd1 vccd1 _17086_/A sky130_fd_sc_hd__o21ai_2
X_10528_ _10528_/A _10626_/A vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__nor2_4
Xinput69 i_wb_we vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_6
X_14296_ _14297_/A _14297_/B vssd1 vssd1 vccd1 vccd1 _14296_/X sky130_fd_sc_hd__and2b_1
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _16035_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _16036_/B sky130_fd_sc_hd__xor2_4
X_13247_ _13248_/A _13248_/B _13248_/C vssd1 vssd1 vccd1 vccd1 _13249_/C sky130_fd_sc_hd__o21ai_4
X_10459_ _10459_/A _10459_/B _10459_/C vssd1 vssd1 vccd1 vccd1 _10459_/Y sky130_fd_sc_hd__nand3_2
XFILLER_108_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13178_ _13178_/A _13178_/B _13178_/C vssd1 vssd1 vccd1 vccd1 _13312_/B sky130_fd_sc_hd__and3_4
XFILLER_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12129_ _12620_/A _12129_/B vssd1 vssd1 vccd1 vccd1 _12131_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16937_ _16937_/A _16937_/B vssd1 vssd1 vccd1 vccd1 _16943_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16868_ _16868_/A _16868_/B vssd1 vssd1 vccd1 vccd1 _16872_/A sky130_fd_sc_hd__nor2_1
X_15819_ _16127_/A _15726_/D _15817_/X _15726_/A vssd1 vssd1 vccd1 vccd1 _15821_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16799_ _16796_/B _17162_/A2 _16974_/B _14863_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16799_/X sky130_fd_sc_hd__a221o_1
X_09340_ _09391_/B _09391_/C _09391_/A vssd1 vssd1 vccd1 vccd1 _09395_/B sky130_fd_sc_hd__a21oi_4
XFILLER_179_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09271_ _12243_/B _09030_/D _09414_/C _12243_/A vssd1 vssd1 vccd1 vccd1 _09273_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _08985_/A _09074_/A vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__and2b_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09607_/A _09735_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__nor2_4
XFILLER_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09538_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__xor2_2
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ _09473_/A _09591_/A _09473_/C vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__o21ai_4
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _11499_/A _11539_/A _11456_/X _11490_/Y vssd1 vssd1 vccd1 vccd1 _11502_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__and3_1
XFILLER_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11431_ _11430_/A _11475_/A vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__nand2b_4
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14150_ _14150_/A _14150_/B _14150_/C vssd1 vssd1 vccd1 vccd1 _14151_/B sky130_fd_sc_hd__nor3_1
XFILLER_171_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11362_ _11362_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__xnor2_4
XFILLER_193_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _13101_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _13103_/B sky130_fd_sc_hd__xnor2_2
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10313_ _10314_/B _10314_/A vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__and2b_1
XFILLER_180_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14081_ _14081_/A _14173_/A vssd1 vssd1 vccd1 vccd1 _14084_/A sky130_fd_sc_hd__nor2_2
X_11293_ _11293_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _13033_/A _13033_/B _13033_/C vssd1 vssd1 vccd1 vccd1 _13046_/A sky130_fd_sc_hd__a21o_4
XFILLER_79_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10244_ _11026_/A _10911_/B vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__nand2_4
XFILLER_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10175_ _10288_/A _10296_/A _10288_/C vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__o21ai_4
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout180 _15687_/B vssd1 vssd1 vccd1 vccd1 _16747_/A sky130_fd_sc_hd__buf_6
X_14983_ _15095_/B _14981_/Y _14982_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _14983_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout191 _15263_/Y vssd1 vssd1 vccd1 vccd1 _16352_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16722_ _16722_/A _17153_/B vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__nor2_1
X_13934_ _13935_/A _13935_/B vssd1 vssd1 vccd1 vccd1 _13934_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16653_ _16653_/A _16653_/B vssd1 vssd1 vccd1 vccd1 _16653_/X sky130_fd_sc_hd__or2_1
X_13865_ _14213_/B _13866_/C _13764_/C _14213_/A vssd1 vssd1 vccd1 vccd1 _13867_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15604_ _15604_/A _15604_/B vssd1 vssd1 vccd1 vccd1 _15607_/A sky130_fd_sc_hd__xnor2_4
X_12816_ _12816_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__xnor2_2
X_16584_ _17169_/A1 _16577_/X _16583_/X _16569_/X vssd1 vssd1 vccd1 vccd1 _16584_/X
+ sky130_fd_sc_hd__o211a_1
X_13796_ _14326_/A _14485_/D _13796_/C vssd1 vssd1 vccd1 vccd1 _13906_/B sky130_fd_sc_hd__nand3_2
XFILLER_37_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15535_ _16485_/A _15535_/B vssd1 vssd1 vccd1 vccd1 _15535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12747_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__xnor2_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12678_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__o21ai_1
X_15466_ _16115_/A _15541_/B _15463_/Y _15465_/Y _15462_/Y vssd1 vssd1 vccd1 vccd1
+ _15467_/D sky130_fd_sc_hd__o311a_1
XFILLER_147_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ _17545_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__and2_1
X_14417_ _14284_/B _14534_/A _14415_/X vssd1 vssd1 vccd1 vccd1 _14419_/B sky130_fd_sc_hd__a21o_1
XFILLER_128_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ _11629_/A _11629_/B _11629_/C _14794_/B vssd1 vssd1 vccd1 vccd1 _11632_/A
+ sky130_fd_sc_hd__and4_1
X_15397_ _15397_/A _16246_/A vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__nand2_8
XFILLER_156_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17136_ _17099_/Y _17102_/X _17133_/Y _17134_/X vssd1 vssd1 vccd1 vccd1 _17136_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14348_ _14348_/A _14348_/B vssd1 vssd1 vccd1 vccd1 _14350_/C sky130_fd_sc_hd__xnor2_1
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14279_ _14279_/A _14279_/B vssd1 vssd1 vccd1 vccd1 _14279_/Y sky130_fd_sc_hd__nor2_1
X_17067_ _17018_/Y _17066_/X _17065_/X _17064_/X vssd1 vssd1 vccd1 vccd1 _17067_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_143_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16018_ _15996_/Y _15998_/X _16017_/X _14871_/Y _16014_/A vssd1 vssd1 vccd1 vccd1
+ _16019_/A sky130_fd_sc_hd__a32o_1
XFILLER_170_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _12275_/A _12107_/B _12088_/D _11881_/D vssd1 vssd1 vccd1 vccd1 _08843_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08771_ _09023_/B _12166_/B _12158_/C _09023_/A vssd1 vssd1 vccd1 vccd1 _08772_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09328_/C sky130_fd_sc_hd__nor2_2
XFILLER_167_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09254_ _09255_/B _09255_/C vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__nand2_2
XFILLER_166_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ _11953_/B _12338_/D _12174_/D _11953_/A vssd1 vssd1 vccd1 vccd1 _09189_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_181_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08969_ _12845_/S _08969_/B _08969_/C vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__and3_4
XFILLER_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11980_ _11980_/A _11980_/B vssd1 vssd1 vccd1 vccd1 _11982_/B sky130_fd_sc_hd__xnor2_2
XFILLER_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10931_ _14788_/A _11335_/B _10922_/X _14806_/A _10800_/C vssd1 vssd1 vccd1 vccd1
+ _10938_/A sky130_fd_sc_hd__a32o_4
XFILLER_16_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13650_ _13648_/X _13650_/B vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__and2b_1
X_10862_ _10861_/A _10861_/B _10861_/C vssd1 vssd1 vccd1 vccd1 _10863_/C sky130_fd_sc_hd__a21oi_4
XFILLER_182_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12446_/A _12448_/B _12446_/B vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__o21ba_2
X_13581_ _14153_/A _14153_/B _13866_/C _13764_/C vssd1 vssd1 vccd1 vccd1 _13582_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ _11629_/B _10791_/C _10640_/D _11561_/A vssd1 vssd1 vccd1 vccd1 _10794_/B
+ sky130_fd_sc_hd__a22oi_4
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__nand2b_1
X_15320_ _15386_/A _15313_/Y _15319_/X _17164_/C vssd1 vssd1 vccd1 vccd1 _15321_/D
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12463_ _12618_/A _12770_/B _12618_/D _12463_/D vssd1 vssd1 vccd1 vccd1 _12662_/A
+ sky130_fd_sc_hd__and4_1
X_15251_ _16485_/A _15243_/Y _15244_/X _15250_/X vssd1 vssd1 vccd1 vccd1 _15257_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14202_ _14202_/A _14202_/B _14202_/C vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__and3_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _11299_/B _11299_/C _11299_/A vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__o21ai_2
X_15182_ _11321_/X _14790_/Y _14798_/Y vssd1 vssd1 vccd1 vccd1 _15182_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ _12394_/A vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__inv_2
X_14133_ _13947_/Y _14042_/Y _14218_/A vssd1 vssd1 vccd1 vccd1 _14134_/C sky130_fd_sc_hd__a21o_1
XFILLER_152_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11345_ _11345_/A _11345_/B vssd1 vssd1 vccd1 vccd1 _11357_/A sky130_fd_sc_hd__xor2_4
XFILLER_153_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14064_ _14064_/A _14064_/B vssd1 vssd1 vccd1 vccd1 _14066_/A sky130_fd_sc_hd__nor2_1
XFILLER_165_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11276_ _11137_/C _11276_/B vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__and2b_2
XFILLER_141_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _17371_/A _13015_/B vssd1 vssd1 vccd1 vccd1 _13015_/Y sky130_fd_sc_hd__nor2_1
X_10227_ _10219_/A _10219_/C _10219_/B vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__o21ai_4
XFILLER_121_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10158_ _10157_/C _10157_/Y _10028_/B _10104_/X vssd1 vssd1 vccd1 vccd1 _10193_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14966_ _17612_/Q _15208_/C _14877_/Y vssd1 vssd1 vccd1 vccd1 _14966_/X sky130_fd_sc_hd__a21o_1
X_10089_ _10081_/A _10084_/A _10090_/A _10088_/X vssd1 vssd1 vccd1 vccd1 _10101_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_82_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16705_ _16705_/A _16705_/B vssd1 vssd1 vccd1 vccd1 _16706_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _13918_/A _13918_/B vssd1 vssd1 vccd1 vccd1 _14018_/B sky130_fd_sc_hd__nand2_1
X_14897_ _14897_/A _15208_/C _15208_/D _14897_/D vssd1 vssd1 vccd1 vccd1 _14899_/C
+ sky130_fd_sc_hd__or4_4
X_16636_ _16636_/A _16636_/B _16636_/C vssd1 vssd1 vccd1 vccd1 _16637_/B sky130_fd_sc_hd__and3_1
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13848_ _13848_/A _13848_/B vssd1 vssd1 vccd1 vccd1 _13849_/C sky130_fd_sc_hd__xnor2_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16567_ _16566_/A _16566_/B _17063_/A vssd1 vssd1 vccd1 vccd1 _16567_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ _13779_/A _13779_/B vssd1 vssd1 vccd1 vccd1 _13781_/A sky130_fd_sc_hd__nor2_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15518_ _15518_/A _15518_/B vssd1 vssd1 vccd1 vccd1 _15520_/C sky130_fd_sc_hd__xnor2_1
XFILLER_175_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16498_ _16498_/A _16609_/A vssd1 vssd1 vccd1 vccd1 _16499_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15449_ _15532_/A vssd1 vssd1 vccd1 vccd1 _15449_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _17119_/A _17119_/B _17119_/C vssd1 vssd1 vccd1 vccd1 _17121_/A sky130_fd_sc_hd__and3_1
Xmax_cap122 _10500_/Y vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_144_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__nor2_2
XFILLER_143_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout905 _17270_/B1 vssd1 vssd1 vccd1 vccd1 _17231_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_135_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout916 _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17414_/C1 sky130_fd_sc_hd__buf_4
Xfanout927 fanout929/X vssd1 vssd1 vccd1 vccd1 fanout927/X sky130_fd_sc_hd__clkbuf_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__nor2_2
XFILLER_174_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout938 fanout940/X vssd1 vssd1 vccd1 vccd1 fanout938/X sky130_fd_sc_hd__clkbuf_4
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _12088_/A _12088_/B _11867_/C _11867_/D vssd1 vssd1 vccd1 vccd1 _08826_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_100_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _09025_/C _12166_/B _08754_/C _08754_/D vssd1 vssd1 vccd1 vccd1 _08768_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09306_ _09306_/A _09306_/B vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__nor2_1
XFILLER_179_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09237_ _09238_/A _09238_/B _09238_/C vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__o21a_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09168_/A _09168_/B vssd1 vssd1 vccd1 vccd1 _09333_/B sky130_fd_sc_hd__xnor2_4
XFILLER_135_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09099_ _09780_/A _09350_/B _14978_/A vssd1 vssd1 vccd1 vccd1 _09099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _11130_/A _11130_/B _11130_/C vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__nand3_2
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11061_ _11061_/A _11077_/A _11061_/C vssd1 vssd1 vccd1 vccd1 _11065_/B sky130_fd_sc_hd__nand3_4
XFILLER_103_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10012_ _10018_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__nor2_2
XFILLER_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14820_ _16729_/B _16730_/A _13459_/A vssd1 vssd1 vccd1 vccd1 _16797_/A sky130_fd_sc_hd__a21o_1
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14751_/A _14751_/B vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11963_ _12169_/B _11963_/B vssd1 vssd1 vccd1 vccd1 _11966_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13702_/A _13702_/B _13702_/C vssd1 vssd1 vccd1 vccd1 _13703_/B sky130_fd_sc_hd__and3_1
X_17470_ fanout928/X _17543_/Q vssd1 vssd1 vccd1 vccd1 _17470_/Q sky130_fd_sc_hd__dfxtp_1
X_10914_ _10914_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10915_/B sky130_fd_sc_hd__nor2_2
XTAP_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14682_ _14682_/A _14682_/B vssd1 vssd1 vccd1 vccd1 _14719_/A sky130_fd_sc_hd__xnor2_4
X_11894_ _12270_/B _12102_/D _12734_/C _11895_/A vssd1 vssd1 vccd1 vccd1 _11894_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16421_ _16422_/A _16422_/B vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__or2_1
X_13633_ _14775_/A _14002_/B vssd1 vssd1 vccd1 vccd1 _13635_/C sky130_fd_sc_hd__nand2_2
X_10845_ _10846_/A _10846_/B vssd1 vssd1 vccd1 vccd1 _10943_/B sky130_fd_sc_hd__nand2_2
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16352_ _16352_/A _16352_/B _16352_/C vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__and3_1
XFILLER_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13564_ _13895_/A _13895_/B _13564_/C _13564_/D vssd1 vssd1 vccd1 vccd1 _13695_/A
+ sky130_fd_sc_hd__and4_2
X_10776_ _10678_/B _10691_/X _10774_/A _11722_/A vssd1 vssd1 vccd1 vccd1 _10777_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15303_ _15303_/A _15303_/B vssd1 vssd1 vccd1 vccd1 _15303_/Y sky130_fd_sc_hd__nand2_1
X_12515_ _12670_/A _12515_/B vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__nor2_4
X_16283_ _16283_/A _16283_/B vssd1 vssd1 vccd1 vccd1 _16285_/A sky130_fd_sc_hd__xor2_4
XFILLER_158_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13495_ _13495_/A _13495_/B vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__nor2_1
XFILLER_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12446_ _12446_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12448_/A sky130_fd_sc_hd__nor2_2
X_15234_ _15233_/A _15233_/B _14836_/A vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _12377_/A _12377_/B vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__nor2_2
X_15165_ _15165_/A _15230_/A vssd1 vssd1 vccd1 vccd1 _15166_/B sky130_fd_sc_hd__nand2_4
XFILLER_176_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14116_ _14117_/A _14117_/B vssd1 vssd1 vccd1 vccd1 _14202_/B sky130_fd_sc_hd__nand2b_1
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _11369_/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11331_/C sky130_fd_sc_hd__nand2_2
XFILLER_153_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15096_ _14978_/Y _14981_/Y _15096_/S vssd1 vssd1 vccd1 vccd1 _15097_/B sky130_fd_sc_hd__mux2_1
XFILLER_180_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14047_ _14047_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14048_/B sky130_fd_sc_hd__and2_1
X_11259_ _11258_/B _11561_/D _15402_/A _11314_/A vssd1 vssd1 vccd1 vccd1 _11259_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_140_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15998_ _16207_/B _15998_/B _11707_/Y vssd1 vssd1 vccd1 vccd1 _15998_/X sky130_fd_sc_hd__or3b_4
XFILLER_54_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ _14949_/A _14949_/B vssd1 vssd1 vccd1 vccd1 _14949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16619_ _16619_/A _16827_/D _16695_/C vssd1 vssd1 vccd1 vccd1 _16774_/A sky130_fd_sc_hd__or3_4
X_17599_ fanout943/X _17599_/D vssd1 vssd1 vccd1 vccd1 _17599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09924_ _09928_/C _09926_/B _09783_/A _09781_/Y vssd1 vssd1 vccd1 vccd1 _09930_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout702 _16651_/A vssd1 vssd1 vccd1 vccd1 _14052_/B sky130_fd_sc_hd__buf_6
XFILLER_160_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout713 _12077_/C vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout724 _17496_/Q vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__buf_6
Xfanout735 _12068_/C vssd1 vssd1 vccd1 vccd1 _16298_/A sky130_fd_sc_hd__buf_8
Xfanout746 fanout757/X vssd1 vssd1 vccd1 vccd1 _12068_/D sky130_fd_sc_hd__clkbuf_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _10254_/A _10254_/B _10738_/D _10736_/C vssd1 vssd1 vccd1 vccd1 _09855_/X
+ sky130_fd_sc_hd__and4_1
Xfanout757 _17493_/Q vssd1 vssd1 vccd1 vccd1 fanout757/X sky130_fd_sc_hd__buf_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout768 _17492_/Q vssd1 vssd1 vccd1 vccd1 _13434_/C sky130_fd_sc_hd__buf_6
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout779 _17491_/Q vssd1 vssd1 vccd1 vccd1 _13196_/B sky130_fd_sc_hd__buf_12
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _09023_/B _11961_/B _12340_/B _09023_/A vssd1 vssd1 vccd1 vccd1 _08806_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09786_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__or2_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _14929_/A vssd1 vssd1 vccd1 vccd1 _08737_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10630_ _10499_/Y _10589_/X _10598_/X _10611_/Y vssd1 vssd1 vccd1 vccd1 _10632_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10561_ _10561_/A _11749_/A vssd1 vssd1 vccd1 vccd1 _10671_/B sky130_fd_sc_hd__or2_1
XFILLER_182_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12300_ _12508_/B _12300_/B vssd1 vssd1 vccd1 vccd1 _12307_/A sky130_fd_sc_hd__nor2_4
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13280_ _13280_/A _13280_/B vssd1 vssd1 vccd1 vccd1 _13282_/A sky130_fd_sc_hd__nor2_2
XFILLER_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10492_ _11006_/B _10490_/C _10490_/D _11006_/A vssd1 vssd1 vccd1 vccd1 _10493_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _11849_/A _12227_/X _12230_/X _17165_/A1 vssd1 vssd1 vccd1 vccd1 _12231_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12162_ _12162_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12163_/C sky130_fd_sc_hd__nor2_2
XFILLER_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11113_ _11112_/A _11112_/C _11112_/B vssd1 vssd1 vccd1 vccd1 _11113_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_111_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16970_ _16970_/A _16970_/B vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__nand2_1
X_12093_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__or3_1
XFILLER_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15921_ _15921_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15923_/B sky130_fd_sc_hd__xnor2_2
X_11044_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__nand2b_2
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15852_ _15853_/A _15853_/B vssd1 vssd1 vccd1 vccd1 _15852_/Y sky130_fd_sc_hd__nand2_1
XTAP_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14803_ _14803_/A _14803_/B vssd1 vssd1 vccd1 vccd1 _14803_/Y sky130_fd_sc_hd__nor2_1
XTAP_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15783_ _15784_/A _15784_/B vssd1 vssd1 vccd1 vccd1 _15883_/B sky130_fd_sc_hd__and2_2
XFILLER_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _12800_/A _12950_/B _12801_/A _12799_/A vssd1 vssd1 vccd1 vccd1 _12996_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17522_ fanout931/X _17522_/D vssd1 vssd1 vccd1 vccd1 _17522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14734_/A _14734_/B vssd1 vssd1 vccd1 vccd1 _14734_/Y sky130_fd_sc_hd__nand2_1
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11946_ _11943_/Y _11944_/X _09006_/X _09010_/A vssd1 vssd1 vccd1 vccd1 _11947_/D
+ sky130_fd_sc_hd__o211ai_4
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17453_ fanout941/X _17453_/D vssd1 vssd1 vccd1 vccd1 _17453_/Q sky130_fd_sc_hd__dfxtp_2
X_14665_ _14756_/A1 _14663_/Y _14664_/X _14636_/Y _14637_/X vssd1 vssd1 vccd1 vccd1
+ _17602_/D sky130_fd_sc_hd__a32o_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11877_/A _11877_/B _11877_/C vssd1 vssd1 vccd1 vccd1 _11891_/B sky130_fd_sc_hd__and3_2
XFILLER_189_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16404_ _16404_/A _16404_/B _16404_/C vssd1 vssd1 vccd1 vccd1 _16404_/X sky130_fd_sc_hd__and3_1
X_13616_ _13618_/B _13618_/A vssd1 vssd1 vccd1 vccd1 _13616_/Y sky130_fd_sc_hd__nand2b_1
X_10828_ _10828_/A _10828_/B vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__xnor2_4
X_17384_ input37/X _17384_/A2 _17383_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17520_/D
+ sky130_fd_sc_hd__o211a_1
X_14596_ _14676_/A _14641_/C vssd1 vssd1 vccd1 vccd1 _14596_/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16335_ _16333_/X _16335_/B vssd1 vssd1 vccd1 vccd1 _16337_/A sky130_fd_sc_hd__nand2b_1
X_13547_ _13662_/A _13545_/X _13418_/A _13419_/Y vssd1 vssd1 vccd1 vccd1 _13547_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_146_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _11726_/A _10759_/B vssd1 vssd1 vccd1 vccd1 _10760_/C sky130_fd_sc_hd__and2_2
XFILLER_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16266_ _16266_/A _16266_/B vssd1 vssd1 vccd1 vccd1 _16268_/B sky130_fd_sc_hd__xor2_2
X_13478_ _13479_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__or2_2
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15217_ _15218_/A _15218_/B vssd1 vssd1 vccd1 vccd1 _15283_/A sky130_fd_sc_hd__or2_4
XFILLER_126_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12429_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__nor3_2
X_16197_ _16197_/A _16197_/B _16195_/Y vssd1 vssd1 vccd1 vccd1 _16198_/B sky130_fd_sc_hd__or3b_1
XFILLER_127_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15148_ _15262_/C _15270_/B vssd1 vssd1 vccd1 vccd1 _17083_/A sky130_fd_sc_hd__nand2_8
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15079_ _14898_/Y _15077_/Y _11377_/D vssd1 vssd1 vccd1 vccd1 _15734_/B sky130_fd_sc_hd__o21ai_4
XFILLER_113_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09640_ _09640_/A _09795_/A vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09571_ _10255_/A _10791_/C _09570_/B _09567_/Y vssd1 vssd1 vccd1 vccd1 _09573_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_167_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09005_ _08946_/A _08946_/B _08944_/X vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__a21oi_2
XFILLER_152_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout510 _10036_/B vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__buf_4
Xfanout521 _10640_/C vssd1 vssd1 vccd1 vccd1 _11260_/C sky130_fd_sc_hd__clkbuf_16
Xfanout532 _10419_/A vssd1 vssd1 vccd1 vccd1 _14789_/A sky130_fd_sc_hd__buf_6
X_09907_ _09784_/A _09784_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09908_/B sky130_fd_sc_hd__o21ai_1
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout543 _12847_/A vssd1 vssd1 vccd1 vccd1 _14839_/A sky130_fd_sc_hd__buf_2
XFILLER_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout554 _17514_/Q vssd1 vssd1 vccd1 vccd1 fanout554/X sky130_fd_sc_hd__buf_6
Xfanout565 _10299_/C vssd1 vssd1 vccd1 vccd1 _10647_/C sky130_fd_sc_hd__buf_6
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout576 _17164_/B vssd1 vssd1 vccd1 vccd1 _12845_/S sky130_fd_sc_hd__buf_6
XFILLER_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _09838_/A _10235_/A _10490_/D _17469_/D vssd1 vssd1 vccd1 vccd1 _09841_/A
+ sky130_fd_sc_hd__and4_2
Xfanout587 _12398_/S vssd1 vssd1 vccd1 vccd1 _14982_/A sky130_fd_sc_hd__clkbuf_8
Xfanout598 _11839_/S vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09769_ _09769_/A _09769_/B _09776_/B _09769_/D vssd1 vssd1 vccd1 vccd1 _09812_/C
+ sky130_fd_sc_hd__and4_2
XFILLER_6_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11800_ _14888_/A _14876_/C _11800_/C _11800_/D vssd1 vssd1 vccd1 vccd1 _11800_/Y
+ sky130_fd_sc_hd__nor4_4
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12780_ _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12782_/C sky130_fd_sc_hd__xnor2_4
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11731_/A _11731_/B _11736_/A vssd1 vssd1 vccd1 vccd1 _11732_/C sky130_fd_sc_hd__nor3_4
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14450_ _14450_/A _14708_/C _14509_/A vssd1 vssd1 vccd1 vccd1 _14567_/A sky130_fd_sc_hd__and3_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A _11662_/B vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__xnor2_1
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _13526_/B _13401_/B _13401_/C vssd1 vssd1 vccd1 vccd1 _13403_/A sky130_fd_sc_hd__nand3_1
X_10613_ _10613_/A _10613_/B vssd1 vssd1 vccd1 vccd1 _10615_/C sky130_fd_sc_hd__xnor2_2
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14381_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__nor2_1
X_11593_ _11595_/A _14796_/A vssd1 vssd1 vccd1 vccd1 _11593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_128_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16120_ _16108_/C _17119_/A _17075_/A2 _16119_/X vssd1 vssd1 vccd1 vccd1 _16120_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_183_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13332_ _13332_/A _13332_/B _13332_/C vssd1 vssd1 vccd1 vccd1 _13373_/B sky130_fd_sc_hd__and3_2
X_10544_ _15126_/A _10753_/B _10309_/C vssd1 vssd1 vccd1 vccd1 _10544_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16051_ _16051_/A _16051_/B vssd1 vssd1 vccd1 vccd1 _16077_/A sky130_fd_sc_hd__xnor2_1
X_10475_ _10385_/A _10385_/C _10385_/B vssd1 vssd1 vccd1 vccd1 _10475_/Y sky130_fd_sc_hd__a21oi_2
X_13263_ _13263_/A _13263_/B vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__nand2_1
XFILLER_182_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15002_ _14794_/A _15373_/B _11675_/B vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__a21o_1
X_12214_ _12214_/A _12546_/C vssd1 vssd1 vccd1 vccd1 _12214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_170_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ _17425_/A _17423_/A _13321_/D _13194_/D vssd1 vssd1 vccd1 vccd1 _13195_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12145_ _12145_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__or2_1
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16953_ _16953_/A _16953_/B vssd1 vssd1 vccd1 vccd1 _16955_/A sky130_fd_sc_hd__nor2_4
X_12076_ _11867_/B _12077_/C _12950_/B _09030_/A vssd1 vssd1 vccd1 vccd1 _12078_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11027_ _11027_/A _11027_/B _11027_/C _11027_/D vssd1 vssd1 vccd1 vccd1 _11032_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15904_ _14924_/A _12401_/A _13516_/X _15900_/Y _15903_/X vssd1 vssd1 vccd1 vccd1
+ _15904_/X sky130_fd_sc_hd__o311a_1
X_16884_ _16939_/B _16884_/B vssd1 vssd1 vccd1 vccd1 _16886_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15835_ _15836_/B _15836_/A vssd1 vssd1 vccd1 vccd1 _15966_/B sky130_fd_sc_hd__nand2b_1
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15868_/B _15765_/C _15765_/A vssd1 vssd1 vccd1 vccd1 _15767_/B sky130_fd_sc_hd__o21a_1
XFILLER_45_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _12978_/A _12978_/B vssd1 vssd1 vccd1 vccd1 _12979_/B sky130_fd_sc_hd__and2_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17505_ fanout933/X _17505_/D vssd1 vssd1 vccd1 vccd1 _17505_/Q sky130_fd_sc_hd__dfxtp_4
X_14717_ _14717_/A _14717_/B vssd1 vssd1 vccd1 vccd1 _14718_/B sky130_fd_sc_hd__nand2_1
X_11929_ _11930_/B _12752_/B _12270_/C _17373_/A vssd1 vssd1 vccd1 vccd1 _11931_/A
+ sky130_fd_sc_hd__a22oi_2
X_15697_ _15786_/B _15695_/X _15603_/Y _15606_/Y vssd1 vssd1 vccd1 vccd1 _15698_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17436_ fanout936/X _17436_/D vssd1 vssd1 vccd1 vccd1 _17436_/Q sky130_fd_sc_hd__dfxtp_4
X_14648_ _14680_/A _14708_/C _14679_/B vssd1 vssd1 vccd1 vccd1 _14649_/B sky130_fd_sc_hd__and3_2
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_17 _17473_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _17464_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_39 _11027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _17367_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17367_/Y sky130_fd_sc_hd__nand2_1
X_14579_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _14580_/B sky130_fd_sc_hd__and2_1
XFILLER_119_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16318_ _16318_/A _16504_/B vssd1 vssd1 vccd1 vccd1 _16321_/A sky130_fd_sc_hd__xnor2_1
XFILLER_186_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17298_ _10560_/D _17322_/A2 _17297_/X _17428_/B vssd1 vssd1 vccd1 vccd1 _17478_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16249_ _16250_/A _16250_/B _16250_/C vssd1 vssd1 vccd1 vccd1 _16251_/A sky130_fd_sc_hd__o21a_2
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 _17460_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[26] sky130_fd_sc_hd__clkbuf_2
Xoutput113 _17441_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09623_ _09616_/Y _09621_/X _09629_/A _09601_/Y vssd1 vssd1 vccd1 vccd1 _09629_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _12243_/B _10839_/D _12338_/C _12243_/A vssd1 vssd1 vccd1 vccd1 _09556_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09485_ _09458_/X _09628_/A _09391_/C _09399_/Y vssd1 vssd1 vccd1 vccd1 _09485_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10260_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10262_/B sky130_fd_sc_hd__xnor2_4
XFILLER_106_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ _10028_/B _10104_/X _10157_/C _10157_/Y vssd1 vssd1 vccd1 vccd1 _10192_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout340 _14599_/A vssd1 vssd1 vccd1 vccd1 _14153_/A sky130_fd_sc_hd__buf_6
XFILLER_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout351 _12176_/A vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__buf_4
Xfanout362 _17413_/A vssd1 vssd1 vccd1 vccd1 _16913_/C sky130_fd_sc_hd__buf_8
X_13950_ _13950_/A _14181_/B vssd1 vssd1 vccd1 vccd1 _13951_/B sky130_fd_sc_hd__nand2_2
Xfanout373 _10321_/A vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__clkbuf_4
Xfanout384 _14248_/A vssd1 vssd1 vccd1 vccd1 _14326_/A sky130_fd_sc_hd__buf_6
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout395 _17531_/Q vssd1 vssd1 vccd1 vccd1 _16644_/C sky130_fd_sc_hd__buf_6
X_12901_ _12902_/A _12902_/B _12902_/C vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__a21o_2
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13881_ _13882_/A _13882_/B vssd1 vssd1 vccd1 vccd1 _13986_/A sky130_fd_sc_hd__and2b_1
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15620_ _15620_/A _15620_/B vssd1 vssd1 vccd1 vccd1 _15621_/B sky130_fd_sc_hd__and2_1
X_12832_ _12685_/A _12685_/B _12681_/Y vssd1 vssd1 vccd1 vccd1 _12834_/C sky130_fd_sc_hd__o21ba_2
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_931 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15551_/A _15552_/B vssd1 vssd1 vccd1 vccd1 _15551_/Y sky130_fd_sc_hd__nor2_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12764_/A _12764_/B _12764_/C vssd1 vssd1 vccd1 vccd1 _12928_/B sky130_fd_sc_hd__a21oi_4
XFILLER_188_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14502_ _14502_/A _14562_/B vssd1 vssd1 vccd1 vccd1 _14505_/A sky130_fd_sc_hd__nand2_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16294_/B sky130_fd_sc_hd__and2_1
X_15482_ _14898_/Y _15077_/Y _16533_/A _11377_/D vssd1 vssd1 vccd1 vccd1 _15567_/A
+ sky130_fd_sc_hd__o211a_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12694_/A _12694_/B vssd1 vssd1 vccd1 vccd1 _13003_/A sky130_fd_sc_hd__xnor2_2
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _17441_/Q _17233_/A2 _17219_/X _17220_/X _17372_/C1 vssd1 vssd1 vccd1 vccd1
+ _17441_/D sky130_fd_sc_hd__o221a_1
X_14433_ _14680_/A _14593_/C vssd1 vssd1 vccd1 vccd1 _14492_/A sky130_fd_sc_hd__nand2_8
X_11645_ _11641_/A _11664_/A _11644_/X vssd1 vssd1 vccd1 vccd1 _11646_/C sky130_fd_sc_hd__a21o_1
XFILLER_174_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ _17153_/B _17167_/C vssd1 vssd1 vccd1 vccd1 _17152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14364_ _14364_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _14365_/B sky130_fd_sc_hd__and2_1
XFILLER_155_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput15 i_wb_addr[20] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
Xinput26 i_wb_addr[30] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_2
X_11576_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__and2_1
XFILLER_183_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput37 i_wb_data[10] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
X_16103_ _16100_/B _16101_/Y _16102_/X vssd1 vssd1 vccd1 vccd1 _16103_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 i_wb_data[20] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13315_ _13442_/A _13315_/B vssd1 vssd1 vccd1 vccd1 _13317_/C sky130_fd_sc_hd__and2_2
Xinput59 i_wb_data[30] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10527_ _10528_/A _10526_/Y _10970_/A _10743_/C vssd1 vssd1 vccd1 vccd1 _10626_/A
+ sky130_fd_sc_hd__and4bb_2
X_17083_ _17083_/A _17083_/B _17083_/C vssd1 vssd1 vccd1 vccd1 _17085_/C sky130_fd_sc_hd__and3_2
X_14295_ _14372_/B _14295_/B vssd1 vssd1 vccd1 vccd1 _14297_/B sky130_fd_sc_hd__nor2_4
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16034_ _16034_/A _16034_/B vssd1 vssd1 vccd1 vccd1 _16035_/B sky130_fd_sc_hd__xnor2_4
X_10458_ _10459_/A _10459_/B _10459_/C vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__and3_2
X_13246_ _13246_/A _13246_/B vssd1 vssd1 vccd1 vccd1 _13248_/C sky130_fd_sc_hd__and2_1
XFILLER_182_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13177_ _13178_/A _13178_/B _13178_/C vssd1 vssd1 vccd1 vccd1 _13177_/Y sky130_fd_sc_hd__a21oi_4
X_10389_ _10390_/A _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__a21o_4
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12128_ _12128_/A _12343_/A vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__or2_1
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16936_ _16935_/A _16935_/B _16935_/C vssd1 vssd1 vccd1 vccd1 _16937_/B sky130_fd_sc_hd__a21oi_1
X_12059_ _14942_/A _15553_/A _14911_/B vssd1 vssd1 vccd1 vccd1 _12397_/B sky130_fd_sc_hd__or3b_2
XFILLER_38_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16867_ _14864_/A _14864_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _16868_/B sky130_fd_sc_hd__o21ai_1
X_15818_ _16809_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16030_/B sky130_fd_sc_hd__nand2_2
XFILLER_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16798_ _14863_/B _16652_/B _14863_/A vssd1 vssd1 vccd1 vccd1 _16798_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15749_ _15749_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _15751_/B sky130_fd_sc_hd__nand2_2
XFILLER_178_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09270_ _12245_/A _12637_/D vssd1 vssd1 vccd1 vccd1 _16982_/A sky130_fd_sc_hd__nand2_8
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17419_ _17419_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17419_/X sky130_fd_sc_hd__or2_1
XFILLER_193_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08985_ _08985_/A _08985_/B _08985_/C vssd1 vssd1 vccd1 vccd1 _09074_/A sky130_fd_sc_hd__or3_2
XFILLER_180_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09606_ _09607_/A _09605_/Y _09750_/C _10308_/B vssd1 vssd1 vccd1 vccd1 _09735_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09537_ _12800_/A _09414_/C _09213_/B _09212_/A vssd1 vssd1 vccd1 vccd1 _09538_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ _09468_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09473_/C sky130_fd_sc_hd__nor2_2
XFILLER_184_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09399_ _09339_/A _09344_/B _09339_/C vssd1 vssd1 vccd1 vccd1 _09399_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11430_ _11430_/A _11430_/B _11430_/C vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__or3_4
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11361_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__nand2_4
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10312_ _10312_/A _10429_/A vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__nor2_4
X_13100_ _17415_/A _13100_/B vssd1 vssd1 vccd1 vccd1 _13101_/B sky130_fd_sc_hd__nand2_2
XFILLER_164_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14080_ _14318_/B _14545_/D _14080_/C vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__and3_2
X_11292_ _11293_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__or2_4
X_13031_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13033_/C sky130_fd_sc_hd__xnor2_4
X_10243_ _10243_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__nor2_2
XFILLER_180_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10174_ _10174_/A _10174_/B vssd1 vssd1 vccd1 vccd1 _10288_/C sky130_fd_sc_hd__xnor2_2
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14982_ _14982_/A _14982_/B _14982_/C vssd1 vssd1 vccd1 vccd1 _14982_/Y sky130_fd_sc_hd__nor3_1
Xfanout170 _15820_/C vssd1 vssd1 vccd1 vccd1 _16662_/C sky130_fd_sc_hd__buf_4
Xfanout181 _15581_/B vssd1 vssd1 vccd1 vccd1 _16589_/B sky130_fd_sc_hd__buf_6
X_16721_ _16791_/A vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__inv_2
Xfanout192 _15932_/B vssd1 vssd1 vccd1 vccd1 _16410_/A sky130_fd_sc_hd__buf_12
X_13933_ _13936_/A _13936_/B vssd1 vssd1 vccd1 vccd1 _13935_/B sky130_fd_sc_hd__or2_1
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16652_ _16652_/A _16652_/B _16652_/C vssd1 vssd1 vccd1 vccd1 _16652_/X sky130_fd_sc_hd__or3_1
X_13864_ _13862_/X _13864_/B vssd1 vssd1 vccd1 vccd1 _13870_/A sky130_fd_sc_hd__nand2b_1
XFILLER_62_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15603_ _15604_/B _15604_/A vssd1 vssd1 vccd1 vccd1 _15603_/Y sky130_fd_sc_hd__nand2b_2
X_12815_ _12816_/A _12816_/B vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_76_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16583_ _16583_/A1 _14209_/X _16581_/Y _16582_/X vssd1 vssd1 vccd1 vccd1 _16583_/X
+ sky130_fd_sc_hd__o211a_1
X_13795_ _13795_/A _13906_/A vssd1 vssd1 vccd1 vccd1 _13796_/C sky130_fd_sc_hd__and2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _10716_/A _14785_/X _14806_/X vssd1 vssd1 vccd1 vccd1 _15535_/B sky130_fd_sc_hd__a21o_1
XFILLER_163_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12746_ _12747_/A _12747_/B vssd1 vssd1 vccd1 vccd1 _12920_/A sky130_fd_sc_hd__nand2_2
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15465_ _14806_/A _15804_/A2 _15464_/X vssd1 vssd1 vccd1 vccd1 _15465_/Y sky130_fd_sc_hd__a21oi_1
X_12677_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12677_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17204_ _17577_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__a21o_1
X_14416_ _14283_/B _14416_/B vssd1 vssd1 vccd1 vccd1 _14534_/A sky130_fd_sc_hd__and2b_1
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11628_ _11628_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__xnor2_4
XFILLER_191_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15396_ _15396_/A _15396_/B _15472_/B vssd1 vssd1 vccd1 vccd1 _16041_/B sky130_fd_sc_hd__nand3_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17135_ _17133_/Y _17134_/X _17099_/Y _17102_/X vssd1 vssd1 vccd1 vccd1 _17135_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_190_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14347_ _14348_/B _14348_/A vssd1 vssd1 vccd1 vccd1 _14413_/B sky130_fd_sc_hd__and2b_1
XFILLER_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _11520_/C _11561_/C _11521_/A _11519_/Y vssd1 vssd1 vccd1 vccd1 _11565_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_156_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17066_ _17066_/A _17066_/B vssd1 vssd1 vccd1 vccd1 _17066_/X sky130_fd_sc_hd__and2_2
X_14278_ _14278_/A _14278_/B vssd1 vssd1 vccd1 vccd1 _14281_/B sky130_fd_sc_hd__nor2_1
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16017_ _16017_/A _16017_/B _16017_/C vssd1 vssd1 vccd1 vccd1 _16017_/X sky130_fd_sc_hd__and3_1
X_13229_ _17415_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _13230_/B sky130_fd_sc_hd__nand2_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08770_ _08773_/A vssd1 vssd1 vccd1 vccd1 _08772_/C sky130_fd_sc_hd__inv_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16919_ _16918_/A _16918_/B _16918_/C vssd1 vssd1 vccd1 vccd1 _16919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _15538_/A _09652_/B _09317_/A _09086_/Y vssd1 vssd1 vccd1 vccd1 _09323_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09253_ _09250_/Y _09251_/X _09182_/Y _09342_/A vssd1 vssd1 vccd1 vccd1 _09255_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_178_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09184_ _12800_/A _09414_/C vssd1 vssd1 vccd1 vccd1 _09213_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_923 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08968_ _10542_/A _08968_/B vssd1 vssd1 vccd1 vccd1 _08969_/C sky130_fd_sc_hd__and2_4
XFILLER_75_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08899_ _12088_/B _11867_/D _12645_/B _12088_/A vssd1 vssd1 vccd1 vccd1 _08900_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10930_ _11124_/C _11132_/C _10842_/B _10841_/A vssd1 vssd1 vccd1 vccd1 _10940_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _10861_/A _10861_/B _10861_/C vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__and3_4
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12600_/A _12755_/B vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__nor2_4
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _14153_/B _13866_/C _13764_/C _14153_/A vssd1 vssd1 vccd1 vccd1 _13582_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10792_ _10899_/C _10932_/B vssd1 vssd1 vccd1 vccd1 _10884_/A sky130_fd_sc_hd__nand2_2
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12531_ _12526_/B _12361_/B _12361_/C _12366_/A vssd1 vssd1 vccd1 vccd1 _12534_/B
+ sky130_fd_sc_hd__a31o_4
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ _15244_/A _15804_/A2 _15249_/X _14944_/A vssd1 vssd1 vccd1 vccd1 _15250_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _12770_/B _12618_/D _12463_/D _12618_/A vssd1 vssd1 vccd1 vccd1 _12464_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_166_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14201_ _14276_/B _14201_/B vssd1 vssd1 vccd1 vccd1 _14202_/C sky130_fd_sc_hd__nand2b_1
XFILLER_138_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11413_ _11416_/B _11413_/B _11413_/C vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__nor3_4
XFILLER_138_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15181_ _12858_/Y _15180_/B _15179_/X _13837_/A vssd1 vssd1 vccd1 vccd1 _16582_/B
+ sky130_fd_sc_hd__o22a_2
X_12393_ _12865_/S _12393_/B vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__nor2_2
X_14132_ _13951_/B _14042_/Y _13947_/Y vssd1 vssd1 vccd1 vccd1 _14218_/A sky130_fd_sc_hd__a21oi_4
XFILLER_181_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11344_ _11352_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__or2_1
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ _14153_/A _14153_/B _14063_/C _14213_/C vssd1 vssd1 vccd1 vccd1 _14064_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_180_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11275_ _11520_/C _15703_/A _11135_/C vssd1 vssd1 vccd1 vccd1 _11276_/B sky130_fd_sc_hd__a21o_1
XFILLER_106_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13014_ _11805_/X _11810_/X _11838_/X _11843_/X _15384_/S _15538_/A vssd1 vssd1 vccd1
+ vccd1 _13015_/B sky130_fd_sc_hd__mux4_2
X_10226_ _10226_/A _10226_/B vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__xnor2_4
XFILLER_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10157_ _10155_/Y _10157_/B _10157_/C vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _09959_/X _09972_/Y _10060_/Y _10216_/A vssd1 vssd1 vccd1 vccd1 _10088_/X
+ sky130_fd_sc_hd__o211a_2
X_14965_ _15553_/A _16977_/A _14910_/X _14964_/Y vssd1 vssd1 vccd1 vccd1 _17543_/D
+ sky130_fd_sc_hd__o22a_1
X_16704_ _16705_/A _16705_/B vssd1 vssd1 vccd1 vccd1 _16784_/A sky130_fd_sc_hd__or2_1
X_13916_ _14021_/A _13916_/B vssd1 vssd1 vccd1 vccd1 _13918_/B sky130_fd_sc_hd__nor2_1
X_14896_ _15530_/A _14896_/B _15143_/A vssd1 vssd1 vccd1 vccd1 _14897_/D sky130_fd_sc_hd__or3b_1
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16635_ _16636_/A _16636_/B _16636_/C vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__a21oi_2
X_13847_ _13950_/A _13948_/D _13848_/A vssd1 vssd1 vccd1 vccd1 _13954_/B sky130_fd_sc_hd__and3_1
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16566_ _16566_/A _16566_/B vssd1 vssd1 vccd1 vccd1 _16566_/Y sky130_fd_sc_hd__nor2_2
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13778_ _13778_/A _13778_/B _13778_/C vssd1 vssd1 vccd1 vccd1 _13779_/B sky130_fd_sc_hd__nor3_1
XFILLER_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15517_ _15518_/B _15518_/A vssd1 vssd1 vccd1 vccd1 _15609_/B sky130_fd_sc_hd__and2b_1
XFILLER_176_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12729_ _12730_/A _12730_/B _12730_/C vssd1 vssd1 vccd1 vccd1 _12902_/A sky130_fd_sc_hd__a21o_2
X_16497_ _16667_/A _16814_/A _16662_/C _16662_/D vssd1 vssd1 vccd1 vccd1 _16609_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15448_ _15396_/A _15373_/B _15450_/A vssd1 vssd1 vccd1 vccd1 _15532_/A sky130_fd_sc_hd__a21bo_2
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15379_ _10799_/Y _14803_/Y _16304_/A _15378_/X vssd1 vssd1 vccd1 vccd1 _15379_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17118_ _17118_/A _17118_/B vssd1 vssd1 vccd1 vccd1 _17127_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17049_ _17049_/A _17049_/B vssd1 vssd1 vccd1 vccd1 _17050_/B sky130_fd_sc_hd__nor2_1
X_09940_ _10062_/A _10067_/B _09801_/B _09798_/Y vssd1 vssd1 vccd1 vccd1 _09941_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap189 _16505_/A vssd1 vssd1 vccd1 vccd1 _15667_/B sky130_fd_sc_hd__buf_6
Xfanout906 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17291_/B1 sky130_fd_sc_hd__buf_4
XFILLER_131_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _11902_/A _09892_/D _09731_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _09872_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_48_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout917 _17322_/C1 vssd1 vssd1 vccd1 vccd1 _17406_/C1 sky130_fd_sc_hd__buf_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout928 fanout929/X vssd1 vssd1 vccd1 vccd1 fanout928/X sky130_fd_sc_hd__buf_6
XFILLER_98_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout939 fanout944/X vssd1 vssd1 vccd1 vccd1 fanout939/X sky130_fd_sc_hd__clkbuf_4
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08822_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__xnor2_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08753_ _09023_/B _12171_/B _11961_/B _09023_/A vssd1 vssd1 vccd1 vccd1 _08754_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09305_ _09750_/C _10180_/B _09081_/A _09079_/Y vssd1 vssd1 vccd1 vccd1 _09306_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09236_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09238_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _09167_/A _09167_/B vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__or2_4
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09098_ _09926_/A _17139_/A _14981_/A vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__and3_2
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11060_ _11051_/A _11051_/C _11051_/B vssd1 vssd1 vccd1 vccd1 _11061_/C sky130_fd_sc_hd__a21o_2
XFILLER_122_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10011_ _10508_/C _10036_/D _09876_/A _09874_/Y vssd1 vssd1 vccd1 vccd1 _10018_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14750_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14751_/B sky130_fd_sc_hd__nand2_1
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11962_ _12166_/A _11961_/B _11961_/C vssd1 vssd1 vccd1 vccd1 _11963_/B sky130_fd_sc_hd__a21o_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13701_ _13702_/A _13702_/B _13702_/C vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__a21oi_2
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10913_ _10963_/B _10912_/C _11005_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _10914_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_189_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14682_/A _14682_/B vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _11890_/X _11891_/Y _08801_/A _08801_/Y vssd1 vssd1 vccd1 vccd1 _11915_/B
+ sky130_fd_sc_hd__o211a_1
X_16420_ _16420_/A vssd1 vssd1 vccd1 vccd1 _16422_/B sky130_fd_sc_hd__inv_2
X_13632_ _13844_/A _13844_/B _14089_/B _13903_/B vssd1 vssd1 vccd1 vccd1 _13741_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10846_/B sky130_fd_sc_hd__xnor2_4
XFILLER_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _16619_/A _16681_/C vssd1 vssd1 vccd1 vccd1 _16352_/C sky130_fd_sc_hd__nor2_2
X_13563_ _14383_/A _13564_/C _13564_/D _13895_/A vssd1 vssd1 vccd1 vccd1 _13565_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10775_ _10774_/A _11722_/A _10678_/B _10691_/X vssd1 vssd1 vccd1 vccd1 _10778_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15302_ _15302_/A _15302_/B vssd1 vssd1 vccd1 vccd1 _15303_/B sky130_fd_sc_hd__or2_1
X_12514_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12515_/B sky130_fd_sc_hd__and2_1
X_16282_ _16282_/A _16282_/B vssd1 vssd1 vccd1 vccd1 _16283_/B sky130_fd_sc_hd__xor2_4
XFILLER_160_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ _13494_/A _13494_/B _13494_/C vssd1 vssd1 vccd1 vccd1 _13495_/B sky130_fd_sc_hd__nor3_1
XFILLER_173_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/X sky130_fd_sc_hd__or2_2
X_12445_ _17385_/A _17383_/A _12736_/B _12578_/B vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15164_ _15774_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__nand2_2
X_12376_ _12015_/Y _12377_/B _12375_/Y _12208_/B vssd1 vssd1 vccd1 vccd1 _13005_/A
+ sky130_fd_sc_hd__o22ai_4
XFILLER_181_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14115_ _14115_/A _14115_/B vssd1 vssd1 vccd1 vccd1 _14117_/B sky130_fd_sc_hd__nand2_1
XFILLER_154_997 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11327_ _11331_/B _11327_/B vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__and2_2
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15095_ _15097_/A _15095_/B _14979_/B vssd1 vssd1 vccd1 vccd1 _17164_/D sky130_fd_sc_hd__or3b_4
XFILLER_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _14047_/A _14047_/B vssd1 vssd1 vccd1 vccd1 _14150_/A sky130_fd_sc_hd__nor2_1
X_11258_ _11314_/A _11258_/B _11561_/D _15402_/A vssd1 vssd1 vccd1 vccd1 _11261_/A
+ sky130_fd_sc_hd__and4_2
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10210_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11189_ _11218_/B _11187_/X _11053_/Y _11055_/X vssd1 vssd1 vccd1 vccd1 _11190_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15997_ _15997_/A _15997_/B vssd1 vssd1 vccd1 vccd1 _15998_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14948_ _15096_/S _14948_/B _14948_/C vssd1 vssd1 vccd1 vccd1 _14948_/Y sky130_fd_sc_hd__nor3_1
XFILLER_75_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14879_ _15147_/C _17614_/Q vssd1 vssd1 vccd1 vccd1 _14879_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16618_ _16695_/A _16533_/B _16695_/B _16533_/A vssd1 vssd1 vccd1 vccd1 _16620_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17598_ fanout943/X _17598_/D vssd1 vssd1 vccd1 vccd1 _17598_/Q sky130_fd_sc_hd__dfxtp_1
X_16549_ _16550_/A _16550_/B _16550_/C vssd1 vssd1 vccd1 vccd1 _16636_/A sky130_fd_sc_hd__a21o_1
XFILLER_176_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09021_ _09025_/C _09555_/C _08882_/A _08880_/Y vssd1 vssd1 vccd1 vccd1 _09027_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09956_/A sky130_fd_sc_hd__and2_1
Xfanout703 _17499_/Q vssd1 vssd1 vccd1 vccd1 _16651_/A sky130_fd_sc_hd__buf_8
Xfanout714 _10545_/D vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout725 _16399_/A vssd1 vssd1 vccd1 vccd1 _13966_/D sky130_fd_sc_hd__buf_8
Xfanout736 _17495_/Q vssd1 vssd1 vccd1 vccd1 _12068_/C sky130_fd_sc_hd__buf_6
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__xnor2_4
Xfanout747 fanout757/X vssd1 vssd1 vccd1 vccd1 _13664_/D sky130_fd_sc_hd__buf_6
XFILLER_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout758 _17492_/Q vssd1 vssd1 vccd1 vccd1 _12171_/B sky130_fd_sc_hd__buf_12
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout769 _12637_/D vssd1 vssd1 vccd1 vccd1 _12166_/B sky130_fd_sc_hd__buf_6
XFILLER_140_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08805_ _09023_/A _09023_/B _11961_/B _12340_/B vssd1 vssd1 vccd1 vccd1 _08808_/A
+ sky130_fd_sc_hd__and4_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09785_ _09502_/A _10321_/C _17466_/D _09172_/A vssd1 vssd1 vccd1 vccd1 _09786_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _17607_/Q _17608_/Q vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__nand2_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10560_ _10560_/A _10560_/B _11370_/C _10560_/D vssd1 vssd1 vccd1 vccd1 _11749_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_167_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _09219_/A _11958_/A _09219_/C vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__nor3_2
XFILLER_148_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10491_ _11005_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12230_ _15457_/B _12230_/B vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__or2_1
XFILLER_108_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _12161_/A _12325_/A _12161_/C vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__nor3_2
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11112_/A _11112_/B _11112_/C vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__or3_4
XFILLER_122_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12092_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__o21ai_4
XFILLER_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15920_ _16315_/C _16499_/B vssd1 vssd1 vccd1 vccd1 _15921_/B sky130_fd_sc_hd__nor2_1
X_11043_ _11043_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15851_ _16446_/A _16041_/A vssd1 vssd1 vccd1 vccd1 _15853_/B sky130_fd_sc_hd__nor2_8
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14802_ _14801_/B _14801_/C _11100_/A vssd1 vssd1 vccd1 vccd1 _14803_/B sky130_fd_sc_hd__o21a_1
XTAP_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15782_ _15782_/A _15782_/B vssd1 vssd1 vccd1 vccd1 _15784_/B sky130_fd_sc_hd__nand2_1
XTAP_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12994_ _12993_/A _12993_/B _12991_/X vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__o21ba_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17521_ fanout931/X _17521_/D vssd1 vssd1 vccd1 vccd1 _17521_/Q sky130_fd_sc_hd__dfxtp_4
X_14733_ _13624_/B _13627_/X _14840_/A vssd1 vssd1 vccd1 vccd1 _14734_/B sky130_fd_sc_hd__mux2_2
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11945_ _09006_/X _09010_/A _11943_/Y _11944_/X vssd1 vssd1 vccd1 vccd1 _12156_/B
+ sky130_fd_sc_hd__a211o_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ fanout941/X _17452_/D vssd1 vssd1 vccd1 vccd1 _17452_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _14664_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14664_/X sky130_fd_sc_hd__or2_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11876_ _11877_/A _11877_/B _11877_/C vssd1 vssd1 vccd1 vccd1 _11891_/A sky130_fd_sc_hd__a21oi_4
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ _16735_/A _14036_/X _14926_/X _15040_/X vssd1 vssd1 vccd1 vccd1 _16404_/C
+ sky130_fd_sc_hd__o22a_1
X_13615_ _13501_/B _13503_/B _13501_/A vssd1 vssd1 vccd1 vccd1 _13618_/B sky130_fd_sc_hd__o21ba_2
XFILLER_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10827_ _10827_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__nor2_2
X_17383_ _17383_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17383_/X sky130_fd_sc_hd__or2_1
X_14595_ _14676_/A _14641_/C vssd1 vssd1 vccd1 vccd1 _14597_/B sky130_fd_sc_hd__and2_4
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ _16814_/A _16827_/A _16747_/A _16827_/B vssd1 vssd1 vccd1 vccd1 _16335_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13546_ _13418_/A _13419_/Y _13662_/A _13545_/X vssd1 vssd1 vccd1 vccd1 _13662_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10758_ _10757_/A _10757_/B _10757_/C vssd1 vssd1 vccd1 vccd1 _10759_/B sky130_fd_sc_hd__o21ai_1
XFILLER_185_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16265_ _16172_/A _16172_/B _16170_/A vssd1 vssd1 vccd1 vccd1 _16266_/B sky130_fd_sc_hd__o21ai_4
XFILLER_187_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13477_ _13477_/A _13477_/B vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10689_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10689_/X sky130_fd_sc_hd__and2_1
XFILLER_127_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ _15216_/A _15216_/B vssd1 vssd1 vccd1 vccd1 _15218_/B sky130_fd_sc_hd__xor2_4
XFILLER_127_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12428_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__o21a_2
X_16196_ _16197_/A _16197_/B _16195_/Y vssd1 vssd1 vccd1 vccd1 _16290_/B sky130_fd_sc_hd__o21ba_1
XFILLER_127_986 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15147_ _15147_/A _17614_/Q _15147_/C _15270_/A vssd1 vssd1 vccd1 vccd1 _15147_/Y
+ sky130_fd_sc_hd__nor4_2
X_12359_ _12526_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__a21o_2
XFILLER_126_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15078_ _14898_/Y _15077_/Y _11377_/D vssd1 vssd1 vccd1 vccd1 _15647_/A sky130_fd_sc_hd__o21a_4
XFILLER_102_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14029_ _14030_/A _14030_/B _14030_/C vssd1 vssd1 vccd1 vccd1 _14029_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09570_ _09567_/Y _09570_/B vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__and2b_2
XFILLER_64_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09004_ _09004_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09007_/A sky130_fd_sc_hd__xnor2_2
XFILLER_192_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout500 _17518_/Q vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__buf_6
XFILLER_116_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout511 _15373_/C vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__buf_6
X_09906_ _09906_/A _09906_/B _10035_/A vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__nand3_1
Xfanout522 _10640_/C vssd1 vssd1 vccd1 vccd1 _15305_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_120_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout533 _10419_/A vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__buf_6
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout544 _09470_/B vssd1 vssd1 vccd1 vccd1 _12847_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout555 _15538_/A vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__buf_6
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout566 _10299_/C vssd1 vssd1 vccd1 vccd1 _16011_/A sky130_fd_sc_hd__buf_4
X_09837_ _09842_/A _09842_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__nor2_2
XFILLER_47_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout577 _17164_/B vssd1 vssd1 vccd1 vccd1 _16011_/B sky130_fd_sc_hd__buf_4
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout588 _12398_/S vssd1 vssd1 vccd1 vccd1 _14958_/A sky130_fd_sc_hd__buf_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout599 _10430_/A vssd1 vssd1 vccd1 vccd1 _11839_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _09768_/A _09768_/B _09832_/A vssd1 vssd1 vccd1 vccd1 _09769_/D sky130_fd_sc_hd__or3_1
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _12135_/B vssd1 vssd1 vccd1 vccd1 _08719_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09699_ _09699_/A _09706_/A vssd1 vssd1 vccd1 vccd1 _09701_/C sky130_fd_sc_hd__nor2_1
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _11731_/B _11736_/A _11731_/A vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__o21a_2
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11662_/A _11662_/B vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__and2b_1
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _13950_/A _13895_/C _13282_/A _13280_/B vssd1 vssd1 vccd1 vccd1 _13401_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_186_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10612_ _10598_/X _10611_/Y _10499_/Y _10589_/X vssd1 vssd1 vccd1 vccd1 _10632_/A
+ sky130_fd_sc_hd__a211o_4
X_14380_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__and2_2
X_11592_ _11629_/A _14792_/B vssd1 vssd1 vccd1 vccd1 _14796_/A sky130_fd_sc_hd__nand2_2
XFILLER_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13332_/A _13332_/B _13332_/C vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__a21oi_4
X_10543_ _15126_/A _10543_/B _10543_/C vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__and3_1
XFILLER_127_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16050_ _16051_/B _16051_/A vssd1 vssd1 vccd1 vccd1 _16183_/A sky130_fd_sc_hd__and2b_1
X_13262_ _13261_/A _13261_/B _13261_/C vssd1 vssd1 vccd1 vccd1 _13263_/B sky130_fd_sc_hd__a21o_1
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _10405_/B _10405_/C _10405_/D _10405_/A vssd1 vssd1 vccd1 vccd1 _10474_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_183_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15001_ _14995_/X _15538_/B _15538_/A vssd1 vssd1 vccd1 vccd1 _15001_/X sky130_fd_sc_hd__mux2_2
XFILLER_68_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12213_ _12211_/X _12212_/X _15384_/S vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__mux2_1
X_13193_ _17423_/A _13321_/D _13194_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _13195_/A
+ sky130_fd_sc_hd__a22oi_2
X_12144_ _12145_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__nand2_2
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16952_ _16952_/A _16952_/B _16952_/C vssd1 vssd1 vccd1 vccd1 _16953_/B sky130_fd_sc_hd__and3_1
X_12075_ _12075_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11026_ _11026_/A _11605_/B vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__nand2_4
X_15903_ _14666_/S _15901_/X _15902_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15903_/X
+ sky130_fd_sc_hd__a211o_1
X_16883_ _16938_/B _16938_/D _16883_/C vssd1 vssd1 vccd1 vccd1 _16884_/B sky130_fd_sc_hd__or3_1
XFILLER_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15834_ _15834_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15836_/B sky130_fd_sc_hd__xnor2_4
XTAP_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_951 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _15765_/A _15868_/B _15765_/C vssd1 vssd1 vccd1 vccd1 _15866_/B sky130_fd_sc_hd__nor3_2
X_12977_ _12976_/A _12976_/B _12975_/X vssd1 vssd1 vccd1 vccd1 _12978_/B sky130_fd_sc_hd__o21bai_2
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ fanout933/X _17504_/D vssd1 vssd1 vccd1 vccd1 _17504_/Q sky130_fd_sc_hd__dfxtp_2
X_14716_ _14717_/A _14717_/B vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__or2_1
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11928_ _11930_/B _12752_/B vssd1 vssd1 vccd1 vccd1 _12470_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15696_ _15603_/Y _15606_/Y _15786_/B _15695_/X vssd1 vssd1 vccd1 vccd1 _15698_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _14594_/A _14596_/Y _14594_/B vssd1 vssd1 vccd1 vccd1 _14649_/A sky130_fd_sc_hd__o21bai_4
X_17435_ fanout925/X _17435_/D vssd1 vssd1 vccd1 vccd1 _17435_/Q sky130_fd_sc_hd__dfxtp_4
X_11859_ _12068_/A _12068_/B _11859_/C _12637_/C vssd1 vssd1 vccd1 vccd1 _11860_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 _17542_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_29 _17465_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _14627_/B sky130_fd_sc_hd__nor2_1
X_17366_ input47/X _17377_/B _17365_/Y _17372_/C1 vssd1 vssd1 vccd1 vccd1 _17511_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13529_ _13527_/X _13529_/B vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__and2b_2
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16317_ _16317_/A _16317_/B vssd1 vssd1 vccd1 vccd1 _16504_/B sky130_fd_sc_hd__nand2_4
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17297_ input36/X _17362_/C _17429_/C vssd1 vssd1 vccd1 vccd1 _17297_/X sky130_fd_sc_hd__or3_1
XFILLER_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16248_ _16248_/A _16248_/B vssd1 vssd1 vccd1 vccd1 _16250_/C sky130_fd_sc_hd__nor2_1
XFILLER_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 _17461_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[27] sky130_fd_sc_hd__clkbuf_2
X_16179_ _16179_/A _16179_/B vssd1 vssd1 vccd1 vccd1 _16180_/B sky130_fd_sc_hd__nor2_1
Xoutput114 _17442_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09622_ _09629_/A _09601_/Y _09616_/Y _09621_/X vssd1 vssd1 vccd1 vccd1 _09626_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09553_ _09559_/B _09559_/A vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__and2b_1
XFILLER_110_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ _09484_/A _09484_/B _09484_/C vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__and3_4
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10190_ _10188_/A _10188_/Y _10207_/A _10161_/X vssd1 vssd1 vccd1 vccd1 _10207_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout330 _12620_/A vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__buf_12
Xfanout341 _14599_/A vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__clkbuf_16
Xfanout352 _12659_/A vssd1 vssd1 vccd1 vccd1 _12176_/A sky130_fd_sc_hd__clkbuf_8
Xfanout363 _17413_/A vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__buf_4
XFILLER_28_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1041 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout374 _12488_/A vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__buf_4
Xfanout385 _17407_/A vssd1 vssd1 vccd1 vccd1 _14248_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout396 _17530_/Q vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__buf_6
XFILLER_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _12900_/A _13049_/B vssd1 vssd1 vccd1 vccd1 _12902_/C sky130_fd_sc_hd__nand2_1
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13880_ _13880_/A _13880_/B vssd1 vssd1 vccd1 vccd1 _13882_/B sky130_fd_sc_hd__xnor2_4
XFILLER_143_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12831_ _12991_/A _12829_/Y _12672_/X _12674_/Y vssd1 vssd1 vccd1 vccd1 _12834_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15550_ _15071_/A _14888_/B _15262_/B vssd1 vssd1 vccd1 vccd1 _15552_/B sky130_fd_sc_hd__a21bo_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12928_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _12764_/C sky130_fd_sc_hd__or2_2
XFILLER_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14500_/B _14501_/B vssd1 vssd1 vccd1 vccd1 _14562_/B sky130_fd_sc_hd__nand2b_1
XFILLER_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _16206_/B sky130_fd_sc_hd__xor2_2
X_15481_ _15481_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15504_/A sky130_fd_sc_hd__xnor2_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12694_/A _12694_/B vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__or2_1
XFILLER_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _13977_/B _14593_/C _17028_/A _14599_/A vssd1 vssd1 vccd1 vccd1 _14432_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17550_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__and2_1
X_11644_ _11607_/B _11648_/A _11644_/C vssd1 vssd1 vccd1 vccd1 _11644_/X sky130_fd_sc_hd__and3b_1
XFILLER_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17151_ _17151_/A _17151_/B vssd1 vssd1 vccd1 vccd1 _17167_/C sky130_fd_sc_hd__nand2_1
X_14363_ _14364_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _14440_/B sky130_fd_sc_hd__nor2_1
XFILLER_168_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 i_wb_addr[21] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_2
X_11575_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__nor2_2
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput27 i_wb_addr[31] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16102_ _15991_/X _15994_/X _16100_/Y _16911_/A vssd1 vssd1 vccd1 vccd1 _16102_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ _13314_/A _13314_/B _13314_/C vssd1 vssd1 vccd1 vccd1 _13315_/B sky130_fd_sc_hd__or3_1
Xinput38 i_wb_data[11] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10526_ _10971_/A _10640_/D _10933_/D _10525_/A vssd1 vssd1 vccd1 vccd1 _10526_/Y
+ sky130_fd_sc_hd__a22oi_2
X_17082_ _11026_/A _10791_/C _17038_/B _10254_/A _10036_/D vssd1 vssd1 vccd1 vccd1
+ _17083_/C sky130_fd_sc_hd__a32o_1
Xinput49 i_wb_data[21] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
X_14294_ _14294_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _14295_/B sky130_fd_sc_hd__and2_1
XFILLER_182_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16033_ _16136_/B _16745_/B vssd1 vssd1 vccd1 vccd1 _16034_/B sky130_fd_sc_hd__nand2_4
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ _13244_/B _13244_/C _13244_/A vssd1 vssd1 vccd1 vccd1 _13246_/B sky130_fd_sc_hd__a21o_1
X_10457_ _10319_/Y _10354_/X _10407_/Y _10442_/Y vssd1 vssd1 vccd1 vccd1 _10459_/C
+ sky130_fd_sc_hd__a211o_4
XFILLER_123_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _13176_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _13178_/C sky130_fd_sc_hd__xnor2_4
X_10388_ _10388_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10390_/C sky130_fd_sc_hd__or2_2
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12127_ _12618_/A _12770_/B _12127_/C _12127_/D vssd1 vssd1 vccd1 vccd1 _12343_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16935_ _16935_/A _16935_/B _16935_/C vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__and3_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12058_ _12038_/X _12057_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ _11009_/A _11009_/B vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__xor2_4
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16866_ _16866_/A _16866_/B vssd1 vssd1 vccd1 vccd1 _16866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_92_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15817_ _16809_/A _16020_/B vssd1 vssd1 vccd1 vccd1 _15817_/X sky130_fd_sc_hd__and2_2
XFILLER_34_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16797_ _16797_/A _16797_/B vssd1 vssd1 vccd1 vccd1 _16797_/X sky130_fd_sc_hd__xor2_1
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15748_ _15414_/B _15746_/X _15747_/X vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__o21a_2
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15679_ _15679_/A _15772_/B _15679_/C vssd1 vssd1 vccd1 vccd1 _15769_/B sky130_fd_sc_hd__and3_2
XFILLER_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17418_ input55/X _17426_/A2 _17417_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17537_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_178_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17349_ input54/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17349_/X sky130_fd_sc_hd__or3_1
XFILLER_186_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08984_ _09242_/B _08984_/B vssd1 vssd1 vccd1 vccd1 _08985_/C sky130_fd_sc_hd__nand2_1
XFILLER_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09605_ _09748_/B _10545_/D _10753_/B _09748_/A vssd1 vssd1 vccd1 vccd1 _09605_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09536_ _09536_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__nor2_2
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09467_ _15538_/A _11808_/B _09462_/A _09326_/Y vssd1 vssd1 vccd1 vccd1 _09468_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_157_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09398_ _09393_/B _09393_/C _09393_/D _09395_/B vssd1 vssd1 vccd1 vccd1 _09398_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11360_ _11354_/A _11354_/C _11354_/B vssd1 vssd1 vccd1 vccd1 _11361_/B sky130_fd_sc_hd__o21ai_2
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10311_ _10312_/A _10310_/Y _12398_/S _10311_/D vssd1 vssd1 vccd1 vccd1 _10429_/A
+ sky130_fd_sc_hd__and4bb_4
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11293_/B sky130_fd_sc_hd__and2_1
XFILLER_180_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13030_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13165_/B sky130_fd_sc_hd__nand2_2
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10242_ _10694_/B _10912_/C _10479_/B _10694_/A vssd1 vssd1 vccd1 vccd1 _10243_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_65_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10173_ _10288_/A _10172_/Y _15711_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _10296_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout160 _17419_/B vssd1 vssd1 vccd1 vccd1 _17397_/B sky130_fd_sc_hd__clkbuf_4
X_14981_ _14981_/A _14981_/B vssd1 vssd1 vccd1 vccd1 _14981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout171 _15726_/D vssd1 vssd1 vccd1 vccd1 _16743_/C sky130_fd_sc_hd__buf_6
XFILLER_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout182 _15472_/Y vssd1 vssd1 vccd1 vccd1 _16827_/A sky130_fd_sc_hd__buf_6
X_16720_ _16723_/A _16644_/B _16722_/A vssd1 vssd1 vccd1 vccd1 _16791_/A sky130_fd_sc_hd__a21bo_1
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ _13932_/A _13932_/B vssd1 vssd1 vccd1 vccd1 _14122_/A sky130_fd_sc_hd__xnor2_2
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13863_ _13964_/A _13862_/C _13862_/A vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16651_ _16651_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16652_/C sky130_fd_sc_hd__nor2_1
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12814_ _12976_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__xor2_4
X_15602_ _15505_/A _15505_/B _15511_/X vssd1 vssd1 vccd1 vccd1 _15604_/B sky130_fd_sc_hd__a21oi_4
X_13794_ _13793_/A _13793_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__o21ai_2
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16582_ _16582_/A _16582_/B vssd1 vssd1 vccd1 vccd1 _16582_/X sky130_fd_sc_hd__or2_1
XFILLER_188_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12585_/B _12585_/C _12585_/A vssd1 vssd1 vccd1 vccd1 _12747_/B sky130_fd_sc_hd__a21bo_4
X_15533_ _15533_/A _15533_/B vssd1 vssd1 vccd1 vccd1 _15533_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15464_ _14805_/B _15899_/A2 _15713_/B1 _15463_/A _14944_/A vssd1 vssd1 vccd1 vccd1
+ _15464_/X sky130_fd_sc_hd__a221o_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__or3_2
XFILLER_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _14352_/A _14349_/X _14351_/B vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__o21a_1
X_17203_ _17435_/Q _17233_/A2 _17201_/X _17202_/X _17428_/B vssd1 vssd1 vccd1 vccd1
+ _17435_/D sky130_fd_sc_hd__o221a_1
X_11627_ _11613_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__a21o_1
X_15395_ _15396_/A _15396_/B _15472_/B vssd1 vssd1 vccd1 vccd1 _16152_/A sky130_fd_sc_hd__and3_4
XFILLER_11_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14346_ _14254_/A _14554_/B _14255_/A _14253_/A vssd1 vssd1 vccd1 vccd1 _14348_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_155_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17134_ _17134_/A _17134_/B _17134_/C vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__and3_1
XFILLER_184_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _11558_/A _11558_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__nand3_1
XFILLER_183_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _17065_/A _17153_/B _14765_/A vssd1 vssd1 vccd1 vccd1 _17065_/X sky130_fd_sc_hd__or3b_4
XFILLER_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _10509_/A _10617_/A vssd1 vssd1 vccd1 vccd1 _10511_/B sky130_fd_sc_hd__nor2_2
XFILLER_170_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14277_ _14352_/A _14277_/B vssd1 vssd1 vccd1 vccd1 _14283_/B sky130_fd_sc_hd__nand2b_1
X_11489_ _11496_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__or2_4
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16016_ _15309_/B _16004_/Y _16007_/X _16015_/X vssd1 vssd1 vccd1 vccd1 _16017_/C
+ sky130_fd_sc_hd__o211a_1
X_13228_ _13228_/A _13228_/B vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13159_ _13159_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13161_/B sky130_fd_sc_hd__xnor2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16918_ _16918_/A _16918_/B _16918_/C vssd1 vssd1 vccd1 vccd1 _16918_/X sky130_fd_sc_hd__and3_1
XFILLER_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16849_ _16850_/A _16850_/B vssd1 vssd1 vccd1 vccd1 _16851_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _09328_/A _09320_/Y _09750_/C _10309_/B vssd1 vssd1 vccd1 vccd1 _09451_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_179_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _09182_/Y _09342_/A _09250_/Y _09251_/X vssd1 vssd1 vccd1 vccd1 _09255_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09183_ _09155_/Y _09156_/X _09179_/A _09346_/A vssd1 vssd1 vccd1 vccd1 _09214_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_159_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08967_ _09779_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _12700_/C sky130_fd_sc_hd__and2_4
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08898_ _12258_/A _12950_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__nand2_4
XFILLER_5_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _10860_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10861_/C sky130_fd_sc_hd__xnor2_4
X_09519_ _09519_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09520_/C sky130_fd_sc_hd__xnor2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10791_ _11561_/A _11629_/B _10791_/C _10791_/D vssd1 vssd1 vccd1 vccd1 _10794_/A
+ sky130_fd_sc_hd__and4_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12530_ _12530_/A _12530_/B vssd1 vssd1 vccd1 vccd1 _12534_/A sky130_fd_sc_hd__or2_4
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12307_/A _12307_/B _12306_/A vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__a21o_4
XFILLER_138_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ _14200_/A _14200_/B _14198_/X vssd1 vssd1 vccd1 vccd1 _14201_/B sky130_fd_sc_hd__or3b_1
X_11412_ _11419_/A _11419_/B _11410_/Y vssd1 vssd1 vccd1 vccd1 _11413_/C sky130_fd_sc_hd__a21oi_4
X_15180_ _16011_/B _15180_/B vssd1 vssd1 vccd1 vccd1 _15180_/X sky130_fd_sc_hd__or2_2
X_12392_ _12035_/C _12033_/Y _15095_/B vssd1 vssd1 vccd1 vccd1 _12393_/B sky130_fd_sc_hd__mux2_2
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14131_ _14131_/A vssd1 vssd1 vccd1 vccd1 _14138_/A sky130_fd_sc_hd__inv_2
XFILLER_153_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11343_ _11343_/A _11349_/A vssd1 vssd1 vccd1 vccd1 _11352_/B sky130_fd_sc_hd__and2_2
XFILLER_193_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14062_ _13977_/B _14063_/C _14213_/C _14599_/A vssd1 vssd1 vccd1 vccd1 _14064_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_180_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11274_ _11274_/A _11274_/B _11274_/C vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__nand3_2
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _15457_/B _13012_/X _17165_/A1 vssd1 vssd1 vccd1 vccd1 _13013_/Y sky130_fd_sc_hd__o21ai_1
X_10225_ _10348_/A _10348_/B _10348_/C vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__o21ai_4
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ _10005_/X _10105_/Y _10134_/A _10134_/Y vssd1 vssd1 vccd1 vccd1 _10157_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _10060_/Y _10216_/A _09959_/X _09972_/Y vssd1 vssd1 vccd1 vccd1 _10090_/A
+ sky130_fd_sc_hd__a211oi_4
X_14964_ _14961_/X _14963_/X _14927_/X _14945_/X vssd1 vssd1 vccd1 vccd1 _14964_/Y
+ sky130_fd_sc_hd__o211ai_4
X_16703_ _16628_/A _16628_/B _16617_/A vssd1 vssd1 vccd1 vccd1 _16705_/B sky130_fd_sc_hd__a21oi_1
X_13915_ _13915_/A _13915_/B _13915_/C vssd1 vssd1 vccd1 vccd1 _13916_/B sky130_fd_sc_hd__nor3_1
XFILLER_81_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14895_ _15530_/A _15450_/A vssd1 vssd1 vccd1 vccd1 _14905_/C sky130_fd_sc_hd__or2_1
XFILLER_48_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16634_ _16634_/A _16634_/B vssd1 vssd1 vccd1 vccd1 _16636_/C sky130_fd_sc_hd__xnor2_1
X_13846_ _13950_/A _13948_/D vssd1 vssd1 vccd1 vccd1 _13848_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16565_ _16203_/X _16293_/A _16561_/X _16562_/Y _16564_/Y vssd1 vssd1 vccd1 vccd1
+ _16566_/B sky130_fd_sc_hd__o311a_4
X_13777_ _13778_/A _13778_/B _13778_/C vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__o21a_1
XFILLER_188_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__a21o_1
X_15516_ _15774_/A _15667_/B _15431_/A _15428_/X vssd1 vssd1 vccd1 vccd1 _15518_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ _12886_/B _12728_/B vssd1 vssd1 vccd1 vccd1 _12730_/C sky130_fd_sc_hd__or2_2
X_16496_ _16814_/A _16662_/C _16662_/D _16667_/A vssd1 vssd1 vccd1 vccd1 _16498_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12659_ _12659_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__nand2_2
X_15447_ _15447_/A _16207_/B vssd1 vssd1 vccd1 vccd1 _15447_/X sky130_fd_sc_hd__or2_1
XFILLER_157_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15378_ _10800_/C _14803_/A _14803_/B vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17117_ _17096_/A _17096_/B _17093_/Y _17095_/B vssd1 vssd1 vccd1 vccd1 _17130_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14329_ _14330_/A _14330_/B _14330_/C vssd1 vssd1 vccd1 vccd1 _14409_/A sky130_fd_sc_hd__a21oi_4
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ _17049_/A _17049_/B vssd1 vssd1 vccd1 vccd1 _17088_/B sky130_fd_sc_hd__and2_1
XFILLER_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__nand3_2
Xfanout907 _17270_/B1 vssd1 vssd1 vccd1 vccd1 _17288_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout918 _17372_/C1 vssd1 vssd1 vccd1 vccd1 _17428_/B sky130_fd_sc_hd__buf_4
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout929 input2/X vssd1 vssd1 vccd1 vccd1 fanout929/X sky130_fd_sc_hd__buf_4
XFILLER_86_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A _08822_/A _08821_/C vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__or3_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08755_/A vssd1 vssd1 vccd1 vccd1 _08754_/C sky130_fd_sc_hd__inv_2
XFILLER_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09304_ _09304_/A _09304_/B vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09235_ _12176_/A _12174_/D vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09166_ _12772_/A _09172_/B _17466_/D _11920_/B vssd1 vssd1 vccd1 vccd1 _09167_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_147_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _10542_/A _17508_/Q vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__and2_2
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10010_ _10010_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09999_ _10254_/B _10736_/C _10392_/D _10254_/A vssd1 vssd1 vccd1 vccd1 _10000_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_49_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ _12166_/A _11961_/B _11961_/C vssd1 vssd1 vccd1 vccd1 _12169_/B sky130_fd_sc_hd__nand3_1
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13700_ _13800_/B _13700_/B vssd1 vssd1 vccd1 vccd1 _13702_/C sky130_fd_sc_hd__nand2_1
X_10912_ _11095_/A _11240_/A _10912_/C _11005_/B vssd1 vssd1 vccd1 vccd1 _10914_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14680_/A _14708_/C _14680_/C vssd1 vssd1 vccd1 vccd1 _14682_/B sky130_fd_sc_hd__nand3_4
XFILLER_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11892_ _08801_/A _08801_/Y _11890_/X _11891_/Y vssd1 vssd1 vccd1 vccd1 _11915_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13631_ _13844_/B _14089_/B _13523_/B _13844_/A vssd1 vssd1 vccd1 vccd1 _13635_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10843_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10943_/A sky130_fd_sc_hd__nand2b_2
XFILLER_73_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16350_ _16252_/A _16252_/B _16251_/A vssd1 vssd1 vccd1 vccd1 _16362_/A sky130_fd_sc_hd__a21o_2
X_13562_ _13562_/A _13562_/B vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__nor2_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10774_ _10774_/A _10774_/B _10774_/C vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__nor3_4
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12513_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__nor2_4
X_15301_ _15233_/X _15299_/Y _15300_/Y vssd1 vssd1 vccd1 vccd1 _15301_/Y sky130_fd_sc_hd__o21ai_1
X_16281_ _16281_/A _16695_/B vssd1 vssd1 vccd1 vccd1 _16282_/B sky130_fd_sc_hd__nand2_4
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13493_ _13494_/A _13494_/B _13494_/C vssd1 vssd1 vccd1 vccd1 _13495_/A sky130_fd_sc_hd__o21a_2
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12444_ _17383_/A _12736_/B _12578_/B _17385_/A vssd1 vssd1 vccd1 vccd1 _12446_/A
+ sky130_fd_sc_hd__a22oi_4
X_15232_ _15171_/A _15171_/B _15168_/Y vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__a21boi_1
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15163_ _15821_/A _15774_/A _15164_/B vssd1 vssd1 vccd1 vccd1 _15165_/A sky130_fd_sc_hd__a21o_1
X_12375_ _12375_/A _12375_/B vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14114_ _14202_/A _14114_/B vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11326_ _11320_/A _11320_/C _11320_/B vssd1 vssd1 vccd1 vccd1 _11327_/B sky130_fd_sc_hd__o21ai_1
XFILLER_180_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15094_ _15094_/A _15170_/C vssd1 vssd1 vccd1 vccd1 _15094_/X sky130_fd_sc_hd__xor2_2
XFILLER_180_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14045_ _14134_/B _14045_/B vssd1 vssd1 vccd1 vccd1 _14047_/B sky130_fd_sc_hd__xnor2_1
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11274_/A sky130_fd_sc_hd__xnor2_4
XFILLER_80_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__and2_1
XFILLER_192_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11188_ _11053_/Y _11055_/X _11218_/B _11187_/X vssd1 vssd1 vccd1 vccd1 _11222_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10139_ _10508_/C _10745_/D _10017_/A _10015_/Y vssd1 vssd1 vccd1 vccd1 _10140_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15996_ _15994_/A _15993_/X _15995_/Y vssd1 vssd1 vccd1 vccd1 _15996_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14947_ _15100_/A _14947_/B vssd1 vssd1 vccd1 vccd1 _15180_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14878_ _15147_/C _14888_/B _14877_/Y vssd1 vssd1 vccd1 vccd1 _14878_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16617_ _16617_/A _16617_/B vssd1 vssd1 vccd1 vccd1 _16628_/A sky130_fd_sc_hd__nor2_4
XFILLER_51_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ _13936_/B _13830_/B vssd1 vssd1 vccd1 vccd1 _13829_/Y sky130_fd_sc_hd__nand2_1
X_17597_ fanout943/X _17597_/D vssd1 vssd1 vccd1 vccd1 _17597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16548_ _16630_/B _16548_/B vssd1 vssd1 vccd1 vccd1 _16550_/C sky130_fd_sc_hd__nand2_1
XFILLER_189_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16479_ _14775_/A _16644_/B _16480_/A vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__a21bo_1
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__xnor2_4
XFILLER_176_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__or2_1
Xfanout704 _13094_/B vssd1 vssd1 vccd1 vccd1 _11881_/D sky130_fd_sc_hd__buf_6
XFILLER_59_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout715 _12077_/C vssd1 vssd1 vccd1 vccd1 _10545_/D sky130_fd_sc_hd__clkbuf_8
Xfanout726 _16399_/A vssd1 vssd1 vccd1 vccd1 _13866_/C sky130_fd_sc_hd__buf_6
XFILLER_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09853_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__nand2b_1
Xfanout737 _17494_/Q vssd1 vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__buf_12
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 fanout757/X vssd1 vssd1 vccd1 vccd1 _13100_/B sky130_fd_sc_hd__buf_4
XFILLER_140_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout759 _17492_/Q vssd1 vssd1 vccd1 vccd1 _12637_/C sky130_fd_sc_hd__buf_12
XFILLER_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08804_ _08804_/A _08804_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__nor2_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09784_ _09784_/A _09784_/B _09784_/C vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__or3_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08735_ _15147_/A _14836_/B _17131_/A vssd1 vssd1 vccd1 vccd1 _17613_/D sky130_fd_sc_hd__mux2_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ _09219_/A _11958_/A _09219_/C vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__o21a_1
XFILLER_10_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10490_ _11006_/A _11006_/B _10490_/C _10490_/D vssd1 vssd1 vccd1 vccd1 _10493_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09149_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09245_/B sky130_fd_sc_hd__nand2b_2
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _12161_/A _12325_/A _12161_/C vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__o21a_1
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _10893_/A _10893_/B _10893_/C vssd1 vssd1 vccd1 vccd1 _11112_/C sky130_fd_sc_hd__a21oi_4
X_12091_ _12091_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12093_/C sky130_fd_sc_hd__xnor2_4
X_11042_ _11041_/A _11041_/B _11041_/C vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__a21o_1
XFILLER_77_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15850_ _15850_/A _15850_/B vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__xor2_4
XTAP_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14801_ _14801_/A _14801_/B _14801_/C vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__or3_1
XTAP_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15781_ _15781_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15784_/A sky130_fd_sc_hd__xnor2_1
XTAP_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _12993_/A _12993_/B _12991_/X vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__or3b_2
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17520_ fanout931/X _17520_/D vssd1 vssd1 vccd1 vccd1 _17520_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _14763_/S _14730_/Y _14731_/X _14705_/Y _14706_/X vssd1 vssd1 vccd1 vccd1
+ _17604_/D sky130_fd_sc_hd__a32o_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11944_ _11940_/X _11941_/Y _08868_/X _08873_/C vssd1 vssd1 vccd1 vccd1 _11944_/X
+ sky130_fd_sc_hd__o211a_2
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17451_ fanout938/X _17451_/D vssd1 vssd1 vccd1 vccd1 _17451_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_17_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14663_ _14664_/A _14669_/B vssd1 vssd1 vccd1 vccd1 _14663_/Y sky130_fd_sc_hd__nand2_1
X_11875_ _12085_/B _11875_/B vssd1 vssd1 vccd1 vccd1 _11877_/C sky130_fd_sc_hd__nand2_2
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16402_ _12235_/C _17075_/A2 _16401_/X vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__a21oi_1
XFILLER_189_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13614_ _13614_/A _13614_/B vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__xor2_4
X_10826_ _11258_/B _10911_/B _10912_/C _11115_/A vssd1 vssd1 vccd1 vccd1 _10827_/B
+ sky130_fd_sc_hd__a22oi_4
X_17382_ input67/X _17396_/A2 _17381_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17519_/D
+ sky130_fd_sc_hd__o211a_1
X_14594_ _14594_/A _14594_/B vssd1 vssd1 vccd1 vccd1 _14597_/A sky130_fd_sc_hd__or2_1
XFILLER_158_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16333_ _16827_/A _16747_/A _16827_/B _16814_/A vssd1 vssd1 vccd1 vccd1 _16333_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_185_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13545_ _13545_/A _13545_/B _13545_/C vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__and3_2
X_10757_ _10757_/A _10757_/B _10757_/C vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__or3_2
XFILLER_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16264_ _16358_/B _16264_/B vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__nor2_2
XFILLER_158_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13476_ _13476_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__xor2_1
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _10688_/A _10688_/B vssd1 vssd1 vccd1 vccd1 _10784_/A sky130_fd_sc_hd__nand2_4
XFILLER_173_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12427_ _12427_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12429_/C sky130_fd_sc_hd__xnor2_2
X_15215_ _15662_/A _16136_/B vssd1 vssd1 vccd1 vccd1 _15216_/B sky130_fd_sc_hd__nand2_2
X_16195_ _16195_/A _16195_/B vssd1 vssd1 vccd1 vccd1 _16195_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15146_ _15553_/A _15553_/B _15948_/A vssd1 vssd1 vccd1 vccd1 _15155_/A sky130_fd_sc_hd__or3_4
X_12358_ _12526_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12526_/B sky130_fd_sc_hd__nand3_4
XFILLER_99_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__nand2b_2
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15077_ _15143_/A _15077_/B vssd1 vssd1 vccd1 vccd1 _15077_/Y sky130_fd_sc_hd__nor2_4
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12289_ _12267_/Y _12268_/X _12476_/B _12290_/D vssd1 vssd1 vccd1 vccd1 _12289_/Y
+ sky130_fd_sc_hd__a2bb2oi_4
XFILLER_114_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _14119_/B _14028_/B vssd1 vssd1 vccd1 vccd1 _14030_/C sky130_fd_sc_hd__nand2b_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15979_ _15980_/A _15980_/B _15980_/C vssd1 vssd1 vccd1 vccd1 _15979_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09004_/B sky130_fd_sc_hd__xnor2_4
XFILLER_118_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout501 _14786_/A vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__buf_6
X_09905_ _09909_/A vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__inv_2
Xfanout512 _15373_/C vssd1 vssd1 vccd1 vccd1 _11258_/B sky130_fd_sc_hd__buf_6
XFILLER_99_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout523 _10640_/C vssd1 vssd1 vccd1 vccd1 _11423_/B sky130_fd_sc_hd__buf_2
XFILLER_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout534 _11322_/A vssd1 vssd1 vccd1 vccd1 _10419_/A sky130_fd_sc_hd__buf_6
XFILLER_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout545 fanout554/X vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__buf_4
XFILLER_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout556 _11268_/A vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__buf_6
X_09836_ _10366_/A _10490_/D _09695_/A _09693_/Y vssd1 vssd1 vccd1 vccd1 _09842_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout567 _10299_/C vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__buf_4
Xfanout578 _17512_/Q vssd1 vssd1 vccd1 vccd1 _17164_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 _12398_/S vssd1 vssd1 vccd1 vccd1 _15095_/B sky130_fd_sc_hd__buf_4
XFILLER_101_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09767_ _09761_/A _09765_/X _09776_/A _09745_/Y vssd1 vssd1 vccd1 vccd1 _09776_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08718_/A vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__clkinv_4
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09698_ _10115_/A _10241_/B _10392_/D _10377_/B vssd1 vssd1 vccd1 vccd1 _09706_/A
+ sky130_fd_sc_hd__and4_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11660_ _11678_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11662_/B sky130_fd_sc_hd__nor2_1
XFILLER_187_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _10711_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__nand2_2
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11591_ _11629_/A _14792_/B vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__and2_4
X_13330_ _13330_/A _13330_/B vssd1 vssd1 vccd1 vccd1 _13332_/C sky130_fd_sc_hd__nand2_2
X_10542_ _10542_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _10543_/C sky130_fd_sc_hd__and2_2
XFILLER_168_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _13261_/A _13261_/B _13261_/C vssd1 vssd1 vccd1 vccd1 _13263_/A sky130_fd_sc_hd__nand3_2
XFILLER_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10473_ _10473_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__xnor2_4
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _11809_/Y _11814_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__mux2_1
X_15000_ _14998_/Y _14999_/Y _15254_/S vssd1 vssd1 vccd1 vccd1 _15538_/B sky130_fd_sc_hd__mux2_1
X_13192_ _13188_/X _13190_/Y _13061_/A _13063_/A vssd1 vssd1 vccd1 vccd1 _13202_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_108_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _12143_/A _12143_/B vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__xor2_2
XFILLER_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16951_ _16952_/A _16952_/B _16952_/C vssd1 vssd1 vccd1 vccd1 _16953_/A sky130_fd_sc_hd__a21oi_4
XFILLER_2_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12074_ _12075_/B _12075_/A vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__and2b_2
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11025_ _11025_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11025_/Y sky130_fd_sc_hd__xnor2_1
X_15902_ _13390_/S _15252_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _15902_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16882_ _16882_/A _16882_/B vssd1 vssd1 vccd1 vccd1 _16886_/A sky130_fd_sc_hd__or2_1
XFILLER_49_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ _15834_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15966_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15764_/A _15764_/B _15764_/C vssd1 vssd1 vccd1 vccd1 _15765_/C sky130_fd_sc_hd__and3_1
XFILLER_46_963 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12976_ _12976_/A _12976_/B _12975_/X vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__or3b_2
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17503_ fanout933/X _17503_/D vssd1 vssd1 vccd1 vccd1 _17503_/Q sky130_fd_sc_hd__dfxtp_1
X_14715_ _14742_/A _14715_/B vssd1 vssd1 vccd1 vccd1 _14717_/B sky130_fd_sc_hd__nand2_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ _17375_/A _12102_/D _08856_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _11935_/A
+ sky130_fd_sc_hd__a31o_1
X_15695_ _15786_/A _15693_/Y _15595_/A _15599_/A vssd1 vssd1 vccd1 vccd1 _15695_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ fanout926/X _17434_/D vssd1 vssd1 vccd1 vccd1 _17434_/Q sky130_fd_sc_hd__dfxtp_4
X_14646_ _14646_/A _14646_/B vssd1 vssd1 vccd1 vccd1 _14710_/C sky130_fd_sc_hd__nand2_4
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _12068_/B _11859_/C _12637_/C _12068_/A vssd1 vssd1 vccd1 vccd1 _11860_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 _17434_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _11095_/A _11240_/A _10957_/D _10809_/D vssd1 vssd1 vccd1 vccd1 _10812_/A
+ sky130_fd_sc_hd__and4_1
X_17365_ _17365_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17365_/Y sky130_fd_sc_hd__nand2_1
X_14577_ _14577_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14579_/B sky130_fd_sc_hd__xnor2_1
X_11789_ _15069_/A _11791_/B _16809_/A vssd1 vssd1 vccd1 vccd1 _11789_/X sky130_fd_sc_hd__or3_4
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16316_ _16316_/A _16316_/B vssd1 vssd1 vccd1 vccd1 _16318_/A sky130_fd_sc_hd__nand2_2
X_13528_ _13637_/B _13527_/B _13527_/C vssd1 vssd1 vccd1 vccd1 _13529_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17296_ _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17296_/Y sky130_fd_sc_hd__nor2_2
X_16247_ _16246_/A _16589_/B _16246_/C vssd1 vssd1 vccd1 vccd1 _16248_/B sky130_fd_sc_hd__a21oi_1
X_13459_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__or2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 _17462_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_127_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16178_ _16179_/A _16179_/B vssd1 vssd1 vccd1 vccd1 _16279_/C sky130_fd_sc_hd__and2_2
Xoutput115 _17443_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15129_ _11629_/C _14848_/B _14848_/A _15314_/A _14942_/A _10993_/C vssd1 vssd1 vccd1
+ vccd1 _15129_/X sky130_fd_sc_hd__mux4_1
XFILLER_130_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__and3_4
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09552_ _09552_/A _09696_/A vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__nor2_4
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _09483_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09484_/C sky130_fd_sc_hd__xnor2_4
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout320 _14832_/A vssd1 vssd1 vccd1 vccd1 _14738_/A sky130_fd_sc_hd__buf_6
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout331 _14215_/A vssd1 vssd1 vccd1 vccd1 _14676_/A sky130_fd_sc_hd__buf_6
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout342 _17538_/Q vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout353 _14226_/A vssd1 vssd1 vccd1 vccd1 _16965_/C sky130_fd_sc_hd__buf_6
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout364 _17535_/Q vssd1 vssd1 vccd1 vccd1 _17413_/A sky130_fd_sc_hd__buf_6
XFILLER_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout375 _17533_/Q vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__buf_8
XFILLER_115_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout386 _16723_/A vssd1 vssd1 vccd1 vccd1 _17407_/A sky130_fd_sc_hd__buf_6
X_09819_ _09819_/A _09819_/B _09819_/C vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__nor3_1
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout397 _17530_/Q vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _12672_/X _12674_/Y _12991_/A _12829_/Y vssd1 vssd1 vccd1 vccd1 _12991_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12761_/A _12761_/B _12761_/C vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__nor3_1
XFILLER_188_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14501_/B _14500_/B vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__nand2b_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11713_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _16294_/A sky130_fd_sc_hd__and2_1
X_15480_ _15913_/A _15832_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15590_/A sky130_fd_sc_hd__or3_4
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12533_/X _12536_/B _12532_/Y vssd1 vssd1 vccd1 vccd1 _12694_/B sky130_fd_sc_hd__o21a_1
XFILLER_188_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14497_/B _14431_/B vssd1 vssd1 vccd1 vccd1 _14463_/A sky130_fd_sc_hd__nor2_2
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11607_/B _11644_/C vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__nand2b_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17150_ _17125_/A _17128_/A _17131_/B _17149_/X _14836_/A vssd1 vssd1 vccd1 vccd1
+ _17150_/X sky130_fd_sc_hd__a41o_2
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14362_ _14676_/A _14769_/B vssd1 vssd1 vccd1 vccd1 _14364_/B sky130_fd_sc_hd__nand2_1
X_11574_ _11574_/A _11607_/A _11574_/C vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__or3_4
Xinput17 i_wb_addr[22] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16101_ _15991_/X _15994_/X _16203_/A vssd1 vssd1 vccd1 vccd1 _16101_/Y sky130_fd_sc_hd__o21bai_4
Xinput28 i_wb_addr[3] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_6
X_13313_ _13314_/B _13314_/C _13314_/A vssd1 vssd1 vccd1 vccd1 _13442_/A sky130_fd_sc_hd__o21ai_4
X_10525_ _10525_/A _10971_/A _10640_/D _10933_/D vssd1 vssd1 vccd1 vccd1 _10528_/A
+ sky130_fd_sc_hd__and4_2
Xinput39 i_wb_data[12] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
X_14293_ _14294_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__nor2_2
X_17081_ _17081_/A _17081_/B _17038_/B vssd1 vssd1 vccd1 vccd1 _17083_/B sky130_fd_sc_hd__or3b_1
XFILLER_156_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16032_ _16032_/A _16032_/B vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__or2_4
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13244_ _13244_/A _13244_/B _13244_/C vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__nand3_4
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _10564_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__xor2_4
XFILLER_136_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ _13176_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _13314_/C sky130_fd_sc_hd__and2b_1
XFILLER_184_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10387_ _10387_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10388_/B sky130_fd_sc_hd__nor2_1
XFILLER_123_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12126_ _12770_/B _12127_/C _12127_/D _12618_/A vssd1 vssd1 vccd1 vccd1 _12128_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16934_ _16990_/A _09852_/A _17083_/A _16933_/Y vssd1 vssd1 vccd1 vccd1 _16935_/C
+ sky130_fd_sc_hd__o211a_4
X_12057_ _12047_/X _12056_/X _13838_/S vssd1 vssd1 vccd1 vccd1 _12057_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11008_ _10957_/D _11006_/X _11007_/X vssd1 vssd1 vccd1 vccd1 _11009_/B sky130_fd_sc_hd__a21bo_2
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16865_ _16865_/A _16865_/B vssd1 vssd1 vccd1 vccd1 _16865_/Y sky130_fd_sc_hd__xnor2_1
X_15816_ _15816_/A _16168_/B vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__nor2_4
XFILLER_93_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16796_ _16796_/A _16796_/B vssd1 vssd1 vccd1 vccd1 _16797_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15747_ _16055_/A _15956_/B _16165_/B _16056_/A vssd1 vssd1 vccd1 vccd1 _15747_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _12959_/A _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15678_ _15674_/X _15676_/A _15572_/Y _15583_/Y vssd1 vssd1 vccd1 vccd1 _15679_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_61_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17417_ _17417_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17417_/X sky130_fd_sc_hd__or2_1
X_14629_ _14629_/A _14629_/B _14629_/C vssd1 vssd1 vccd1 vccd1 _14631_/A sky130_fd_sc_hd__and3_2
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17348_ _12734_/D _17354_/A2 _17347_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17503_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17279_ _17602_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17279_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08983_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__or2_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09748_/A _09748_/B _10545_/D _10753_/B vssd1 vssd1 vccd1 vccd1 _09607_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _12005_/B _09397_/X _09531_/X _09540_/A vssd1 vssd1 vccd1 vccd1 _09536_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09466_ _09473_/A _09465_/Y _09750_/C _10311_/D vssd1 vssd1 vccd1 vccd1 _09591_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_184_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09397_ _12005_/A _09395_/X _09343_/X _09392_/B vssd1 vssd1 vccd1 vccd1 _09397_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10310_ _09780_/A _10308_/B _09926_/C vssd1 vssd1 vccd1 vccd1 _10310_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ _11295_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11290_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_98_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ _10694_/A _10241_/B _10912_/C _10805_/C vssd1 vssd1 vccd1 vccd1 _10243_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_191_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _10171_/B _10659_/D _10755_/D _14789_/A vssd1 vssd1 vccd1 vccd1 _10172_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_191_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14980_ _15096_/S _14978_/Y _14979_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _15252_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout150 _15059_/A vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__buf_4
Xfanout161 _17419_/B vssd1 vssd1 vccd1 vccd1 _17425_/B sky130_fd_sc_hd__clkbuf_4
Xfanout172 _16352_/B vssd1 vssd1 vccd1 vccd1 _16809_/C sky130_fd_sc_hd__buf_4
XFILLER_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout183 _15472_/Y vssd1 vssd1 vccd1 vccd1 _16039_/B sky130_fd_sc_hd__clkbuf_4
X_13931_ _13932_/A _13932_/B vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__nor2_1
XFILLER_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout194 _15151_/X vssd1 vssd1 vccd1 vccd1 _16136_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _16649_/A _16649_/B _16649_/C vssd1 vssd1 vccd1 vccd1 _16650_/Y sky130_fd_sc_hd__a21oi_1
X_13862_ _13862_/A _13964_/A _13862_/C vssd1 vssd1 vccd1 vccd1 _13862_/X sky130_fd_sc_hd__and3_2
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ _15601_/A _15601_/B vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__xor2_4
XFILLER_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12813_ _12663_/B _12665_/B _12663_/A vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__o21ba_4
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16581_ _12869_/C _17075_/A2 _16580_/X vssd1 vssd1 vccd1 vccd1 _16581_/Y sky130_fd_sc_hd__a21oi_1
X_13793_ _13793_/A _13793_/B _13793_/C vssd1 vssd1 vccd1 vccd1 _13795_/A sky130_fd_sc_hd__or3_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15532_ _15532_/A _15532_/B vssd1 vssd1 vccd1 vccd1 _15533_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12744_/A _12902_/B vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__and2_4
XFILLER_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15463_/Y sky130_fd_sc_hd__nor2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12675_ _12675_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _12676_/C sky130_fd_sc_hd__xor2_1
XFILLER_169_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17202_ _17544_/Q _17232_/B vssd1 vssd1 vccd1 vccd1 _17202_/X sky130_fd_sc_hd__and2_1
XFILLER_187_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14414_ _14414_/A _14414_/B vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11626_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _15524_/B sky130_fd_sc_hd__and2_1
XFILLER_168_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15394_ _15071_/A _11789_/X _15551_/A vssd1 vssd1 vccd1 vccd1 _15472_/B sky130_fd_sc_hd__a21oi_4
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17133_ _17133_/A vssd1 vssd1 vccd1 vccd1 _17133_/Y sky130_fd_sc_hd__inv_2
X_14345_ _14413_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _14348_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11557_ _11558_/A _11558_/B _11558_/C vssd1 vssd1 vccd1 vccd1 _11557_/X sky130_fd_sc_hd__and3_2
XFILLER_155_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17064_ _14765_/A _16644_/B _17065_/A vssd1 vssd1 vccd1 vccd1 _17064_/X sky130_fd_sc_hd__a21bo_2
X_10508_ _10509_/A _10507_/Y _10508_/C _10970_/B vssd1 vssd1 vccd1 vccd1 _10617_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ _14276_/A _14276_/B _14274_/X vssd1 vssd1 vccd1 vccd1 _14277_/B sky130_fd_sc_hd__or3b_1
X_11488_ _11487_/A _11527_/A _11444_/Y _11466_/X vssd1 vssd1 vccd1 vccd1 _11496_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_171_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16015_ _16015_/A _16114_/B _16015_/C vssd1 vssd1 vccd1 vccd1 _16015_/X sky130_fd_sc_hd__or3_1
X_13227_ _17419_/A _17417_/A _13664_/D _13551_/D vssd1 vssd1 vccd1 vccd1 _13228_/B
+ sky130_fd_sc_hd__and4_1
X_10439_ _10425_/Y _10437_/X _10453_/A _10410_/Y vssd1 vssd1 vccd1 vccd1 _10453_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_170_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _13643_/A _13908_/B vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _17381_/A _12734_/C vssd1 vssd1 vccd1 vccd1 _12110_/B sky130_fd_sc_hd__nand2_2
X_13089_ _17407_/A _13088_/B _13088_/C vssd1 vssd1 vccd1 vccd1 _13090_/B sky130_fd_sc_hd__a21o_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16917_ _16917_/A _16917_/B vssd1 vssd1 vccd1 vccd1 _16917_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16848_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16850_/B sky130_fd_sc_hd__inv_2
XFILLER_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16779_ _16699_/A _16698_/B _16698_/A vssd1 vssd1 vccd1 vccd1 _16781_/B sky130_fd_sc_hd__a21boi_1
XFILLER_92_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09320_ _09748_/B _10311_/D _10308_/B _09748_/A vssd1 vssd1 vccd1 vccd1 _09320_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09251_ _09248_/Y _09249_/X _09115_/A _09114_/Y vssd1 vssd1 vccd1 vccd1 _09251_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_90_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09182_ _09214_/A vssd1 vssd1 vccd1 vccd1 _09182_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ _08993_/C _08965_/Y _08963_/X vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__o21a_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08897_ _12088_/A _12088_/B _11867_/D _12645_/B vssd1 vssd1 vccd1 vccd1 _08900_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09518_ _09519_/B _09519_/A vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__and2b_1
X_10790_ _10901_/B _10796_/B vssd1 vssd1 vccd1 vccd1 _10860_/A sky130_fd_sc_hd__nor2_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__xnor2_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12457_/X _12458_/Y _12267_/Y _12290_/X vssd1 vssd1 vccd1 vccd1 _12481_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_166_930 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11411_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _11419_/B sky130_fd_sc_hd__xor2_4
X_12391_ _12389_/X _12390_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _14130_/A _14134_/B _13958_/C vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__nor3b_1
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11342_ _11329_/Y _11367_/A _11343_/A _11312_/Y vssd1 vssd1 vccd1 vccd1 _11349_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_181_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14061_ _13967_/A _13969_/B _13967_/B vssd1 vssd1 vccd1 vccd1 _14068_/A sky130_fd_sc_hd__o21ba_1
X_11273_ _11274_/B _11274_/C _11274_/A vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__a21o_1
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10224_ _10226_/A _10226_/B _10221_/X vssd1 vssd1 vccd1 vccd1 _10348_/C sky130_fd_sc_hd__a21oi_4
X_13012_ _13627_/S _11833_/X _11854_/C _12858_/Y vssd1 vssd1 vccd1 vccd1 _13012_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10155_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10086_ _10086_/A _10086_/B _10086_/C vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__or3_4
XFILLER_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14963_ _15175_/A _15808_/A vssd1 vssd1 vccd1 vccd1 _14963_/X sky130_fd_sc_hd__or2_4
XFILLER_12_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16702_ _16777_/B _16702_/B vssd1 vssd1 vccd1 vccd1 _16705_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13914_ _13915_/A _13915_/B _13915_/C vssd1 vssd1 vccd1 vccd1 _14021_/A sky130_fd_sc_hd__o21a_1
X_14894_ _14901_/B _15703_/A _15617_/A vssd1 vssd1 vccd1 vccd1 _15208_/D sky130_fd_sc_hd__or3_4
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16633_ _16634_/A _16634_/B vssd1 vssd1 vccd1 vccd1 _16711_/B sky130_fd_sc_hd__nor2_2
X_13845_ _13845_/A _13954_/A vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__nor2_1
X_16564_ _16564_/A _16564_/B vssd1 vssd1 vccd1 vccd1 _16564_/Y sky130_fd_sc_hd__nor2_1
X_13776_ _13776_/A _13776_/B vssd1 vssd1 vccd1 vccd1 _13778_/C sky130_fd_sc_hd__xnor2_1
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10988_ _10990_/A _10990_/B _10990_/C vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_16_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15515_ _15609_/A _15515_/B vssd1 vssd1 vccd1 vccd1 _15518_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ _12727_/A _12727_/B vssd1 vssd1 vccd1 vccd1 _12728_/B sky130_fd_sc_hd__nor2_1
X_16495_ _16495_/A vssd1 vssd1 vccd1 vccd1 _17562_/D sky130_fd_sc_hd__inv_2
XFILLER_148_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15446_ _11672_/Y _11694_/X _11693_/Y _11691_/Y vssd1 vssd1 vccd1 vccd1 _15446_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12658_ _12658_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _12660_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11609_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__or2_2
X_15377_ _15374_/X _15375_/X _15376_/Y vssd1 vssd1 vccd1 vccd1 _15377_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_117_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12589_ _12452_/A _12452_/B _12450_/X vssd1 vssd1 vccd1 vccd1 _12610_/A sky130_fd_sc_hd__a21oi_4
XFILLER_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _14867_/A _17170_/B1 _17103_/X _17115_/X vssd1 vssd1 vccd1 vccd1 _17572_/D
+ sky130_fd_sc_hd__a22oi_1
X_14328_ _14393_/B _14328_/B vssd1 vssd1 vccd1 vccd1 _14330_/C sky130_fd_sc_hd__nand2_2
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17047_ _17088_/A _17047_/B vssd1 vssd1 vccd1 vccd1 _17049_/B sky130_fd_sc_hd__nor2_1
X_14259_ _14164_/X _14186_/A _14257_/Y _14258_/X vssd1 vssd1 vccd1 vccd1 _14340_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 _17172_/Y vssd1 vssd1 vccd1 vccd1 _17270_/B1 sky130_fd_sc_hd__buf_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout919 _17322_/C1 vssd1 vssd1 vccd1 vccd1 _17372_/C1 sky130_fd_sc_hd__buf_6
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08821_/A _08821_/C vssd1 vssd1 vccd1 vccd1 _08822_/B sky130_fd_sc_hd__nor2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _09023_/A _09023_/B _12171_/B _11961_/B vssd1 vssd1 vccd1 vccd1 _08755_/A
+ sky130_fd_sc_hd__and4_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09303_ _09304_/B _09304_/A vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__and2b_2
XFILLER_94_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09165_ _09165_/A _09165_/B _09168_/B vssd1 vssd1 vccd1 vccd1 _09178_/A sky130_fd_sc_hd__or3_4
XFILLER_163_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _10542_/A _09350_/B vssd1 vssd1 vccd1 vccd1 _14981_/A sky130_fd_sc_hd__and2_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09998_ _10255_/A _10738_/D vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__nand2_4
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08949_ _08950_/A _08948_/Y _17375_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _09065_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11960_ _11960_/A _12169_/A vssd1 vssd1 vccd1 vccd1 _11961_/C sky130_fd_sc_hd__and2_1
XFILLER_45_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _10962_/A _10911_/B vssd1 vssd1 vccd1 vccd1 _10915_/A sky130_fd_sc_hd__nand2_4
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _11891_/A _11891_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11891_/Y sky130_fd_sc_hd__nor3_4
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13630_ _14734_/A _13624_/X _13629_/X vssd1 vssd1 vccd1 vccd1 _13630_/Y sky130_fd_sc_hd__a21oi_2
X_10842_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10844_/B sky130_fd_sc_hd__xnor2_4
XFILLER_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13561_ _13557_/Y _13559_/A _13443_/B _13444_/Y vssd1 vssd1 vccd1 vccd1 _13562_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10773_ _10667_/Y _10692_/X _10766_/C _11725_/A vssd1 vssd1 vccd1 vccd1 _10774_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_160_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15300_ _15233_/X _15299_/Y _15523_/A vssd1 vssd1 vccd1 vccd1 _15300_/Y sky130_fd_sc_hd__a21oi_1
X_12512_ _12344_/B _12346_/B _12344_/A vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__o21ba_2
X_16280_ _16280_/A _16280_/B vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__nor2_4
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13492_ _13607_/B _13492_/B vssd1 vssd1 vccd1 vccd1 _13494_/C sky130_fd_sc_hd__nor2_1
XFILLER_160_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15231_ _15231_/A _15231_/B vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__nand2_1
X_12443_ _12443_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__nor2_4
XFILLER_176_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15162_ _15162_/A _15162_/B vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__nand2_4
X_12374_ _12374_/A _12374_/B vssd1 vssd1 vccd1 vccd1 _12377_/B sky130_fd_sc_hd__nand2_2
XFILLER_176_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14113_ _14113_/A _14113_/B _14113_/C vssd1 vssd1 vccd1 vccd1 _14114_/B sky130_fd_sc_hd__nand3_1
XFILLER_126_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11325_ _11325_/A _11376_/A vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nand2_4
XFILLER_181_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15093_ _15093_/A _15093_/B vssd1 vssd1 vccd1 vccd1 _15170_/C sky130_fd_sc_hd__nand2_2
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14044_ _14044_/A _14044_/B vssd1 vssd1 vccd1 vccd1 _14045_/B sky130_fd_sc_hd__nor2_1
XFILLER_125_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11256_ _11255_/A _11255_/C _11255_/B vssd1 vssd1 vccd1 vccd1 _11256_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__nor2_2
XFILLER_80_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11187_ _11202_/B _11186_/B _11218_/A _11186_/D vssd1 vssd1 vccd1 vccd1 _11187_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10138_ _10138_/A _10138_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10138_/Y sky130_fd_sc_hd__nand3_2
X_15995_ _15994_/A _15993_/X _15523_/A vssd1 vssd1 vccd1 vccd1 _15995_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10069_ _10069_/A _10069_/B _10200_/A vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__or3_1
XFILLER_48_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14946_ _09350_/B _12597_/B _17139_/A _12442_/B _15062_/S0 _15095_/B vssd1 vssd1
+ vccd1 vccd1 _14947_/B sky130_fd_sc_hd__mux4_1
XFILLER_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14877_ _17614_/Q _15147_/C _17613_/Q vssd1 vssd1 vccd1 vccd1 _14877_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16616_ _16616_/A _16616_/B _16616_/C vssd1 vssd1 vccd1 vccd1 _16617_/B sky130_fd_sc_hd__nor3_2
X_13828_ _13727_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13830_/B sky130_fd_sc_hd__and2b_1
XFILLER_91_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17596_ fanout943/X _17596_/D vssd1 vssd1 vccd1 vccd1 _17596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16547_ _16547_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _16548_/B sky130_fd_sc_hd__or2_1
X_13759_ _13656_/B _13659_/B _13654_/X vssd1 vssd1 vccd1 vccd1 _13761_/B sky130_fd_sc_hd__a21oi_2
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16478_ _16478_/A _16478_/B vssd1 vssd1 vccd1 vccd1 _16478_/X sky130_fd_sc_hd__or2_4
XFILLER_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15429_ _15429_/A _15429_/B vssd1 vssd1 vccd1 vccd1 _15431_/A sky130_fd_sc_hd__xnor2_4
XFILLER_191_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09921_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__nand2_2
XFILLER_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout705 _15101_/A1 vssd1 vssd1 vccd1 vccd1 _13094_/B sky130_fd_sc_hd__buf_12
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout716 _17497_/Q vssd1 vssd1 vccd1 vccd1 _12077_/C sky130_fd_sc_hd__buf_8
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__xnor2_4
Xfanout727 _17496_/Q vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__buf_6
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout738 _17494_/Q vssd1 vssd1 vccd1 vccd1 _11859_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout749 _09428_/B vssd1 vssd1 vccd1 vccd1 _10036_/D sky130_fd_sc_hd__buf_6
X_08803_ _09025_/C _11961_/B _08772_/C _08772_/D vssd1 vssd1 vccd1 vccd1 _08804_/B
+ sky130_fd_sc_hd__a22oi_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _09930_/A vssd1 vssd1 vccd1 vccd1 _09784_/C sky130_fd_sc_hd__nor2_1
XFILLER_58_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _17608_/Q _17607_/Q vssd1 vssd1 vccd1 vccd1 _14836_/B sky130_fd_sc_hd__and2b_2
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09217_ _12488_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _09219_/C sky130_fd_sc_hd__nand2_1
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09148_ _09148_/A _09148_/B vssd1 vssd1 vccd1 vccd1 _09150_/B sky130_fd_sc_hd__xnor2_4
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_955 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09079_ _09748_/B _12088_/C _12088_/D _09748_/A vssd1 vssd1 vccd1 vccd1 _09079_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _11110_/A _11110_/B _11110_/C vssd1 vssd1 vccd1 vccd1 _11144_/A sky130_fd_sc_hd__nand3_4
XFILLER_162_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _12258_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12091_/B sky130_fd_sc_hd__nand2_4
XFILLER_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ _11041_/A _11041_/B _11041_/C vssd1 vssd1 vccd1 vccd1 _11041_/Y sky130_fd_sc_hd__nand3_4
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14800_ _15244_/B _15244_/C _15244_/A vssd1 vssd1 vccd1 vccd1 _14801_/C sky130_fd_sc_hd__o21ba_1
XTAP_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _15781_/A _15781_/B vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__and2b_1
XTAP_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _12993_/A _12993_/B _12991_/X vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__nor3b_1
XTAP_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _14731_/A _14731_/B vssd1 vssd1 vccd1 vccd1 _14731_/X sky130_fd_sc_hd__or2_1
XFILLER_40_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _12156_/A vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__clkinv_2
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ fanout938/X _17450_/D vssd1 vssd1 vccd1 vccd1 _17450_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14662_/A _14662_/B vssd1 vssd1 vccd1 vccd1 _14669_/B sky130_fd_sc_hd__xnor2_4
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__or2_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16397_/B _16580_/A2 _16733_/B1 _16399_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16401_/X sky130_fd_sc_hd__a221o_1
X_13613_ _17405_/A _16789_/A _13465_/A _13463_/A vssd1 vssd1 vccd1 vccd1 _13614_/B
+ sky130_fd_sc_hd__a31o_2
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _11115_/A _11258_/B _10911_/B _10912_/C vssd1 vssd1 vccd1 vccd1 _10827_/A
+ sky130_fd_sc_hd__and4_1
X_17381_ _17381_/A _17397_/B vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__or2_1
X_14593_ _14593_/A _14593_/B _14593_/C _14593_/D vssd1 vssd1 vccd1 vccd1 _14594_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_186_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16332_ _16245_/A _16245_/B _16248_/A vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__a21oi_2
XFILLER_158_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13544_ _13545_/A _13545_/B _13545_/C vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__a21oi_4
XFILLER_38_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10756_ _10756_/A _11165_/A vssd1 vssd1 vccd1 vccd1 _10757_/C sky130_fd_sc_hd__nor2_1
XFILLER_158_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16263_ _16262_/A _16681_/C _16262_/C vssd1 vssd1 vccd1 vccd1 _16264_/B sky130_fd_sc_hd__o21a_1
XFILLER_158_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _13476_/B _13476_/A vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__and2b_1
X_10687_ _10685_/B _10685_/C _10685_/A vssd1 vssd1 vccd1 vccd1 _10688_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15214_ _15214_/A _15494_/A vssd1 vssd1 vccd1 vccd1 _15216_/A sky130_fd_sc_hd__xnor2_4
X_12426_ _12578_/A _12576_/C vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__nand2_2
X_16194_ _16195_/A _16195_/B vssd1 vssd1 vccd1 vccd1 _16290_/A sky130_fd_sc_hd__nor2_1
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15145_ _14886_/D _15144_/X _15175_/A vssd1 vssd1 vccd1 vccd1 _15145_/X sky130_fd_sc_hd__a21o_4
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12357_ _12357_/A _12357_/B vssd1 vssd1 vccd1 vccd1 _12358_/C sky130_fd_sc_hd__xnor2_4
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__xnor2_4
XFILLER_142_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15076_ _14967_/C _14967_/D _15075_/X _14877_/Y vssd1 vssd1 vccd1 vccd1 _15077_/B
+ sky130_fd_sc_hd__o22a_1
X_12288_ _12476_/A _12286_/Y _12112_/X _12116_/A vssd1 vssd1 vccd1 vccd1 _12290_/D
+ sky130_fd_sc_hd__a211o_2
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14027_ _14027_/A _14027_/B _14025_/Y vssd1 vssd1 vccd1 vccd1 _14028_/B sky130_fd_sc_hd__or3b_1
X_11239_ _15472_/A _11370_/D vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__nand2_4
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15978_ _15980_/A _15980_/B _15980_/C vssd1 vssd1 vccd1 vccd1 _15981_/A sky130_fd_sc_hd__o21a_1
X_14929_ _14929_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__or2_4
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17579_ fanout937/X _17579_/D vssd1 vssd1 vccd1 vccd1 _17579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09002_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09002_/X sky130_fd_sc_hd__and2b_1
XFILLER_118_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_958 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09904_ _09906_/B _10035_/A _09906_/A vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__a21o_1
Xfanout502 _11115_/A vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__buf_6
Xfanout513 _15373_/C vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__buf_2
Xfanout524 _17516_/Q vssd1 vssd1 vccd1 vccd1 _10640_/C sky130_fd_sc_hd__buf_12
XFILLER_99_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout535 _11266_/A vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__buf_6
XFILLER_101_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout546 _10532_/B vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__buf_6
XFILLER_98_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09835_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__xnor2_2
Xfanout557 _14637_/A1 vssd1 vssd1 vccd1 vccd1 _13516_/S sky130_fd_sc_hd__buf_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout568 _11268_/A vssd1 vssd1 vccd1 vccd1 _10299_/C sky130_fd_sc_hd__buf_4
XFILLER_86_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout579 _14922_/S vssd1 vssd1 vccd1 vccd1 _15126_/A sky130_fd_sc_hd__buf_4
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09766_ _09776_/A _09745_/Y _09761_/A _09765_/X vssd1 vssd1 vccd1 vccd1 _09769_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08717_ _17517_/Q vssd1 vssd1 vccd1 vccd1 _17377_/A sky130_fd_sc_hd__inv_4
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09697_ _10241_/B _10392_/D _10377_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _09699_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A _10610_/B vssd1 vssd1 vccd1 vccd1 _10711_/B sky130_fd_sc_hd__xnor2_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__nor2_4
XFILLER_168_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _14982_/A _10543_/B _10434_/A _10432_/Y vssd1 vssd1 vccd1 vccd1 _10547_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13260_ _13260_/A vssd1 vssd1 vccd1 vccd1 _13261_/C sky130_fd_sc_hd__inv_2
X_10472_ _10459_/A _10459_/C _10459_/B vssd1 vssd1 vccd1 vccd1 _10472_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12211_ _11804_/Y _11807_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _12211_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _13061_/A _13063_/A _13188_/X _13190_/Y vssd1 vssd1 vccd1 vccd1 _13332_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_123_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _11937_/A _11937_/B _11936_/A vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__a21oi_4
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16950_ _16950_/A _16950_/B vssd1 vssd1 vccd1 vccd1 _16952_/C sky130_fd_sc_hd__xor2_4
X_12073_ _11860_/A _11862_/B _11860_/B vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__o21ba_1
XFILLER_2_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11024_ _11024_/A _11024_/B _11024_/C vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__or3_2
X_15901_ _15245_/X _15253_/X _15901_/S vssd1 vssd1 vccd1 vccd1 _15901_/X sky130_fd_sc_hd__mux2_1
X_16881_ _16880_/A _16935_/B _16880_/C vssd1 vssd1 vccd1 vccd1 _16882_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _15832_/A _15832_/B vssd1 vssd1 vccd1 vccd1 _15834_/B sky130_fd_sc_hd__xnor2_4
XFILLER_65_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _15764_/A _15764_/B _15764_/C vssd1 vssd1 vccd1 vccd1 _15868_/B sky130_fd_sc_hd__a21oi_4
XTAP_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ _13112_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _12975_/X sky130_fd_sc_hd__and2_1
XTAP_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14714_ _14713_/A _14713_/B _14713_/C vssd1 vssd1 vccd1 vccd1 _14715_/B sky130_fd_sc_hd__a21o_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17502_ fanout932/X _17502_/D vssd1 vssd1 vccd1 vccd1 _17502_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11926_ _11932_/A _12752_/B _09001_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _11937_/A
+ sky130_fd_sc_hd__a31o_4
X_15694_ _15595_/A _15599_/A _15786_/A _15693_/Y vssd1 vssd1 vccd1 vccd1 _15786_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17433_ input61/X _17477_/D _17433_/S vssd1 vssd1 vccd1 vccd1 _17610_/D sky130_fd_sc_hd__mux2_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14645_ _14645_/A _14678_/B vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11857_ _11785_/X _11786_/Y _11856_/X vssd1 vssd1 vccd1 vccd1 _17576_/D sky130_fd_sc_hd__o21ai_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10808_ _10808_/A _10808_/B vssd1 vssd1 vccd1 vccd1 _10814_/A sky130_fd_sc_hd__xnor2_4
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17364_ input36/X _17384_/A2 _17363_/Y _17428_/B vssd1 vssd1 vccd1 vccd1 _17510_/D
+ sky130_fd_sc_hd__o211a_1
X_14576_ _14577_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__nor2_1
X_11788_ _16108_/C _16317_/A vssd1 vssd1 vccd1 vccd1 _14888_/B sky130_fd_sc_hd__or2_4
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16315_ _16315_/A _16315_/B _16315_/C _17038_/C vssd1 vssd1 vccd1 vccd1 _16316_/B
+ sky130_fd_sc_hd__or4_4
X_13527_ _13637_/B _13527_/B _13527_/C vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__and3_1
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10739_ _10739_/A _11018_/A vssd1 vssd1 vccd1 vccd1 _10747_/A sky130_fd_sc_hd__nor2_4
X_17295_ input25/X _17362_/D input28/X _17428_/C vssd1 vssd1 vccd1 vccd1 _17295_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_146_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16246_ _16246_/A _16589_/B _16246_/C vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__and3_1
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13458_ _13459_/A _13459_/B vssd1 vssd1 vccd1 vccd1 _13576_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ _12409_/A _12561_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__nor2_4
X_16177_ _16177_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _16179_/B sky130_fd_sc_hd__xnor2_1
Xoutput105 _17463_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13389_ _16922_/A _13387_/Y _13388_/X _13274_/Y _13277_/X vssd1 vssd1 vccd1 vccd1
+ _17586_/D sky130_fd_sc_hd__a32o_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15128_ _15381_/A _15463_/A _15541_/A _15624_/A _14942_/A _10993_/C vssd1 vssd1 vccd1
+ vccd1 _15131_/B sky130_fd_sc_hd__mux4_1
XFILLER_86_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15059_ _15059_/A _15059_/B vssd1 vssd1 vccd1 vccd1 _15059_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09621_/C sky130_fd_sc_hd__and2_2
X_09551_ _09552_/A _09550_/Y _10366_/A _10490_/C vssd1 vssd1 vccd1 vccd1 _09696_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09482_ _09476_/Y _09480_/X _09460_/X _09461_/Y vssd1 vssd1 vccd1 vccd1 _09484_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout310 _17611_/Q vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__buf_4
Xfanout321 _17541_/Q vssd1 vssd1 vccd1 vccd1 _14832_/A sky130_fd_sc_hd__buf_8
Xfanout332 _12620_/A vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__clkbuf_16
Xfanout343 _12657_/B vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__buf_6
XFILLER_28_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout354 _12659_/A vssd1 vssd1 vccd1 vccd1 _14226_/A sky130_fd_sc_hd__buf_12
Xfanout365 _12487_/B vssd1 vssd1 vccd1 vccd1 _11953_/B sky130_fd_sc_hd__buf_8
XFILLER_8_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout376 _14168_/A vssd1 vssd1 vccd1 vccd1 _14387_/A sky130_fd_sc_hd__clkbuf_8
X_09818_ _09828_/A _09817_/B _09814_/X vssd1 vssd1 vccd1 vccd1 _09819_/C sky130_fd_sc_hd__a21oi_1
Xfanout387 _17532_/Q vssd1 vssd1 vccd1 vccd1 _16723_/A sky130_fd_sc_hd__buf_6
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout398 _09838_/A vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__buf_4
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09749_ _09748_/B _10753_/B _09892_/C _09748_/A vssd1 vssd1 vccd1 vccd1 _09749_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12761_/A _12761_/B _12761_/C vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__o21a_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/A _11711_/B vssd1 vssd1 vccd1 vccd1 _11713_/B sky130_fd_sc_hd__xnor2_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A _12691_/B vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__or2_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _14431_/B sky130_fd_sc_hd__and2_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _15305_/C _11605_/B _11610_/B _11605_/D vssd1 vssd1 vccd1 vccd1 _11644_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14361_ _14361_/A _14440_/A vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__or2_1
XFILLER_168_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ _11534_/B _11530_/B _11530_/C vssd1 vssd1 vccd1 vccd1 _11574_/C sky130_fd_sc_hd__a21oi_4
XFILLER_35_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16100_ _16203_/A _16100_/B vssd1 vssd1 vccd1 vccd1 _16100_/Y sky130_fd_sc_hd__nor2_1
Xinput18 i_wb_addr[23] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
X_13312_ _13312_/A _13312_/B _13312_/C vssd1 vssd1 vccd1 vccd1 _13317_/B sky130_fd_sc_hd__or3_4
X_17080_ _17065_/A _17170_/B1 _17063_/Y _17079_/X vssd1 vssd1 vccd1 vccd1 _17571_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput29 i_wb_addr[4] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_4
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__xnor2_4
X_14292_ _14676_/A _14360_/C vssd1 vssd1 vccd1 vccd1 _14294_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16031_ _16226_/B _16743_/C _16136_/C vssd1 vssd1 vccd1 vccd1 _16032_/B sky130_fd_sc_hd__and3_1
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _13243_/A _13243_/B vssd1 vssd1 vccd1 vccd1 _13244_/C sky130_fd_sc_hd__or2_2
XFILLER_182_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10455_ _10564_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__or2_2
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13174_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13176_/B sky130_fd_sc_hd__xnor2_4
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _10385_/A _10385_/Y _10262_/X _10357_/Y vssd1 vssd1 vccd1 vccd1 _10405_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_184_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12125_ _11939_/A _11939_/B _11940_/X vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__o21ba_4
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16933_ _16933_/A _16989_/A vssd1 vssd1 vccd1 vccd1 _16933_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12056_ _12049_/Y _12051_/Y _12053_/Y _12055_/Y _12390_/S _15312_/S vssd1 vssd1 vccd1
+ vccd1 _12056_/X sky130_fd_sc_hd__mux4_2
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11007_ _11006_/B _10957_/D _11097_/D _11006_/A vssd1 vssd1 vccd1 vccd1 _11007_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16864_ _16864_/A _16864_/B vssd1 vssd1 vccd1 vccd1 _16865_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15815_ _15815_/A vssd1 vssd1 vccd1 vccd1 _17555_/D sky130_fd_sc_hd__inv_2
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16795_ _16795_/A _16795_/B vssd1 vssd1 vccd1 vccd1 _16795_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_93_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15746_ _16055_/A _16681_/C vssd1 vssd1 vccd1 vccd1 _15746_/X sky130_fd_sc_hd__or2_4
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _12959_/A _12959_/B vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__or2_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11909_ _11909_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _11911_/C sky130_fd_sc_hd__or2_2
X_15677_ _15572_/Y _15583_/Y _15674_/X _15676_/A vssd1 vssd1 vccd1 vccd1 _15772_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12889_ _13298_/A _13908_/B _13903_/B _13658_/A vssd1 vssd1 vccd1 vccd1 _12889_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14628_ _14638_/A _14628_/B vssd1 vssd1 vccd1 vccd1 _14633_/A sky130_fd_sc_hd__and2_2
XFILLER_60_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17416_ input54/X _17426_/A2 _17415_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17536_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ input53/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17347_/X sky130_fd_sc_hd__or3_1
X_14559_ _14492_/A _14492_/B _14495_/A vssd1 vssd1 vccd1 vccd1 _14560_/B sky130_fd_sc_hd__o21ba_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _17460_/Q _17293_/A2 _17276_/X _17277_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17460_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16229_ _16229_/A _16229_/B vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__xor2_4
XFILLER_134_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08982_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09603_ _09603_/A _09603_/B vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__nand2_2
XFILLER_58_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09534_ _09531_/X _09540_/A _12005_/B _09397_/X vssd1 vssd1 vccd1 vccd1 _09536_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _09748_/B _10308_/B _10545_/D _09748_/A vssd1 vssd1 vccd1 vccd1 _09465_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09396_ _09343_/X _09392_/B _12005_/A _09395_/X vssd1 vssd1 vccd1 vccd1 _12005_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10240_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10261_/B sky130_fd_sc_hd__nand2_2
XFILLER_191_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _14789_/A _10171_/B _10659_/D _10755_/D vssd1 vssd1 vccd1 vccd1 _10288_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout140 _16281_/A vssd1 vssd1 vccd1 vccd1 _15774_/A sky130_fd_sc_hd__buf_8
Xfanout151 _15059_/A vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__buf_4
XFILLER_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout162 _17361_/Y vssd1 vssd1 vccd1 vccd1 _17419_/B sky130_fd_sc_hd__buf_4
X_13930_ _13930_/A _13930_/B vssd1 vssd1 vccd1 vccd1 _13932_/B sky130_fd_sc_hd__nor2_2
Xfanout173 _15749_/B vssd1 vssd1 vccd1 vccd1 _16352_/B sky130_fd_sc_hd__buf_8
Xfanout184 _15956_/B vssd1 vssd1 vccd1 vccd1 _16814_/A sky130_fd_sc_hd__buf_4
Xfanout195 _15151_/X vssd1 vssd1 vccd1 vccd1 _16317_/B sky130_fd_sc_hd__clkbuf_4
X_13861_ _13861_/A _13861_/B _13861_/C vssd1 vssd1 vccd1 vccd1 _13862_/C sky130_fd_sc_hd__nand3_1
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15600_ _15601_/A _15601_/B vssd1 vssd1 vccd1 vccd1 _15600_/Y sky130_fd_sc_hd__nor2_2
X_12812_ _12812_/A _12812_/B vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__xor2_4
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16580_ _16576_/B _16580_/A2 _16733_/B1 _16571_/A _17074_/C1 vssd1 vssd1 vccd1 vccd1
+ _16580_/X sky130_fd_sc_hd__a221o_1
X_13792_ _13792_/A _13792_/B vssd1 vssd1 vccd1 vccd1 _13793_/C sky130_fd_sc_hd__xnor2_1
XFILLER_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15531_ _15529_/Y _15620_/A vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__and2b_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12902_/A _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _12902_/B sky130_fd_sc_hd__nand3_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15462_ _15458_/Y _15459_/Y _15461_/Y vssd1 vssd1 vccd1 vccd1 _15462_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12674_ _12675_/B _12675_/A vssd1 vssd1 vccd1 vccd1 _12674_/Y sky130_fd_sc_hd__nand2b_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17201_ _17576_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17201_/X sky130_fd_sc_hd__a21o_1
XFILLER_187_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14413_ _14413_/A _14413_/B _14413_/C vssd1 vssd1 vccd1 vccd1 _14414_/B sky130_fd_sc_hd__nor3_1
X_11625_ _11617_/B _11617_/C _11617_/A vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__o21ai_2
XFILLER_169_983 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15393_ _16136_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15396_/B sky130_fd_sc_hd__nand2_2
X_17132_ _17134_/A _17134_/C _17134_/B vssd1 vssd1 vccd1 vccd1 _17133_/A sky130_fd_sc_hd__a21o_1
X_14344_ _14344_/A _14344_/B _14344_/C vssd1 vssd1 vccd1 vccd1 _14345_/B sky130_fd_sc_hd__nor3_1
XFILLER_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11556_ _11512_/A _11512_/C _11512_/B vssd1 vssd1 vccd1 vccd1 _11558_/C sky130_fd_sc_hd__a21o_1
XFILLER_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17063_ _17063_/A _17063_/B vssd1 vssd1 vccd1 vccd1 _17063_/Y sky130_fd_sc_hd__nor2_1
X_10507_ _10963_/B _10971_/B _10920_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _10507_/Y
+ sky130_fd_sc_hd__a22oi_2
X_14275_ _14276_/A _14276_/B _14274_/X vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__o21ba_1
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11487_ _11487_/A _11487_/B _11485_/X vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__nor3b_4
XFILLER_171_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16014_ _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16015_/C sky130_fd_sc_hd__nor2_1
X_13226_ _17417_/A _13664_/D _13551_/D _17419_/A vssd1 vssd1 vccd1 vccd1 _13228_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10438_ _10453_/A _10410_/Y _10425_/Y _10437_/X vssd1 vssd1 vccd1 vccd1 _10440_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ _13157_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__nor2_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10484_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__nand2_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _12108_/A _12108_/B vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__nor2_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _17407_/A _13088_/B _13088_/C vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__nand3_2
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16916_ _16916_/A _16916_/B vssd1 vssd1 vccd1 vccd1 _16917_/B sky130_fd_sc_hd__xnor2_1
X_12039_ _14848_/B _17304_/A1 _12060_/S vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16847_ _16909_/A _16847_/B vssd1 vssd1 vccd1 vccd1 _16848_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16778_ _16846_/A _16778_/B vssd1 vssd1 vccd1 vccd1 _16781_/A sky130_fd_sc_hd__or2_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15729_ _15730_/A _15730_/B vssd1 vssd1 vccd1 vccd1 _15827_/A sky130_fd_sc_hd__nand2_4
XFILLER_34_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _09115_/A _09114_/Y _09248_/Y _09249_/X vssd1 vssd1 vccd1 vccd1 _09250_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09181_ _09179_/A _09346_/A _09155_/Y _09156_/X vssd1 vssd1 vccd1 vccd1 _09214_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08965_ _12845_/S _12592_/C vssd1 vssd1 vccd1 vccd1 _08965_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08896_ _12256_/B _12645_/B vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09517_ _09517_/A _09636_/A vssd1 vssd1 vccd1 vccd1 _09519_/B sky130_fd_sc_hd__nor2_1
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09449_/B _09449_/A vssd1 vssd1 vccd1 vccd1 _09448_/X sky130_fd_sc_hd__and2b_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _09379_/A _09513_/A vssd1 vssd1 vccd1 vccd1 _09381_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11410_ _11411_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _11410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12390_ _12026_/Y _12031_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11341_ _11341_/A _11341_/B _11341_/C vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__and3_4
XFILLER_180_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14060_ _14060_/A _14060_/B vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__xnor2_1
X_11272_ _11274_/B _11274_/C _11274_/A vssd1 vssd1 vccd1 vccd1 _11272_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _16922_/A _13009_/Y _13138_/B _12860_/Y _12867_/X vssd1 vssd1 vccd1 vccd1
+ _17583_/D sky130_fd_sc_hd__a32o_1
X_10223_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10226_/B sky130_fd_sc_hd__xnor2_4
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10154_ _10137_/X _10138_/Y _10149_/A _10152_/X vssd1 vssd1 vccd1 vccd1 _10155_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14962_ _15175_/A _15808_/A vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__nor2_1
X_10085_ _10059_/A _10059_/B _10059_/C vssd1 vssd1 vccd1 vccd1 _10086_/C sky130_fd_sc_hd__o21a_1
XFILLER_43_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16701_ _16701_/A _16701_/B vssd1 vssd1 vccd1 vccd1 _16702_/B sky130_fd_sc_hd__nand2_1
X_13913_ _14013_/B _13913_/B vssd1 vssd1 vccd1 vccd1 _13915_/C sky130_fd_sc_hd__and2_1
XFILLER_47_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14893_ _14901_/B _15703_/A vssd1 vssd1 vccd1 vccd1 _14967_/C sky130_fd_sc_hd__or2_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _13844_/A _13844_/B _14181_/B _13844_/D vssd1 vssd1 vccd1 vccd1 _13954_/A
+ sky130_fd_sc_hd__and4_1
X_16632_ _16543_/A _16543_/B _16544_/X vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__a21oi_2
XFILLER_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16563_ _16563_/A _16563_/B vssd1 vssd1 vccd1 vccd1 _16564_/B sky130_fd_sc_hd__nor2_1
X_13775_ _14226_/A _14213_/D vssd1 vssd1 vccd1 vccd1 _13776_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10987_ _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _10990_/C sky130_fd_sc_hd__xnor2_4
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12726_ _12727_/A _12727_/B vssd1 vssd1 vccd1 vccd1 _12886_/B sky130_fd_sc_hd__and2_2
X_15514_ _15514_/A _15514_/B _15514_/C vssd1 vssd1 vccd1 vccd1 _15515_/B sky130_fd_sc_hd__and3_1
X_16494_ _16475_/X _16478_/X _16493_/X _16806_/A2 _16480_/A vssd1 vssd1 vccd1 vccd1
+ _16495_/A sky130_fd_sc_hd__a32o_1
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15445_ _15442_/Y _15443_/X _15444_/Y vssd1 vssd1 vccd1 vccd1 _15445_/X sky130_fd_sc_hd__a21o_1
X_12657_ _12657_/A _12657_/B _13194_/D _13067_/D vssd1 vssd1 vccd1 vccd1 _12658_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_169_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _11607_/A _11607_/C _11607_/B vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__a21o_1
XFILLER_191_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15376_ _15374_/X _15375_/X _15309_/B vssd1 vssd1 vccd1 vccd1 _15376_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ _12588_/A _12588_/B _12588_/C vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__and3_2
XFILLER_117_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14327_ _14326_/A _14554_/B _14326_/C vssd1 vssd1 vccd1 vccd1 _14328_/B sky130_fd_sc_hd__a21o_1
X_17115_ _17063_/A _17096_/Y _17097_/X _17114_/X vssd1 vssd1 vccd1 vccd1 _17115_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11539_ _11539_/A _11539_/B _11538_/X vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__nor3b_4
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17046_ _17046_/A _17046_/B _17046_/C vssd1 vssd1 vccd1 vccd1 _17047_/B sky130_fd_sc_hd__nor3_1
X_14258_ _14258_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__or2_1
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13209_ _14771_/A _14050_/D vssd1 vssd1 vccd1 vccd1 _13211_/C sky130_fd_sc_hd__nand2_1
X_14189_ _14268_/A _14189_/B vssd1 vssd1 vccd1 vccd1 _14190_/B sky130_fd_sc_hd__nor2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout909 _17266_/A2 vssd1 vssd1 vccd1 vccd1 _17233_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_98_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08750_/B vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__xnor2_4
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _09302_/A _09443_/A vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09233_ _12174_/A _12174_/B _12129_/B _12127_/C vssd1 vssd1 vccd1 vccd1 _09234_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_181_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09164_ _09164_/A _09354_/A vssd1 vssd1 vccd1 vccd1 _09168_/B sky130_fd_sc_hd__nor2_4
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09095_ _09095_/A _09095_/B vssd1 vssd1 vccd1 vccd1 _09103_/A sky130_fd_sc_hd__nor2_2
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09997_ _10254_/A _10254_/B _10736_/C _10392_/D vssd1 vssd1 vccd1 vccd1 _10000_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08948_ _12592_/B _12090_/B _12565_/C _11895_/A vssd1 vssd1 vccd1 vccd1 _08948_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_85_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08879_ _09023_/A _09023_/B _09414_/C _09509_/B vssd1 vssd1 vccd1 vccd1 _08882_/A
+ sky130_fd_sc_hd__and4_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _11107_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11074_/A sky130_fd_sc_hd__nand2_4
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11890_ _11891_/A _11891_/B _11891_/C vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__o21a_2
XFILLER_45_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10841_ _10841_/A _10841_/B vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__nor2_4
XFILLER_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _13443_/B _13444_/Y _13557_/Y _13559_/A vssd1 vssd1 vccd1 vccd1 _13562_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_53_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _10777_/A _10772_/B vssd1 vssd1 vccd1 vccd1 _10774_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12511_ _12511_/A _12511_/B vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__xor2_4
XFILLER_160_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ _13607_/A _13490_/B _13490_/C _13490_/D vssd1 vssd1 vccd1 vccd1 _13492_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15230_ _15230_/A _15230_/B vssd1 vssd1 vccd1 vccd1 _15231_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _12442_/A _12442_/B _12442_/C vssd1 vssd1 vccd1 vccd1 _12616_/B sky130_fd_sc_hd__and3_2
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15162_/B sky130_fd_sc_hd__nand2_1
XFILLER_153_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _12373_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__xnor2_2
XFILLER_181_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14112_ _14113_/A _14113_/B _14113_/C vssd1 vssd1 vccd1 vccd1 _14202_/A sky130_fd_sc_hd__a21o_1
XFILLER_4_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _11553_/B _11518_/C _11325_/A _11324_/D vssd1 vssd1 vccd1 vccd1 _11376_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_176_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15092_ _15170_/A _15170_/B vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _14043_/A _14043_/B vssd1 vssd1 vccd1 vccd1 _14134_/B sky130_fd_sc_hd__xnor2_4
XFILLER_125_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11255_ _11255_/A _11255_/B _11255_/C vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__or3_4
XFILLER_140_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10206_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__and2b_2
X_11186_ _11202_/B _11186_/B _11218_/A _11186_/D vssd1 vssd1 vccd1 vccd1 _11218_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_80_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10137_ _10138_/A _10138_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10137_/X sky130_fd_sc_hd__a21o_4
X_15994_ _15994_/A _15994_/B vssd1 vssd1 vccd1 vccd1 _15994_/X sky130_fd_sc_hd__and2_2
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10068_ _10069_/B _10200_/A _10069_/A vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__o21ai_4
X_14945_ _14924_/A _11853_/Y _14841_/B _14944_/Y vssd1 vssd1 vccd1 vccd1 _14945_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14876_ _15396_/A _14888_/C _14876_/C _14876_/D vssd1 vssd1 vccd1 vccd1 _14876_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_78_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16615_ _16616_/A _16616_/B _16616_/C vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__o21a_2
X_13827_ _13827_/A _13827_/B vssd1 vssd1 vccd1 vccd1 _13936_/B sky130_fd_sc_hd__xor2_2
X_17595_ fanout941/X _17595_/D vssd1 vssd1 vccd1 vccd1 _17595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16546_ _16547_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _16630_/B sky130_fd_sc_hd__nand2_2
X_13758_ _13862_/A _13758_/B vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__or2_1
XFILLER_176_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ _13837_/A _12709_/B vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__or2_4
X_16477_ _11200_/Y _11229_/Y _16389_/C _16207_/B vssd1 vssd1 vccd1 vccd1 _16478_/B
+ sky130_fd_sc_hd__a31o_1
X_13689_ _14771_/A _16789_/A vssd1 vssd1 vccd1 vccd1 _16796_/A sky130_fd_sc_hd__nand2_4
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15428_ _15428_/A _15428_/B _15429_/B vssd1 vssd1 vccd1 vccd1 _15428_/X sky130_fd_sc_hd__and3_1
XFILLER_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15359_ _15359_/A _15359_/B vssd1 vssd1 vccd1 vccd1 _15362_/A sky130_fd_sc_hd__xor2_4
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _09920_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__and2_1
XFILLER_171_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17029_ _17140_/A _17029_/B _17029_/C vssd1 vssd1 vccd1 vccd1 _17033_/B sky130_fd_sc_hd__or3_1
XFILLER_131_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout706 _10308_/B vssd1 vssd1 vccd1 vccd1 _10543_/B sky130_fd_sc_hd__buf_4
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09851_ _09845_/B _09847_/B _09845_/A vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__o21ba_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout717 _14050_/D vssd1 vssd1 vccd1 vccd1 _13450_/D sky130_fd_sc_hd__clkbuf_16
Xfanout728 _12795_/B vssd1 vssd1 vccd1 vccd1 _11867_/D sky130_fd_sc_hd__buf_8
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 _13229_/B vssd1 vssd1 vccd1 vccd1 _13764_/D sky130_fd_sc_hd__buf_8
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__xnor2_2
XFILLER_86_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09783_/A _09781_/Y _09928_/C _09926_/B vssd1 vssd1 vccd1 vccd1 _09930_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08733_ _17476_/D _17477_/D vssd1 vssd1 vccd1 vccd1 _08733_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _11953_/A _11953_/B _12338_/C _12338_/D vssd1 vssd1 vccd1 vccd1 _11958_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_148_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09147_ _09148_/A _09147_/B _09231_/B vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__or3_2
XFILLER_147_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09078_ _12592_/A _09748_/B _12088_/C _12565_/D vssd1 vssd1 vccd1 vccd1 _09081_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_136_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11040_ _11046_/A _11040_/B vssd1 vssd1 vccd1 vccd1 _11041_/C sky130_fd_sc_hd__xnor2_4
XFILLER_131_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _12991_/A _12991_/B vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__or2_1
XFILLER_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730_ _14731_/A _14731_/B vssd1 vssd1 vccd1 vccd1 _14730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11942_ _08868_/X _08873_/C _11940_/X _11941_/Y vssd1 vssd1 vccd1 vccd1 _12156_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14661_ _14661_/A _14662_/A vssd1 vssd1 vccd1 vccd1 _14698_/B sky130_fd_sc_hd__nand2_1
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__nand2_2
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13612_/A _13612_/B vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__nor2_4
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16400_ _16652_/A _16400_/B _16400_/C vssd1 vssd1 vccd1 vccd1 _16404_/A sky130_fd_sc_hd__or3_1
XFILLER_189_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _11260_/C _10962_/B vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__nand2_4
X_14592_ _14593_/B _14593_/C _14593_/D _14593_/A vssd1 vssd1 vccd1 vccd1 _14594_/A
+ sky130_fd_sc_hd__a22oi_4
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17380_ input66/X _17396_/A2 _17379_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17518_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16331_ _16331_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__xor2_1
X_13543_ _13543_/A _13543_/B vssd1 vssd1 vccd1 vccd1 _13545_/C sky130_fd_sc_hd__xnor2_4
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ _10756_/A _10754_/Y _14794_/A _10755_/D vssd1 vssd1 vccd1 vccd1 _11165_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _16262_/A _16681_/C _16262_/C vssd1 vssd1 vccd1 vccd1 _16358_/B sky130_fd_sc_hd__nor3_2
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13474_ _13353_/A _13355_/B _13353_/B vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__o21ba_1
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10686_ _10579_/B _10584_/X _10685_/B _10688_/A vssd1 vssd1 vccd1 vccd1 _11768_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15213_ _15660_/A _15918_/A _15213_/C vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__and3_1
X_12425_ _12425_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__nor2_1
X_16193_ _16089_/A _16089_/B _16081_/A vssd1 vssd1 vccd1 vccd1 _16195_/B sky130_fd_sc_hd__o21a_1
XFILLER_127_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ _11790_/X _14877_/Y _15270_/B _15143_/C _15143_/A vssd1 vssd1 vccd1 vccd1
+ _15144_/X sky130_fd_sc_hd__a2111o_1
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12356_ _12357_/B _12357_/A vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__and2b_1
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__nand2_4
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15075_ _15204_/A _15147_/C vssd1 vssd1 vccd1 vccd1 _15075_/X sky130_fd_sc_hd__and2_1
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12287_ _12112_/X _12116_/A _12476_/A _12286_/Y vssd1 vssd1 vccd1 vccd1 _12476_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_153_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14026_ _14027_/A _14027_/B _14025_/Y vssd1 vssd1 vccd1 vccd1 _14119_/B sky130_fd_sc_hd__o21ba_1
X_11238_ _11238_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11249_/A sky130_fd_sc_hd__xor2_4
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11169_ _11168_/A _11168_/B _11167_/X vssd1 vssd1 vccd1 vccd1 _11169_/X sky130_fd_sc_hd__o21ba_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15977_ _16165_/A _16165_/B _15850_/A _15848_/A vssd1 vssd1 vccd1 vccd1 _15980_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14928_ _14929_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14928_/Y sky130_fd_sc_hd__nor2_2
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _16298_/A _14859_/B _16115_/B vssd1 vssd1 vccd1 vccd1 _16399_/B sky130_fd_sc_hd__and3_1
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_283 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17578_ fanout936/X _17578_/D vssd1 vssd1 vccd1 vccd1 _17578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16529_ _16454_/A _16454_/B _16452_/Y vssd1 vssd1 vccd1 vccd1 _16545_/A sky130_fd_sc_hd__a21bo_1
XFILLER_176_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09001_ _09001_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _09003_/B sky130_fd_sc_hd__xnor2_4
XFILLER_192_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _10034_/A _10042_/A _10034_/C vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__o21ai_2
XFILLER_63_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout503 _11115_/A vssd1 vssd1 vccd1 vccd1 _11314_/A sky130_fd_sc_hd__buf_6
Xfanout514 _17517_/Q vssd1 vssd1 vccd1 vccd1 _15373_/C sky130_fd_sc_hd__buf_6
Xfanout525 _09470_/A vssd1 vssd1 vccd1 vccd1 _17373_/A sky130_fd_sc_hd__buf_6
Xfanout536 _11322_/A vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__buf_6
XFILLER_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09834_ _09866_/A _09866_/B vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__nand2_1
XFILLER_63_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout547 _10532_/B vssd1 vssd1 vccd1 vccd1 _16012_/S sky130_fd_sc_hd__buf_6
XFILLER_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout558 _13390_/S vssd1 vssd1 vccd1 vccd1 _13627_/S sky130_fd_sc_hd__buf_6
XFILLER_59_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout569 _11553_/B vssd1 vssd1 vccd1 vccd1 _11124_/C sky130_fd_sc_hd__buf_6
XFILLER_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A _09765_/B _09765_/C vssd1 vssd1 vccd1 vccd1 _09765_/X sky130_fd_sc_hd__and3_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09696_ _09696_/A _09696_/B _09703_/B vssd1 vssd1 vccd1 vccd1 _09718_/B sky130_fd_sc_hd__or3_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _10540_/A _10540_/B _10540_/C vssd1 vssd1 vccd1 vccd1 _10550_/B sky130_fd_sc_hd__nand3_2
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10463_/A _10461_/X _10454_/A _10455_/X vssd1 vssd1 vccd1 vccd1 _10471_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ _12374_/B _12210_/B vssd1 vssd1 vccd1 vccd1 _12210_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_182_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13190_ _13189_/A _13189_/B _13189_/C vssd1 vssd1 vccd1 vccd1 _13190_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_157_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12141_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12143_/A sky130_fd_sc_hd__xnor2_4
XFILLER_151_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ _12239_/B _12072_/B vssd1 vssd1 vccd1 vccd1 _12075_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11023_ _11024_/A _11024_/B _11024_/C vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__o21ai_4
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15900_ _09424_/X _17075_/A2 _15899_/X vssd1 vssd1 vccd1 vccd1 _15900_/Y sky130_fd_sc_hd__a21oi_1
X_16880_ _16880_/A _16935_/B _16880_/C vssd1 vssd1 vccd1 vccd1 _16882_/A sky130_fd_sc_hd__and3_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15831_ _15829_/X _15831_/B vssd1 vssd1 vccd1 vccd1 _15832_/B sky130_fd_sc_hd__and2b_2
XTAP_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _15762_/A _15762_/B vssd1 vssd1 vccd1 vccd1 _15764_/C sky130_fd_sc_hd__xnor2_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12974_ _12974_/A _12974_/B vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__nand2_1
XTAP_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17501_ fanout932/X _17501_/D vssd1 vssd1 vccd1 vccd1 _17501_/Q sky130_fd_sc_hd__dfxtp_1
X_14713_ _14713_/A _14713_/B _14713_/C vssd1 vssd1 vccd1 vccd1 _14742_/A sky130_fd_sc_hd__nand3_2
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11925_ _12179_/B _11925_/B vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _15779_/B _15691_/Y _15591_/A _15600_/Y vssd1 vssd1 vccd1 vccd1 _15693_/Y
+ sky130_fd_sc_hd__a211oi_4
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17432_ input58/X _17476_/D _17433_/S vssd1 vssd1 vccd1 vccd1 _17609_/D sky130_fd_sc_hd__mux2_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14644_ _14676_/A _14708_/D _14644_/C vssd1 vssd1 vccd1 vccd1 _14678_/B sky130_fd_sc_hd__and3_2
X_11856_ _11849_/A _11845_/X _13625_/B _11855_/X vssd1 vssd1 vccd1 vccd1 _11856_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _10808_/B sky130_fd_sc_hd__nor2_2
X_14575_ _14624_/A _14575_/B vssd1 vssd1 vccd1 vccd1 _14577_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17363_ _17363_/A _17377_/B vssd1 vssd1 vccd1 vccd1 _17363_/Y sky130_fd_sc_hd__nand2_1
X_11787_ _15396_/A _15373_/C vssd1 vssd1 vccd1 vccd1 _14888_/A sky130_fd_sc_hd__or2_4
X_16314_ _15647_/A _17119_/C _16695_/B _16226_/C vssd1 vssd1 vccd1 vccd1 _16316_/A
+ sky130_fd_sc_hd__a22o_1
X_13526_ _13526_/A _13526_/B vssd1 vssd1 vccd1 vccd1 _13527_/C sky130_fd_sc_hd__nand2_1
X_10738_ _10739_/A _10737_/Y _11260_/C _10738_/D vssd1 vssd1 vccd1 vccd1 _11018_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_185_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17294_ input35/X input68/X input69/X vssd1 vssd1 vccd1 vccd1 _17362_/D sky130_fd_sc_hd__nand3_4
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16245_ _16245_/A _16245_/B vssd1 vssd1 vccd1 vccd1 _16246_/C sky130_fd_sc_hd__xor2_1
X_13457_ _13457_/A _13576_/A vssd1 vssd1 vccd1 vccd1 _13459_/B sky130_fd_sc_hd__and2_1
X_10669_ _10669_/A _10669_/B _10661_/A vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__or3b_4
X_12408_ _17401_/A _13966_/D _12408_/C vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__and3_2
XFILLER_173_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16176_ _16177_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _16279_/B sky130_fd_sc_hd__and2b_1
X_13388_ _13508_/B _13388_/B vssd1 vssd1 vccd1 vccd1 _13388_/X sky130_fd_sc_hd__or2_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput106 _17436_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_182_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12339_ _12339_/A _12339_/B vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__nor2_1
X_15127_ _15126_/A _15125_/Y _15126_/Y vssd1 vssd1 vccd1 vccd1 _15711_/B sky130_fd_sc_hd__o21ai_1
XFILLER_154_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15058_ _15624_/A _15709_/A _15811_/A _09712_/B _15062_/S0 _12214_/A vssd1 vssd1
+ vccd1 vccd1 _15059_/B sky130_fd_sc_hd__mux4_1
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14009_ _14008_/A _14089_/B _14008_/C vssd1 vssd1 vccd1 vccd1 _14010_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09550_ _10235_/A _10491_/B _10490_/D _10236_/A vssd1 vssd1 vccd1 vccd1 _09550_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09481_ _09460_/X _09461_/Y _09476_/Y _09480_/X vssd1 vssd1 vccd1 vccd1 _09484_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_64_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout300 _15806_/B1 vssd1 vssd1 vccd1 vccd1 _17371_/A sky130_fd_sc_hd__buf_4
Xfanout311 _17610_/Q vssd1 vssd1 vccd1 vccd1 _17477_/D sky130_fd_sc_hd__buf_8
XFILLER_87_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout322 _17540_/Q vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__buf_6
XFILLER_114_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout333 _12620_/A vssd1 vssd1 vccd1 vccd1 _17421_/A sky130_fd_sc_hd__buf_8
XFILLER_99_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout344 _12657_/B vssd1 vssd1 vccd1 vccd1 _09172_/A sky130_fd_sc_hd__buf_2
XFILLER_28_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout355 _12659_/A vssd1 vssd1 vccd1 vccd1 _17415_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout366 _12487_/B vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__buf_4
XFILLER_87_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout377 _14771_/A vssd1 vssd1 vccd1 vccd1 _14168_/A sky130_fd_sc_hd__buf_4
X_09817_ _09814_/X _09817_/B vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__and2b_1
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout388 _12500_/A vssd1 vssd1 vccd1 vccd1 _12800_/A sky130_fd_sc_hd__buf_8
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout399 _17530_/Q vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__buf_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09748_ _09748_/A _09748_/B _10753_/B _09892_/C vssd1 vssd1 vccd1 vccd1 _09751_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_185_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__nor2_2
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _15997_/A _15997_/B _16105_/A _11709_/Y _11708_/B vssd1 vssd1 vccd1 vccd1
+ _16206_/A sky130_fd_sc_hd__a32o_2
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12689_/A _12689_/B _12689_/C vssd1 vssd1 vccd1 vccd1 _12691_/B sky130_fd_sc_hd__o21a_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11641_ _11641_/A _11664_/A vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__xor2_4
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14360_ _14593_/A _14593_/B _14360_/C _16789_/A vssd1 vssd1 vccd1 vccd1 _14440_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11572_ _11572_/A _11576_/B _11572_/C _11572_/D vssd1 vssd1 vccd1 vccd1 _11607_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13317_/A vssd1 vssd1 vccd1 vccd1 _13431_/A sky130_fd_sc_hd__inv_2
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 i_wb_addr[24] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
X_10523_ _10437_/X _10521_/Y _10517_/A _10502_/X vssd1 vssd1 vccd1 vccd1 _10523_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14291_ _14291_/A _14372_/A vssd1 vssd1 vccd1 vccd1 _14294_/A sky130_fd_sc_hd__or2_1
X_16030_ _16315_/C _16030_/B vssd1 vssd1 vccd1 vccd1 _16136_/C sky130_fd_sc_hd__nor2_1
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13242_ _13243_/A _13243_/B vssd1 vssd1 vccd1 vccd1 _13244_/B sky130_fd_sc_hd__nand2_4
XFILLER_155_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10454_ _10454_/A _10454_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__nand2_2
XFILLER_109_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13173_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13314_/B sky130_fd_sc_hd__and2b_2
XFILLER_184_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10385_ _10385_/A _10385_/B _10385_/C vssd1 vssd1 vccd1 vccd1 _10385_/Y sky130_fd_sc_hd__nand3_2
XFILLER_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _12121_/X _12122_/Y _11915_/A _11916_/Y vssd1 vssd1 vccd1 vccd1 _12151_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16932_ _16909_/A _16851_/A _16909_/B vssd1 vssd1 vccd1 vccd1 _16932_/X sky130_fd_sc_hd__a21bo_1
X_12055_ _10657_/C _14956_/B _14911_/B vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11006_ _11006_/A _11006_/B _11097_/D vssd1 vssd1 vccd1 vccd1 _11006_/X sky130_fd_sc_hd__and3_1
XFILLER_77_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16863_ _16863_/A _16863_/B vssd1 vssd1 vccd1 vccd1 _16863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15814_ _15792_/X _15794_/X _15813_/X _16008_/C1 _15811_/A vssd1 vssd1 vccd1 vccd1
+ _15815_/A sky130_fd_sc_hd__a32o_1
X_16794_ _16794_/A _16794_/B vssd1 vssd1 vccd1 vccd1 _16795_/B sky130_fd_sc_hd__nand2_2
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15745_ _16938_/A _16020_/B vssd1 vssd1 vccd1 vccd1 _16681_/C sky130_fd_sc_hd__nand2_8
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _17405_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _12959_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11908_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11909_/B sky130_fd_sc_hd__nor2_1
XFILLER_178_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15676_ _15676_/A vssd1 vssd1 vccd1 vccd1 _15772_/A sky130_fd_sc_hd__inv_2
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12723_/A _12725_/B _12723_/B vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__o21ba_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17415_ _17415_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17415_/X sky130_fd_sc_hd__or2_1
X_14627_ _14627_/A _14627_/B _14627_/C vssd1 vssd1 vccd1 vccd1 _14628_/B sky130_fd_sc_hd__or3_1
XFILLER_53_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11839_ _10036_/D _10791_/C _11839_/S vssd1 vssd1 vccd1 vccd1 _11840_/B sky130_fd_sc_hd__mux2_1
XFILLER_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17346_ _12576_/D _17354_/A2 _17345_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17502_/D
+ sky130_fd_sc_hd__o211a_1
X_14558_ _14558_/A _14558_/B vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__nor2_1
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13509_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _17569_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17277_/X sky130_fd_sc_hd__and2_1
XFILLER_147_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14489_ _14489_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14490_/B sky130_fd_sc_hd__and2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16228_ _16315_/C _16813_/B vssd1 vssd1 vccd1 vccd1 _16229_/B sky130_fd_sc_hd__nor2_4
XFILLER_173_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16036_/A _16036_/B _16047_/X vssd1 vssd1 vccd1 vccd1 _16161_/B sky130_fd_sc_hd__a21oi_4
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08981_ _08981_/A vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__inv_2
XFILLER_142_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09602_ _09602_/A _09610_/A _09602_/C vssd1 vssd1 vccd1 vccd1 _09603_/B sky130_fd_sc_hd__or3_1
XFILLER_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09533_ _09487_/X _09530_/B _09531_/X _09532_/Y vssd1 vssd1 vccd1 vccd1 _09540_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09464_ _09748_/A _09748_/B _10308_/B _10545_/D vssd1 vssd1 vccd1 vccd1 _09473_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09395_ _09395_/A _09395_/B _09395_/C vssd1 vssd1 vccd1 vccd1 _09395_/X sky130_fd_sc_hd__or3_2
XFILLER_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ _10170_/A _10174_/A _10170_/C vssd1 vssd1 vccd1 vccd1 _10177_/B sky130_fd_sc_hd__or3_4
XFILLER_133_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout130 _17187_/Y vssd1 vssd1 vccd1 vccd1 _17270_/A2 sky130_fd_sc_hd__buf_4
Xfanout141 _15872_/A vssd1 vssd1 vccd1 vccd1 _16281_/A sky130_fd_sc_hd__buf_12
Xfanout152 _15475_/A vssd1 vssd1 vccd1 vccd1 _15726_/A sky130_fd_sc_hd__buf_6
Xfanout163 _17322_/A2 vssd1 vssd1 vccd1 vccd1 _17328_/A2 sky130_fd_sc_hd__buf_4
Xfanout174 _16168_/B vssd1 vssd1 vccd1 vccd1 _16938_/B sky130_fd_sc_hd__buf_4
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout185 _15497_/B vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__buf_12
Xfanout196 _15145_/X vssd1 vssd1 vccd1 vccd1 _15948_/A sky130_fd_sc_hd__buf_12
X_13860_ _13861_/A _13861_/B _13861_/C vssd1 vssd1 vccd1 vccd1 _13964_/A sky130_fd_sc_hd__a21o_2
XFILLER_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _12812_/B _12812_/A vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__and2b_1
X_13791_ _17409_/A _14360_/C vssd1 vssd1 vccd1 vccd1 _13792_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15530_ _15530_/A _15891_/B _15472_/A vssd1 vssd1 vccd1 vccd1 _15620_/A sky130_fd_sc_hd__or3b_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12902_/A _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _12744_/A sky130_fd_sc_hd__a21o_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12673_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__xnor2_1
X_15461_ _16012_/S _15460_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _15461_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_187_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17434_/Q _17233_/A2 _17197_/X _17199_/X _17428_/B vssd1 vssd1 vccd1 vccd1
+ _17434_/D sky130_fd_sc_hd__o221a_1
XFILLER_179_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14412_ _14413_/A _14413_/B _14413_/C vssd1 vssd1 vccd1 vccd1 _14414_/A sky130_fd_sc_hd__o21a_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15392_ _14896_/B _16008_/C1 _15391_/Y vssd1 vssd1 vccd1 vccd1 _17550_/D sky130_fd_sc_hd__a21oi_1
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_995 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17131_ _17131_/A _17131_/B _17131_/C vssd1 vssd1 vccd1 vccd1 _17131_/X sky130_fd_sc_hd__and3_1
X_14343_ _14344_/A _14344_/B _14344_/C vssd1 vssd1 vccd1 vccd1 _14413_/A sky130_fd_sc_hd__o21a_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11555_ _11555_/A _11555_/B _11637_/A vssd1 vssd1 vccd1 vccd1 _11558_/B sky130_fd_sc_hd__nor3b_2
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10506_ _10963_/A _14784_/A _10971_/B _10920_/B vssd1 vssd1 vccd1 vccd1 _10509_/A
+ sky130_fd_sc_hd__and4_1
X_14274_ _14350_/B _14274_/B vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__or2_1
X_17062_ _17062_/A _17062_/B vssd1 vssd1 vccd1 vccd1 _17063_/B sky130_fd_sc_hd__xor2_1
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _11477_/A _11477_/C _11514_/A vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__a21oi_4
XFILLER_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16013_ _16583_/A1 _13624_/X _14926_/B _16012_/X vssd1 vssd1 vccd1 vccd1 _16017_/B
+ sky130_fd_sc_hd__o22a_1
X_13225_ _13068_/A _13070_/B _13068_/B vssd1 vssd1 vccd1 vccd1 _13232_/A sky130_fd_sc_hd__o21ba_1
X_10437_ _10437_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10437_/X sky130_fd_sc_hd__and3_4
XFILLER_171_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13156_ _13852_/A _13745_/B _13903_/B _13897_/B vssd1 vssd1 vccd1 vccd1 _13157_/B
+ sky130_fd_sc_hd__and4_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10484_/B vssd1 vssd1 vccd1 vccd1 _10369_/B sky130_fd_sc_hd__inv_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12107_/A _12107_/B _12734_/D _12258_/B vssd1 vssd1 vccd1 vccd1 _12108_/B
+ sky130_fd_sc_hd__and4_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13087_/A _13220_/A vssd1 vssd1 vccd1 vccd1 _13088_/C sky130_fd_sc_hd__and2_1
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10299_ _10300_/A _10298_/Y _10299_/C _10659_/D vssd1 vssd1 vccd1 vccd1 _10418_/A
+ sky130_fd_sc_hd__and4bb_2
X_16915_ _16863_/A _16863_/B _16858_/Y vssd1 vssd1 vccd1 vccd1 _16916_/B sky130_fd_sc_hd__a21oi_1
X_12038_ _12028_/X _12037_/Y _17369_/A vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16846_ _16846_/A _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _16847_/B sky130_fd_sc_hd__or3_1
XFILLER_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16777_ _16777_/A _16777_/B _16777_/C vssd1 vssd1 vccd1 vccd1 _16778_/B sky130_fd_sc_hd__and3_1
X_13989_ _14077_/A _13989_/B vssd1 vssd1 vccd1 vccd1 _13990_/B sky130_fd_sc_hd__nor2_4
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15728_ _15834_/A _15728_/B vssd1 vssd1 vccd1 vccd1 _15730_/B sky130_fd_sc_hd__nor2_4
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15659_ _15660_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _15661_/B sky130_fd_sc_hd__nand2_2
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09180_ _09358_/A _09345_/B vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__and2_2
XFILLER_159_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ input43/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17329_/X sky130_fd_sc_hd__or3_1
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08964_ _12546_/B _12752_/B vssd1 vssd1 vccd1 vccd1 _08993_/C sky130_fd_sc_hd__nand2_4
XFILLER_88_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__xnor2_4
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09516_ _09517_/A _09515_/Y _10321_/A _09803_/B vssd1 vssd1 vccd1 vccd1 _09636_/A
+ sky130_fd_sc_hd__and4bb_1
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09447_ _09447_/A _09583_/A vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__nor2_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09378_ _09379_/A _09377_/Y _10062_/A _09937_/B vssd1 vssd1 vccd1 vccd1 _09513_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_910 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ _11340_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11341_/C sky130_fd_sc_hd__xnor2_2
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11271_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11274_/C sky130_fd_sc_hd__nand2_2
XFILLER_180_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13010_ _13268_/A _13010_/B vssd1 vssd1 vccd1 vccd1 _13138_/B sky130_fd_sc_hd__nand2b_1
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10222_ _10560_/B _09937_/B _09953_/B _09952_/A vssd1 vssd1 vccd1 vccd1 _10226_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _10149_/A _10152_/X _10137_/X _10138_/Y vssd1 vssd1 vccd1 vccd1 _10155_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14961_ _15460_/B _15458_/B _15458_/A vssd1 vssd1 vccd1 vccd1 _14961_/X sky130_fd_sc_hd__mux2_4
XFILLER_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16700_ _16701_/A _16701_/B vssd1 vssd1 vccd1 vccd1 _16777_/B sky130_fd_sc_hd__or2_2
X_13912_ _13912_/A _13912_/B vssd1 vssd1 vccd1 vccd1 _13913_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14892_ _15204_/A _16683_/A _16807_/A vssd1 vssd1 vccd1 vccd1 _15208_/C sky130_fd_sc_hd__or3_4
XFILLER_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16631_ _16711_/A _16631_/B vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__or2_2
X_13843_ _13844_/B _14181_/B _13844_/D _13844_/A vssd1 vssd1 vccd1 vccd1 _13845_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16562_ _16561_/X _16562_/B _16562_/C vssd1 vssd1 vccd1 vccd1 _16562_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13774_ _13774_/A _13774_/B vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__nand2_2
XFILLER_15_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15513_ _15514_/A _15514_/B _15514_/C vssd1 vssd1 vccd1 vccd1 _15609_/A sky130_fd_sc_hd__a21oi_2
X_12725_ _12725_/A _12725_/B vssd1 vssd1 vccd1 vccd1 _12727_/B sky130_fd_sc_hd__xnor2_1
XFILLER_188_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16493_ _16483_/X _16493_/B _16493_/C vssd1 vssd1 vccd1 vccd1 _16493_/X sky130_fd_sc_hd__and3b_1
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15444_ _15442_/Y _15443_/X _16911_/A vssd1 vssd1 vccd1 vccd1 _15444_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_188_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ _12657_/B _13194_/D _13067_/D _12657_/A vssd1 vssd1 vccd1 vccd1 _12658_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_90_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _11607_/A _11607_/B _11607_/C vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__nand3_2
X_12587_ _12588_/A _12588_/B _12588_/C vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__a21oi_4
X_15375_ _15307_/B _15307_/C _15307_/A vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__o21ba_2
XFILLER_156_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17114_ _14828_/Y _17169_/A1 _17104_/X _17107_/X _17113_/X vssd1 vssd1 vccd1 vccd1
+ _17114_/X sky130_fd_sc_hd__o311a_1
XFILLER_190_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14326_ _14326_/A _14554_/B _14326_/C vssd1 vssd1 vccd1 vccd1 _14393_/B sky130_fd_sc_hd__nand3_2
X_11538_ _11538_/A _11538_/B vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__or2_1
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap116 _13941_/B vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__buf_2
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17045_ _17046_/A _17046_/B _17046_/C vssd1 vssd1 vccd1 vccd1 _17088_/A sky130_fd_sc_hd__o21a_1
X_14257_ _14258_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14257_/Y sky130_fd_sc_hd__nand2_1
Xmax_cap138 _16315_/B vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__buf_6
X_11469_ _14791_/A _11629_/C vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__and2_2
XFILLER_109_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13208_ _14769_/A _14770_/A _13966_/D _13866_/D vssd1 vssd1 vccd1 vccd1 _13339_/A
+ sky130_fd_sc_hd__and4_2
X_14188_ _14188_/A _14188_/B _14188_/C vssd1 vssd1 vccd1 vccd1 _14189_/B sky130_fd_sc_hd__and3_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13139_ _13268_/B _13140_/B vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__or2_1
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16829_ _16829_/A _16829_/B vssd1 vssd1 vccd1 vccd1 _16830_/B sky130_fd_sc_hd__xnor2_2
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09301_ _09302_/A _09300_/Y _11902_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _09443_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_179_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09232_ _12174_/B _12129_/B _12127_/C _12174_/A vssd1 vssd1 vccd1 vccd1 _09234_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ _09164_/A _09163_/B _12546_/B _09350_/B vssd1 vssd1 vccd1 vccd1 _09354_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09094_ _08973_/B _08971_/C _08993_/C vssd1 vssd1 vccd1 vccd1 _09095_/B sky130_fd_sc_hd__o21a_1
XFILLER_108_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__xnor2_4
XFILLER_131_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08947_ _11895_/A _12592_/B _12090_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _08950_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ _08883_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _08889_/A sky130_fd_sc_hd__nor2_2
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _10933_/B _10933_/D _10970_/B _10933_/A vssd1 vssd1 vccd1 vccd1 _10841_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_53_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ _10771_/A _10771_/B _10771_/C vssd1 vssd1 vccd1 vccd1 _10772_/B sky130_fd_sc_hd__or3_1
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _12339_/A _12341_/B _12339_/B vssd1 vssd1 vccd1 vccd1 _12511_/B sky130_fd_sc_hd__o21ba_4
X_13490_ _13607_/A _13490_/B _13490_/C _13490_/D vssd1 vssd1 vccd1 vccd1 _13607_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _12442_/A _12442_/B _12442_/C vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__a21oi_2
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12372_ _12373_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__or2_4
X_15160_ _15161_/A _15161_/B vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__or2_2
XFILLER_138_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14111_ _14197_/B _14111_/B vssd1 vssd1 vccd1 vccd1 _14113_/C sky130_fd_sc_hd__nand2_1
X_11323_ _11377_/B _11561_/C _11563_/D _11322_/A vssd1 vssd1 vccd1 vccd1 _11324_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15091_ _15091_/A _15091_/B vssd1 vssd1 vccd1 vccd1 _15170_/B sky130_fd_sc_hd__or2_2
XFILLER_125_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14042_ _14043_/A _14043_/B vssd1 vssd1 vccd1 vccd1 _14042_/Y sky130_fd_sc_hd__nand2_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11254_ _11139_/A _11139_/B _11139_/C vssd1 vssd1 vccd1 vccd1 _11255_/C sky130_fd_sc_hd__a21oi_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10469_/B _10205_/B vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__nor2_2
XFILLER_69_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11185_ _11182_/Y _11183_/X _11039_/Y _11041_/Y vssd1 vssd1 vccd1 vccd1 _11186_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10138_/C sky130_fd_sc_hd__xnor2_2
XFILLER_121_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15993_ _15991_/X _15994_/B vssd1 vssd1 vccd1 vccd1 _15993_/X sky130_fd_sc_hd__and2b_2
X_10067_ _10067_/A _10067_/B _10067_/C vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__and3_2
XFILLER_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14944_ _14944_/A _14944_/B _14944_/C vssd1 vssd1 vccd1 vccd1 _14944_/Y sky130_fd_sc_hd__nor3_1
XFILLER_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14875_ _14888_/C _14876_/C _14876_/D vssd1 vssd1 vccd1 vccd1 _14875_/X sky130_fd_sc_hd__or3_1
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16614_ _16614_/A _16614_/B vssd1 vssd1 vccd1 vccd1 _16616_/C sky130_fd_sc_hd__xnor2_2
XFILLER_78_1059 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13826_ _13824_/A _13824_/B _13827_/A vssd1 vssd1 vccd1 vccd1 _13826_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17594_ fanout941/X _17594_/D vssd1 vssd1 vccd1 vccd1 _17594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16545_ _16545_/A _16545_/B vssd1 vssd1 vccd1 vccd1 _16547_/B sky130_fd_sc_hd__xnor2_1
X_13757_ _13756_/B _13757_/B vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__and2b_1
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _10969_/A _10969_/B vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__xnor2_4
XFILLER_149_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12708_ _12040_/Y _12042_/Y _12397_/B _12061_/Y _12383_/S _16011_/B vssd1 vssd1 vccd1
+ vccd1 _12709_/B sky130_fd_sc_hd__mux4_2
XFILLER_188_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16476_ _11200_/Y _16389_/C _11229_/Y vssd1 vssd1 vccd1 vccd1 _16478_/A sky130_fd_sc_hd__a21oi_1
XFILLER_148_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13688_ _13688_/A _13688_/B vssd1 vssd1 vccd1 vccd1 _13707_/A sky130_fd_sc_hd__xor2_2
XFILLER_129_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15427_ _15340_/X _15345_/B _15342_/Y vssd1 vssd1 vccd1 vccd1 _15429_/B sky130_fd_sc_hd__o21ai_4
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12639_ _12640_/A _12792_/A _12640_/C vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__o21a_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1051 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15358_ _15358_/A _15358_/B vssd1 vssd1 vccd1 vccd1 _15359_/B sky130_fd_sc_hd__xnor2_4
XFILLER_102_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ _14309_/A _14309_/B vssd1 vssd1 vccd1 vccd1 _14312_/A sky130_fd_sc_hd__xor2_1
X_15289_ _15774_/A _16136_/B vssd1 vssd1 vccd1 vccd1 _15291_/B sky130_fd_sc_hd__nand2_2
XFILLER_176_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17028_ _17028_/A _17028_/B vssd1 vssd1 vccd1 vccd1 _17029_/C sky130_fd_sc_hd__nor2_1
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09850_ _09863_/B _09863_/C _09863_/A vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__a21o_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout707 _15101_/A1 vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__buf_4
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout718 _16480_/A vssd1 vssd1 vccd1 vccd1 _14050_/D sky130_fd_sc_hd__clkbuf_16
XFILLER_124_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 _12068_/C vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__clkbuf_16
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08801_/Y sky130_fd_sc_hd__nand3_4
XFILLER_113_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09926_/A _09928_/D _14949_/A vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_86_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _17609_/Q _17610_/Q vssd1 vssd1 vccd1 vccd1 _08732_/X sky130_fd_sc_hd__and2_1
XFILLER_66_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_27_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _11953_/B _12338_/C _12338_/D _11953_/A vssd1 vssd1 vccd1 vccd1 _09219_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ _09147_/B _09231_/B vssd1 vssd1 vccd1 vccd1 _09148_/B sky130_fd_sc_hd__nor2_2
XFILLER_33_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _09091_/A sky130_fd_sc_hd__xnor2_1
XFILLER_163_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09979_ _10236_/A _10236_/B _10479_/B _17468_/D vssd1 vssd1 vccd1 vccd1 _09982_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_76_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _12987_/X _12988_/Y _12819_/X _12824_/A vssd1 vssd1 vccd1 vccd1 _12993_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11941_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11941_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14661_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _14662_/B sky130_fd_sc_hd__nor2_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__inv_2
XFILLER_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _13718_/B _13609_/X _13495_/A _13497_/X vssd1 vssd1 vccd1 vccd1 _13612_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _10823_/A _10823_/B _10829_/B vssd1 vssd1 vccd1 vccd1 _11072_/B sky130_fd_sc_hd__or3_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14591_ _17164_/A _12037_/A _13625_/Y _12853_/X vssd1 vssd1 vccd1 vccd1 _14591_/X
+ sky130_fd_sc_hd__a31o_2
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16330_ _16239_/A _16239_/B _16231_/Y vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__a21bo_1
XFILLER_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13542_ _13542_/A vssd1 vssd1 vccd1 vccd1 _13543_/B sky130_fd_sc_hd__clkinv_2
XFILLER_164_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _15126_/A _10993_/D _10543_/C vssd1 vssd1 vccd1 vccd1 _10754_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _16358_/A _16261_/B vssd1 vssd1 vccd1 vccd1 _16262_/C sky130_fd_sc_hd__or2_1
X_13473_ _13473_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__xnor2_1
X_10685_ _10685_/A _10685_/B _10685_/C vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__nand3_4
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15212_ _15948_/A _15932_/B vssd1 vssd1 vccd1 vccd1 _15213_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ _17391_/A _17389_/A _12576_/D _12567_/B vssd1 vssd1 vccd1 vccd1 _12425_/B
+ sky130_fd_sc_hd__and4_1
X_16192_ _16192_/A _16192_/B vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__xnor2_2
XFILLER_166_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15143_ _15143_/A _15270_/B _15143_/C vssd1 vssd1 vccd1 vccd1 _15143_/X sky130_fd_sc_hd__or3_4
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12357_/B sky130_fd_sc_hd__xnor2_4
XFILLER_181_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ _11306_/A _11306_/B vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__nor2_2
X_15074_ _15475_/A _16226_/C vssd1 vssd1 vccd1 vccd1 _15913_/A sky130_fd_sc_hd__nand2_8
X_12286_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12286_/Y sky130_fd_sc_hd__nand3_2
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14025_ _14025_/A _14025_/B vssd1 vssd1 vccd1 vccd1 _14025_/Y sky130_fd_sc_hd__xnor2_1
X_11237_ _11237_/A _11237_/B vssd1 vssd1 vccd1 vccd1 _11295_/A sky130_fd_sc_hd__nand2_4
XFILLER_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11168_ _11168_/A _11168_/B _11167_/X vssd1 vssd1 vccd1 vccd1 _11168_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_121_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10119_ _10119_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__xnor2_4
XFILLER_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15976_ _15976_/A _15976_/B vssd1 vssd1 vccd1 vccd1 _15984_/A sky130_fd_sc_hd__xnor2_4
X_11099_ _11099_/A _11099_/B _11101_/B vssd1 vssd1 vccd1 vccd1 _11104_/B sky130_fd_sc_hd__or3_2
X_14927_ _16011_/A _14919_/X _14923_/Y _17164_/C vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_82_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14858_ _16114_/A _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16115_/B sky130_fd_sc_hd__and3_2
XFILLER_64_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13809_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _13810_/B sky130_fd_sc_hd__and2_1
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17577_ fanout936/X _17577_/D vssd1 vssd1 vccd1 vccd1 _17577_/Q sky130_fd_sc_hd__dfxtp_1
X_14789_ _14789_/A _14848_/A vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16528_ _16630_/A _16528_/B vssd1 vssd1 vccd1 vccd1 _16547_/A sky130_fd_sc_hd__and2_1
XFILLER_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16459_ _16459_/A _16459_/B vssd1 vssd1 vccd1 vccd1 _16460_/B sky130_fd_sc_hd__or2_1
XFILLER_192_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09000_ _11932_/A _12752_/B vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__nand2_2
XFILLER_164_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_144_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _09902_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _10034_/C sky130_fd_sc_hd__xnor2_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout504 _15396_/A vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__buf_6
Xfanout515 _12104_/A vssd1 vssd1 vccd1 vccd1 _17375_/A sky130_fd_sc_hd__buf_6
XFILLER_141_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout526 _09470_/A vssd1 vssd1 vccd1 vccd1 _12135_/A sky130_fd_sc_hd__buf_6
X_09833_ _09720_/A _09719_/C _09719_/B vssd1 vssd1 vccd1 vccd1 _09866_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout537 _11322_/A vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__buf_6
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout548 _10532_/B vssd1 vssd1 vccd1 vccd1 _14790_/A sky130_fd_sc_hd__buf_2
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout559 _13390_/S vssd1 vssd1 vccd1 vccd1 _13837_/A sky130_fd_sc_hd__buf_2
XFILLER_100_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09788_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09765_/C sky130_fd_sc_hd__and2_1
XFILLER_101_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09695_ _09695_/A _09842_/A vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__nor2_4
XFILLER_27_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1024 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10470_ _10470_/A _10470_/B vssd1 vssd1 vccd1 vccd1 _10582_/A sky130_fd_sc_hd__or2_1
XFILLER_109_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09129_ _09502_/A _09803_/B _09126_/Y _09139_/A vssd1 vssd1 vccd1 vccd1 _09130_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _12141_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__nand2_2
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12071_ _12237_/A _12645_/B _12070_/C _12070_/D vssd1 vssd1 vccd1 vccd1 _12072_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11022_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11024_/C sky130_fd_sc_hd__xor2_4
XFILLER_173_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15830_ _16315_/C _15932_/A _16039_/B _16150_/B vssd1 vssd1 vccd1 vccd1 _15831_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _15762_/A _15762_/B vssd1 vssd1 vccd1 vccd1 _15868_/A sky130_fd_sc_hd__and2_1
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12973_ _12974_/A _12974_/B vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__or2_2
XTAP_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17500_ fanout932/X _17500_/D vssd1 vssd1 vccd1 vccd1 _17500_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14744_/A _14712_/B vssd1 vssd1 vccd1 vccd1 _14713_/C sky130_fd_sc_hd__xnor2_2
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__and2_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15591_/A _15600_/Y _15779_/B _15691_/Y vssd1 vssd1 vccd1 vccd1 _15786_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_79_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ input47/X _17608_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17608_/D sky130_fd_sc_hd__mux2_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14676_/A _14708_/D _14644_/C vssd1 vssd1 vccd1 vccd1 _14645_/A sky130_fd_sc_hd__a21oi_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11855_ _14356_/S _11854_/X _15457_/A vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__o21a_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _10963_/B _10805_/C _10957_/D _11095_/A vssd1 vssd1 vccd1 vccd1 _10807_/B
+ sky130_fd_sc_hd__a22oi_4
X_17362_ _17362_/A _17362_/B _17362_/C _17362_/D vssd1 vssd1 vccd1 vccd1 _17362_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14574_ _14574_/A vssd1 vssd1 vccd1 vccd1 _14575_/B sky130_fd_sc_hd__inv_2
X_11786_ _12016_/A _09826_/A _14837_/A _16922_/A vssd1 vssd1 vccd1 vccd1 _11786_/Y
+ sky130_fd_sc_hd__o31ai_1
X_16313_ _16313_/A vssd1 vssd1 vccd1 vccd1 _17560_/D sky130_fd_sc_hd__inv_2
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _13524_/C _13637_/A _13523_/Y vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__a21bo_1
X_17293_ _17465_/Q _17293_/A2 _17291_/X _17292_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17465_/D sky130_fd_sc_hd__o221a_1
X_10737_ _11258_/B _10839_/D _10971_/B _11314_/A vssd1 vssd1 vccd1 vccd1 _10737_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_174_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16244_ _16814_/A _16827_/A vssd1 vssd1 vccd1 vccd1 _16245_/B sky130_fd_sc_hd__nor2_1
X_13456_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13576_/A sky130_fd_sc_hd__o21ai_1
XFILLER_185_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ wire120/X _10667_/Y _10556_/B _10587_/Y vssd1 vssd1 vccd1 vccd1 _10678_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _17401_/A _13966_/D _12408_/C vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__a21oi_2
X_16175_ _16175_/A _16175_/B vssd1 vssd1 vccd1 vccd1 _16177_/B sky130_fd_sc_hd__xor2_2
XFILLER_127_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10599_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__xor2_4
X_13387_ _13508_/B _13388_/B vssd1 vssd1 vccd1 vccd1 _13387_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput107 _17464_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15126_ _15126_/A _15126_/B vssd1 vssd1 vccd1 vccd1 _15126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_182_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12338_ _12657_/A _12657_/B _12338_/C _12338_/D vssd1 vssd1 vccd1 vccd1 _12339_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_86_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _15056_/A _14913_/Y _15056_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _15057_/X
+ sky130_fd_sc_hd__a211o_2
X_12269_ _12270_/B _12270_/C _12270_/D _17379_/A vssd1 vssd1 vccd1 vccd1 _12271_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_141_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14008_ _14008_/A _14089_/B _14008_/C vssd1 vssd1 vccd1 vccd1 _14115_/B sky130_fd_sc_hd__nand3_2
XFILLER_96_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_110_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15959_ _16171_/A _16589_/B vssd1 vssd1 vccd1 vccd1 _15960_/B sky130_fd_sc_hd__nand2_4
XFILLER_37_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09480_ _09480_/A _09480_/B _09480_/C vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__and3_4
XFILLER_64_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout301 _14666_/S vssd1 vssd1 vccd1 vccd1 _14840_/A sky130_fd_sc_hd__buf_6
XFILLER_120_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout312 _17609_/Q vssd1 vssd1 vccd1 vccd1 _17476_/D sky130_fd_sc_hd__buf_8
Xfanout323 _17540_/Q vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout334 _17539_/Q vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout345 _17537_/Q vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__buf_8
Xfanout356 _17536_/Q vssd1 vssd1 vccd1 vccd1 _12659_/A sky130_fd_sc_hd__clkbuf_16
X_09816_ _09668_/Y _09683_/X _09772_/X _09813_/X vssd1 vssd1 vccd1 vccd1 _09817_/B
+ sky130_fd_sc_hd__a211o_1
Xfanout367 _17534_/Q vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__buf_12
XFILLER_87_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout378 _17409_/A vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__buf_6
XFILLER_189_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout389 _12500_/A vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_28_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09747_ _09747_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__nand2_2
XFILLER_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09678_/A _09678_/B _09681_/A vssd1 vssd1 vccd1 vccd1 _09679_/B sky130_fd_sc_hd__nor3_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11663_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__nor2_4
XFILLER_168_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11571_ _15305_/C _11423_/C _11605_/B _11423_/A vssd1 vssd1 vccd1 vccd1 _11572_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13312_/A _13312_/B _13312_/C vssd1 vssd1 vccd1 vccd1 _13317_/A sky130_fd_sc_hd__o21ai_4
X_10522_ _10502_/X _10517_/A _10521_/Y _10437_/X vssd1 vssd1 vccd1 vccd1 _10566_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14290_ _14290_/A _14708_/B _16789_/A _16722_/A vssd1 vssd1 vccd1 vccd1 _14372_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10453_ _10453_/A _10453_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10454_/B sky130_fd_sc_hd__nand3_1
X_13241_ _13241_/A _13241_/B vssd1 vssd1 vccd1 vccd1 _13243_/B sky130_fd_sc_hd__xnor2_2
XFILLER_108_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13172_ _13172_/A _13172_/B vssd1 vssd1 vccd1 vccd1 _13174_/B sky130_fd_sc_hd__xnor2_4
X_10384_ _10385_/A _10385_/B _10385_/C vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__and3_1
XFILLER_184_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12123_ _11915_/A _11916_/Y _12121_/X _12122_/Y vssd1 vssd1 vccd1 vccd1 _12316_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_112_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16931_ _16931_/A _16931_/B _16910_/B vssd1 vssd1 vccd1 vccd1 _16931_/X sky130_fd_sc_hd__or3b_2
X_12054_ _12054_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _14956_/B sky130_fd_sc_hd__and2_1
XFILLER_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11005_ _11005_/A _11005_/B vssd1 vssd1 vccd1 vccd1 _11009_/A sky130_fd_sc_hd__nand2_2
XFILLER_120_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16862_ _16863_/A _16863_/B vssd1 vssd1 vccd1 vccd1 _16862_/X sky130_fd_sc_hd__or2_1
XFILLER_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout890 _17479_/Q vssd1 vssd1 vccd1 vccd1 _11027_/C sky130_fd_sc_hd__buf_4
X_15813_ _16304_/A _15802_/Y _15812_/X _15800_/Y vssd1 vssd1 vccd1 vccd1 _15813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16793_ _17156_/B _16793_/B vssd1 vssd1 vccd1 vccd1 _16793_/X sky130_fd_sc_hd__or2_1
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15744_ _16938_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16165_/B sky130_fd_sc_hd__and2_4
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12956_ _12956_/A _12956_/B vssd1 vssd1 vccd1 vccd1 _12959_/A sky130_fd_sc_hd__nand2_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11907_ _11908_/A _11908_/B vssd1 vssd1 vccd1 vccd1 _11909_/A sky130_fd_sc_hd__and2_2
X_15675_ _15675_/A _15675_/B vssd1 vssd1 vccd1 vccd1 _15676_/A sky130_fd_sc_hd__nor2_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12887_ _12735_/A _12737_/B _12735_/B vssd1 vssd1 vccd1 vccd1 _12897_/A sky130_fd_sc_hd__o21ba_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ input53/X _17426_/A2 _17413_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17535_/D
+ sky130_fd_sc_hd__o211a_1
X_14626_ _14627_/A _14627_/B _14627_/C vssd1 vssd1 vccd1 vccd1 _14638_/A sky130_fd_sc_hd__o21ai_2
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _11835_/Y _11837_/Y _15096_/S vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ input52/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17345_/X sky130_fd_sc_hd__or3_1
X_14557_ _14557_/A _14557_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14558_/B sky130_fd_sc_hd__nor3_1
X_11769_ _11768_/A _16866_/A _16866_/B _11767_/X vssd1 vssd1 vccd1 vccd1 _16972_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13508_ _13271_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__and2b_1
XFILLER_159_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17276_ _17601_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17276_/X sky130_fd_sc_hd__a21o_1
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _14489_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14557_/B sky130_fd_sc_hd__nor2_1
XFILLER_147_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16227_ _16227_/A _16227_/B vssd1 vssd1 vccd1 vccd1 _16229_/A sky130_fd_sc_hd__nor2_4
X_13439_ _13586_/B _13439_/B vssd1 vssd1 vccd1 vccd1 _13442_/B sky130_fd_sc_hd__nor2_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _16158_/A _16158_/B vssd1 vssd1 vccd1 vccd1 _16161_/A sky130_fd_sc_hd__xnor2_4
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15109_ _11472_/B _14791_/X _14797_/X _15108_/Y vssd1 vssd1 vccd1 vccd1 _15109_/X
+ sky130_fd_sc_hd__a31o_1
X_16089_ _16089_/A _16089_/B vssd1 vssd1 vccd1 vccd1 _16092_/A sky130_fd_sc_hd__xnor2_4
X_08980_ _09238_/B _08980_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__or2_1
XFILLER_102_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09601_ _09480_/X _09599_/Y _09597_/B _09580_/X vssd1 vssd1 vccd1 vccd1 _09601_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09532_ _09393_/X _09398_/Y _09485_/X _09530_/X vssd1 vssd1 vccd1 vccd1 _09532_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_37_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09463_/A _09463_/B vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09394_ _09395_/B _09395_/C _09395_/A vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__o21ai_4
XFILLER_177_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout131 _16760_/B vssd1 vssd1 vccd1 vccd1 _16246_/A sky130_fd_sc_hd__buf_8
Xfanout142 _15821_/A vssd1 vssd1 vccd1 vccd1 _16226_/B sky130_fd_sc_hd__buf_4
Xfanout153 _16056_/A vssd1 vssd1 vccd1 vccd1 _15660_/A sky130_fd_sc_hd__buf_6
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout164 _17296_/Y vssd1 vssd1 vccd1 vccd1 _17322_/A2 sky130_fd_sc_hd__buf_4
Xfanout175 _15575_/Y vssd1 vssd1 vccd1 vccd1 _16814_/B sky130_fd_sc_hd__buf_6
Xfanout186 _15752_/B vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__buf_4
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout197 _15145_/X vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12810_ _12658_/A _12660_/B _12658_/B vssd1 vssd1 vccd1 vccd1 _12812_/B sky130_fd_sc_hd__o21ba_4
X_13790_ _13790_/A _13790_/B vssd1 vssd1 vccd1 vccd1 _13792_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12743_/C sky130_fd_sc_hd__xnor2_2
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _16011_/A _15460_/B vssd1 vssd1 vccd1 vccd1 _15460_/X sky130_fd_sc_hd__or2_2
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12672_ _12673_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _12672_/X sky130_fd_sc_hd__or2_2
XFILLER_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14411_ _14473_/B _14411_/B vssd1 vssd1 vccd1 vccd1 _14413_/C sky130_fd_sc_hd__and2_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11583_/B _11587_/X _11617_/B _11616_/Y vssd1 vssd1 vccd1 vccd1 _11624_/B
+ sky130_fd_sc_hd__a211o_1
X_15391_ _16911_/A _15369_/Y _15390_/Y vssd1 vssd1 vccd1 vccd1 _15391_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_179_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17130_ _17130_/A _17130_/B vssd1 vssd1 vccd1 vccd1 _17131_/C sky130_fd_sc_hd__or2_1
X_14342_ _14342_/A _14342_/B vssd1 vssd1 vccd1 vccd1 _14344_/C sky130_fd_sc_hd__and2_1
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11554_ _15116_/A _15274_/A _11506_/X _11507_/Y vssd1 vssd1 vccd1 vccd1 _11555_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17061_ _17060_/A _17060_/B _17062_/A vssd1 vssd1 vccd1 vccd1 _17096_/B sky130_fd_sc_hd__o21a_1
XFILLER_7_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10505_ _10505_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__nor2_2
X_14273_ _14273_/A _14273_/B _14273_/C vssd1 vssd1 vccd1 vccd1 _14274_/B sky130_fd_sc_hd__and3_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11485_ _11534_/A _11485_/B vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__and2_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _16010_/X _16011_/X _16012_/S vssd1 vssd1 vccd1 vccd1 _16012_/X sky130_fd_sc_hd__mux2_1
X_13224_ _13224_/A _13224_/B vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__and2_2
XFILLER_183_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10436_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _10437_/C sky130_fd_sc_hd__xnor2_4
X_13155_ _13745_/B _13903_/B _13897_/B _13852_/A vssd1 vssd1 vccd1 vccd1 _13157_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_124_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10367_ _10370_/C _10367_/B vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__xnor2_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12107_/B _12734_/D _12258_/B _12107_/A vssd1 vssd1 vccd1 vccd1 _12108_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10171_/B _10755_/D _10534_/D _10419_/A vssd1 vssd1 vccd1 vccd1 _10298_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13086_ _13085_/A _13085_/B _13085_/C vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__o21ai_2
XFILLER_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16914_ _16914_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16916_/A sky130_fd_sc_hd__nor2_2
X_12037_ _12037_/A vssd1 vssd1 vccd1 vccd1 _12037_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16845_ _16846_/A _16846_/B _16846_/C vssd1 vssd1 vccd1 vccd1 _16909_/A sky130_fd_sc_hd__o21ai_2
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16776_ _16777_/A _16777_/B _16777_/C vssd1 vssd1 vccd1 vccd1 _16846_/A sky130_fd_sc_hd__a21oi_2
X_13988_ _13988_/A _13988_/B vssd1 vssd1 vccd1 vccd1 _13989_/B sky130_fd_sc_hd__and2_1
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _16025_/A _16499_/B _15820_/C _15820_/A vssd1 vssd1 vccd1 vccd1 _15728_/B
+ sky130_fd_sc_hd__o22a_2
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12939_ _12817_/A _12817_/B _12815_/Y vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__a21bo_2
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15658_ _15703_/A _15658_/B vssd1 vssd1 vccd1 vccd1 _15658_/Y sky130_fd_sc_hd__nand2_4
XFILLER_33_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14609_ _14609_/A _14609_/B vssd1 vssd1 vccd1 vccd1 _14610_/B sky130_fd_sc_hd__and2_1
X_15589_ _15590_/A _15590_/B _15590_/C vssd1 vssd1 vccd1 vccd1 _15591_/A sky130_fd_sc_hd__a21oi_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17328_ _13664_/D _17328_/A2 _17327_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17493_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_18_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17259_ _17563_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17259_/X sky130_fd_sc_hd__and2_1
XFILLER_179_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08963_ _12546_/B _12592_/C _12752_/B _12845_/S vssd1 vssd1 vccd1 vccd1 _08963_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__nand2b_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09515_ _09637_/B _09947_/B _10067_/B _11953_/A vssd1 vssd1 vccd1 vccd1 _09515_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09447_/A _09445_/Y _11902_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _09583_/A
+ sky130_fd_sc_hd__and4bb_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09377_ _09637_/B _09803_/B _09947_/B _09942_/A vssd1 vssd1 vccd1 vccd1 _09377_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_149_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _11270_/A _11270_/B vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__xnor2_4
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10221_ _10223_/B _10223_/A vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__and2b_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__and2_2
XFILLER_160_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10083_ _10209_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__or2_1
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14960_ _14955_/X _14959_/X _15035_/S vssd1 vssd1 vccd1 vccd1 _15458_/B sky130_fd_sc_hd__mux2_1
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _13912_/A _13912_/B vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__or2_2
X_14891_ _14881_/X _14889_/X _08723_/Y vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__a21o_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16630_ _16630_/A _16630_/B _16630_/C vssd1 vssd1 vccd1 vccd1 _16631_/B sky130_fd_sc_hd__and3_1
XFILLER_75_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13842_ _14734_/A _13839_/X _13841_/X _14758_/A vssd1 vssd1 vccd1 vccd1 _13842_/X
+ sky130_fd_sc_hd__a22o_2
Xwb_buttons_leds_950 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_950/HI led_enb[3] sky130_fd_sc_hd__conb_1
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16561_ _16563_/B _16564_/A _16385_/A vssd1 vssd1 vccd1 vccd1 _16561_/X sky130_fd_sc_hd__or3b_2
XFILLER_16_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13773_ _14153_/A _14153_/B _14141_/D _14050_/D vssd1 vssd1 vccd1 vccd1 _13774_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10985_ _10985_/A _10985_/B vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__xnor2_4
XFILLER_188_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15512_ _15512_/A _15512_/B vssd1 vssd1 vccd1 vccd1 _15514_/C sky130_fd_sc_hd__xor2_2
X_12724_ _17393_/A _14153_/C vssd1 vssd1 vccd1 vccd1 _12725_/B sky130_fd_sc_hd__nand2_1
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16492_ _16492_/A _16492_/B _16492_/C vssd1 vssd1 vccd1 vccd1 _16493_/C sky130_fd_sc_hd__and3_1
XFILLER_188_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15443_ _15367_/B _15369_/B _15365_/X vssd1 vssd1 vccd1 vccd1 _15443_/X sky130_fd_sc_hd__a21o_1
X_12655_ _12655_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__and2_1
XFILLER_169_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11606_ _11576_/B _11572_/C _11572_/D _11572_/A vssd1 vssd1 vccd1 vccd1 _11607_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _15374_/X sky130_fd_sc_hd__or2_1
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12586_ _12586_/A _12586_/B vssd1 vssd1 vccd1 vccd1 _12588_/C sky130_fd_sc_hd__or2_2
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17113_ _17113_/A _17113_/B _17113_/C vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__and3_1
X_14325_ _14325_/A _14325_/B vssd1 vssd1 vccd1 vccd1 _14326_/C sky130_fd_sc_hd__xnor2_2
XFILLER_157_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11537_ _11538_/A _11537_/B _11537_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__nor3_4
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17044_ _17044_/A _17085_/B vssd1 vssd1 vccd1 vccd1 _17046_/C sky130_fd_sc_hd__nor2_1
Xmax_cap117 _09393_/B vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__buf_2
X_14256_ _14258_/A _14258_/B vssd1 vssd1 vccd1 vccd1 _14256_/X sky130_fd_sc_hd__and2_2
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ _11506_/A _11553_/A _15401_/A _11506_/C vssd1 vssd1 vccd1 vccd1 _11468_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1050 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13207_ _14770_/A _13966_/D _13866_/D _14769_/A vssd1 vssd1 vccd1 vccd1 _13211_/A
+ sky130_fd_sc_hd__a22oi_4
X_10419_ _10419_/A _10532_/B _10534_/D _10647_/D vssd1 vssd1 vccd1 vccd1 _10422_/A
+ sky130_fd_sc_hd__and4_1
X_14187_ _14188_/A _14188_/B _14188_/C vssd1 vssd1 vccd1 vccd1 _14268_/A sky130_fd_sc_hd__a21oi_4
XFILLER_171_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11400_/C sky130_fd_sc_hd__xnor2_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13002_/A _13138_/B vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__and2b_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _17421_/A _13321_/D vssd1 vssd1 vccd1 vccd1 _13070_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16828_ _16828_/A _16828_/B vssd1 vssd1 vccd1 vccd1 _16829_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16759_ _16759_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16761_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09300_ _12595_/B _11867_/C _12795_/B _09584_/A vssd1 vssd1 vccd1 vccd1 _09300_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_34_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ _09231_/A _09231_/B vssd1 vssd1 vccd1 vccd1 _09240_/A sky130_fd_sc_hd__or2_1
XFILLER_181_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09162_ _12845_/S _11813_/B _08969_/C vssd1 vssd1 vccd1 vccd1 _09163_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ _09093_/A _09093_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__nand2_2
XFILLER_175_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09995_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _09025_/C _12158_/C _08808_/A _08806_/Y vssd1 vssd1 vccd1 vccd1 _08883_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_57_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _10771_/A _10771_/B _10771_/C vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__o21ai_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09429_ _16990_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__nand2_2
XFILLER_185_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ _12440_/A _12616_/A vssd1 vssd1 vccd1 vccd1 _12442_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _12371_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12373_/B sky130_fd_sc_hd__nor2_4
XFILLER_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ _14015_/B _14110_/B vssd1 vssd1 vccd1 vccd1 _14111_/B sky130_fd_sc_hd__nand2b_1
XFILLER_176_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11322_ _11322_/A _11377_/B _11561_/C _11563_/D vssd1 vssd1 vccd1 vccd1 _11325_/A
+ sky130_fd_sc_hd__nand4_4
X_15090_ _15091_/A _15091_/B vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14041_ _13947_/Y _13951_/B _14040_/X vssd1 vssd1 vccd1 vccd1 _14043_/B sky130_fd_sc_hd__o21a_2
XFILLER_153_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11253_ _11348_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__xor2_4
XFILLER_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _10559_/A _10805_/C _10203_/C vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__a21oi_1
X_11184_ _11039_/Y _11041_/Y _11182_/Y _11183_/X vssd1 vssd1 vccd1 vccd1 _11218_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_192_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10135_ _10134_/A _10134_/Y _10005_/X _10105_/Y vssd1 vssd1 vccd1 vccd1 _10157_/C
+ sky130_fd_sc_hd__a211o_4
XFILLER_121_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15992_ _15992_/A _15992_/B _15990_/Y vssd1 vssd1 vccd1 vccd1 _15994_/B sky130_fd_sc_hd__or3b_1
XFILLER_122_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10066_ _10198_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10067_/C sky130_fd_sc_hd__xor2_1
X_14943_ _14941_/X _14942_/X _15309_/B vssd1 vssd1 vccd1 vccd1 _14944_/C sky130_fd_sc_hd__a21oi_1
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14874_ _15262_/B _14888_/C _14876_/D vssd1 vssd1 vccd1 vccd1 _14874_/X sky130_fd_sc_hd__or3_2
XFILLER_35_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16613_ _16697_/B _16613_/B vssd1 vssd1 vccd1 vccd1 _16614_/B sky130_fd_sc_hd__nor2_2
X_13825_ _13827_/B _13827_/A vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__nand2b_1
X_17593_ fanout943/X _17593_/D vssd1 vssd1 vccd1 vccd1 _17593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16544_ _16545_/B _16545_/A vssd1 vssd1 vccd1 vccd1 _16544_/X sky130_fd_sc_hd__and2b_1
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13756_ _13757_/B _13756_/B vssd1 vssd1 vccd1 vccd1 _13862_/A sky130_fd_sc_hd__and2b_1
X_10968_ _10969_/B _10969_/A vssd1 vssd1 vccd1 vccd1 _11024_/A sky130_fd_sc_hd__and2b_1
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12707_ _12703_/X _12706_/X _14356_/S vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__mux2_1
X_16475_ _16475_/A _16475_/B vssd1 vssd1 vccd1 vccd1 _16475_/X sky130_fd_sc_hd__or2_4
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _13787_/A _13687_/B vssd1 vssd1 vccd1 vccd1 _13688_/B sky130_fd_sc_hd__and2_2
X_10899_ _10995_/A _10898_/Y _10899_/C _10899_/D vssd1 vssd1 vccd1 vccd1 _10995_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_188_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15426_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15433_/A sky130_fd_sc_hd__xor2_4
X_12638_ _14771_/A _12638_/B vssd1 vssd1 vccd1 vccd1 _12640_/C sky130_fd_sc_hd__nand2_1
XFILLER_157_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ _15774_/A _15397_/A vssd1 vssd1 vccd1 vccd1 _15358_/B sky130_fd_sc_hd__nand2_4
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ _12570_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__nand2_1
XFILLER_157_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14308_ _14309_/B _14309_/A vssd1 vssd1 vccd1 vccd1 _14378_/B sky130_fd_sc_hd__nand2b_2
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15288_ _15278_/A _16136_/B _15216_/A _15213_/X vssd1 vssd1 vccd1 vccd1 _15291_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17027_ _11771_/Y _17025_/Y _17026_/Y vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__a21o_2
X_14239_ _14239_/A _14239_/B vssd1 vssd1 vccd1 vccd1 _14258_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout708 _17498_/Q vssd1 vssd1 vccd1 vccd1 _15101_/A1 sky130_fd_sc_hd__buf_8
Xfanout719 _17497_/Q vssd1 vssd1 vccd1 vccd1 _16480_/A sky130_fd_sc_hd__buf_8
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08800_/X sky130_fd_sc_hd__a21o_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09780_/A _11808_/B _14952_/A vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__and3_1
XFILLER_105_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08731_/A vssd1 vssd1 vccd1 vccd1 _15262_/C sky130_fd_sc_hd__clkinv_4
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09214_ _09214_/A _09214_/B _09214_/C vssd1 vssd1 vccd1 vccd1 _09342_/A sky130_fd_sc_hd__and3_2
XFILLER_33_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09145_ _12176_/A _12129_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09231_/B sky130_fd_sc_hd__and3_1
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ _09076_/A _09076_/B _09076_/C vssd1 vssd1 vccd1 vccd1 _09115_/B sky130_fd_sc_hd__and3_4
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09978_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__nor2_2
XFILLER_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08929_ _08929_/A _08930_/B _08930_/C vssd1 vssd1 vccd1 vccd1 _08929_/Y sky130_fd_sc_hd__nor3_4
XTAP_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11940_ _11941_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11940_/X sky130_fd_sc_hd__and2_2
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11871_ _11871_/A _11871_/B vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__xor2_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13495_/A _13497_/X _13718_/B _13609_/X vssd1 vssd1 vccd1 vccd1 _13612_/A
+ sky130_fd_sc_hd__o211a_2
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _10822_/A _11099_/A vssd1 vssd1 vccd1 vccd1 _10829_/B sky130_fd_sc_hd__nor2_4
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14667_/A _14590_/B vssd1 vssd1 vccd1 vccd1 _14590_/Y sky130_fd_sc_hd__nand2_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _13542_/A sky130_fd_sc_hd__xor2_1
XFILLER_125_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10753_ _15126_/A _10753_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__and3_1
XFILLER_186_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_1036 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16260_ _16352_/A _16352_/B _16259_/C vssd1 vssd1 vccd1 vccd1 _16261_/B sky130_fd_sc_hd__a21oi_1
XFILLER_13_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13472_ _13473_/A _13473_/B vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__and2b_1
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10684_ _10575_/Y _10585_/X _10679_/X _10682_/Y vssd1 vssd1 vccd1 vccd1 _10685_/C
+ sky130_fd_sc_hd__a211o_2
X_15211_ _14881_/X _14889_/X _16410_/A _11841_/A vssd1 vssd1 vccd1 vccd1 _15494_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_127_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _17389_/A _12576_/D _12567_/B _17391_/A vssd1 vssd1 vccd1 vccd1 _12425_/A
+ sky130_fd_sc_hd__a22oi_2
X_16191_ _16191_/A _16191_/B vssd1 vssd1 vccd1 vccd1 _16192_/B sky130_fd_sc_hd__xnor2_2
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15142_ _15069_/A _16317_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _15143_/C sky130_fd_sc_hd__o21a_1
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12354_ _12354_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__xnor2_4
XFILLER_154_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _10962_/A _11370_/C _11370_/D _11240_/A vssd1 vssd1 vccd1 vccd1 _11306_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15073_ _14887_/Y _15071_/Y _14791_/A vssd1 vssd1 vccd1 vccd1 _16315_/B sky130_fd_sc_hd__o21ai_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__a21o_4
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14024_ _14025_/A _14025_/B vssd1 vssd1 vccd1 vccd1 _14119_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11236_ _11146_/B _11143_/C _11143_/D _11144_/A vssd1 vssd1 vccd1 vccd1 _11237_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11167_ _11204_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11167_/X sky130_fd_sc_hd__and2_1
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__xnor2_4
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15975_ _15976_/B _15976_/A vssd1 vssd1 vccd1 vccd1 _15975_/Y sky130_fd_sc_hd__nand2b_1
X_11098_ _11098_/A _11242_/A vssd1 vssd1 vccd1 vccd1 _11101_/B sky130_fd_sc_hd__nor2_4
XFILLER_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10049_ _10053_/A vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__inv_2
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14926_ _16012_/S _14926_/B vssd1 vssd1 vccd1 vccd1 _14926_/X sky130_fd_sc_hd__or2_4
XFILLER_152_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14857_ _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16114_/B sky130_fd_sc_hd__and2_1
XFILLER_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13808_ _13809_/A _13809_/B vssd1 vssd1 vccd1 vccd1 _13923_/A sky130_fd_sc_hd__nor2_2
XFILLER_90_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17576_ fanout925/X _17576_/D vssd1 vssd1 vccd1 vccd1 _17576_/Q sky130_fd_sc_hd__dfxtp_1
X_14788_ _14788_/A _15314_/A vssd1 vssd1 vccd1 vccd1 _14801_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ _13739_/A _13739_/B vssd1 vssd1 vccd1 vccd1 _13741_/C sky130_fd_sc_hd__xnor2_2
XFILLER_177_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16527_ _16527_/A _16527_/B _16527_/C vssd1 vssd1 vccd1 vccd1 _16528_/B sky130_fd_sc_hd__or3_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _16459_/A _16459_/B vssd1 vssd1 vccd1 vccd1 _16550_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15409_ _15501_/A _15418_/B vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__nand2b_4
XFILLER_191_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16389_ _16389_/A _16389_/B _16389_/C vssd1 vssd1 vccd1 vccd1 _16389_/Y sky130_fd_sc_hd__nand3_4
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _10034_/A _09900_/Y _15711_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10042_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_99_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout505 _17518_/Q vssd1 vssd1 vccd1 vccd1 _15396_/A sky130_fd_sc_hd__buf_8
XFILLER_99_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout516 _12104_/A vssd1 vssd1 vccd1 vccd1 _09750_/C sky130_fd_sc_hd__clkbuf_4
X_09832_ _09832_/A _09832_/B vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__nor2_1
Xfanout527 _14667_/A vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__buf_6
Xfanout538 _17515_/Q vssd1 vssd1 vccd1 vccd1 _11322_/A sky130_fd_sc_hd__buf_8
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout549 fanout554/X vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__buf_6
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09763_ _09656_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__o21ai_1
XFILLER_100_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _09695_/A _09693_/Y _10366_/A _10490_/D vssd1 vssd1 vccd1 vccd1 _09842_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_132_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09128_ _09139_/A _09803_/B _09502_/A _09128_/D vssd1 vssd1 vccd1 vccd1 _09139_/B
+ sky130_fd_sc_hd__and4b_2
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09059_ _11900_/B _11870_/B _11867_/C _12107_/A vssd1 vssd1 vccd1 vccd1 _09059_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_68_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_991 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _12237_/A _12645_/B _12070_/C _12070_/D vssd1 vssd1 vccd1 vccd1 _12239_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__or2_2
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ _15760_/A _15760_/B vssd1 vssd1 vccd1 vccd1 _15762_/B sky130_fd_sc_hd__xor2_4
XTAP_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _12972_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _12974_/B sky130_fd_sc_hd__nor2_1
XTAP_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_79_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14736_/A _14744_/B vssd1 vssd1 vccd1 vccd1 _14712_/B sky130_fd_sc_hd__nor2_1
X_11923_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _12179_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _15690_/A _15690_/B _15690_/C vssd1 vssd1 vccd1 vccd1 _15691_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14642_/A _14678_/A vssd1 vssd1 vccd1 vccd1 _14644_/C sky130_fd_sc_hd__nor2_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17430_ input36/X _17607_/Q _17433_/S vssd1 vssd1 vccd1 vccd1 _17607_/D sky130_fd_sc_hd__mux2_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ _13627_/S _16011_/B _11854_/C vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__or3_4
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ _11095_/A _10963_/B _10805_/C _10805_/D vssd1 vssd1 vccd1 vccd1 _10807_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14573_ _14621_/B _14571_/X _14517_/Y _14519_/X vssd1 vssd1 vccd1 vccd1 _14574_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_159_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17361_ _17362_/A _17362_/B _17362_/C _17362_/D vssd1 vssd1 vccd1 vccd1 _17361_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11785_ _09826_/A _14837_/A _12016_/A vssd1 vssd1 vccd1 vccd1 _11785_/X sky130_fd_sc_hd__o21a_1
X_13524_ _13523_/Y _13637_/A _13524_/C vssd1 vssd1 vccd1 vccd1 _13637_/B sky130_fd_sc_hd__nand3b_2
X_16312_ _16298_/A _16806_/A2 _16296_/Y _16311_/X vssd1 vssd1 vccd1 vccd1 _16313_/A
+ sky130_fd_sc_hd__a22o_1
X_17292_ _17574_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__and2_1
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10736_ _11314_/A _11258_/B _10736_/C _10971_/B vssd1 vssd1 vccd1 vccd1 _10739_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16243_ _16149_/X _16153_/B _16245_/A _16040_/B vssd1 vssd1 vccd1 vccd1 _16252_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13455_ _13455_/A _13455_/B _13455_/C vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__or3_1
XFILLER_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ wire120/X _10667_/B _10667_/C vssd1 vssd1 vccd1 vccd1 _10667_/Y sky130_fd_sc_hd__nor3_4
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ _12406_/A _12561_/A vssd1 vssd1 vccd1 vccd1 _12408_/C sky130_fd_sc_hd__nor2_1
XFILLER_173_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16174_ _16174_/A _16174_/B vssd1 vssd1 vccd1 vccd1 _16175_/B sky130_fd_sc_hd__xor2_4
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13386_ _13509_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13388_/B sky130_fd_sc_hd__nand2_1
X_10598_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__or2_2
XFILLER_182_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15125_ _15131_/A _15125_/B vssd1 vssd1 vccd1 vccd1 _15125_/Y sky130_fd_sc_hd__nand2_1
Xoutput108 _17465_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[31] sky130_fd_sc_hd__clkbuf_2
X_12337_ _12657_/B _12338_/C _09647_/B _12657_/A vssd1 vssd1 vccd1 vccd1 _12339_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15056_ _15056_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _15056_/Y sky130_fd_sc_hd__nor2_1
XFILLER_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12268_ _12268_/A _12268_/B _12268_/C vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__and3_2
X_14007_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14008_/C sky130_fd_sc_hd__xnor2_2
X_11219_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11219_/Y sky130_fd_sc_hd__nand2_1
X_12199_ _12198_/A _12198_/B _12198_/C vssd1 vssd1 vccd1 vccd1 _12201_/B sky130_fd_sc_hd__o21ai_4
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput90 _17449_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15958_ _15853_/B _15955_/Y _15957_/X vssd1 vssd1 vccd1 vccd1 _15960_/A sky130_fd_sc_hd__a21o_4
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14909_ _15553_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15820_/A sky130_fd_sc_hd__or2_4
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15889_ _15889_/A _15889_/B vssd1 vssd1 vccd1 vccd1 _15889_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17559_ fanout938/X _17559_/D vssd1 vssd1 vccd1 vccd1 _17559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout302 _15806_/B1 vssd1 vssd1 vccd1 vccd1 _14666_/S sky130_fd_sc_hd__buf_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout313 _17541_/Q vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout324 _17134_/A vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__buf_6
Xfanout335 _12657_/A vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__buf_6
XFILLER_59_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout346 _14766_/A vssd1 vssd1 vccd1 vccd1 _17417_/A sky130_fd_sc_hd__buf_6
X_09815_ _09811_/A _09811_/B _09777_/A vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__a21o_2
Xfanout357 _12487_/A vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__buf_4
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout368 _17411_/A vssd1 vssd1 vccd1 vccd1 _14770_/A sky130_fd_sc_hd__buf_8
Xfanout379 _17533_/Q vssd1 vssd1 vccd1 vccd1 _17409_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_87_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09746_ _09746_/A _09754_/A _09746_/C vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__or3_1
XFILLER_101_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09677_/A vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__clkinv_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11570_ _11526_/B _11552_/X _11557_/X _11603_/A vssd1 vssd1 vccd1 vccd1 _11572_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_168_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ _10437_/A _10437_/B _10437_/C vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13240_ _13241_/A _13241_/B vssd1 vssd1 vccd1 vccd1 _13240_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10452_ _10453_/A _10453_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10454_/A sky130_fd_sc_hd__a21o_2
XFILLER_136_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13171_ _17387_/A _13300_/C vssd1 vssd1 vccd1 vccd1 _13172_/B sky130_fd_sc_hd__nand2_4
X_10383_ _10383_/A _10383_/B _10383_/C vssd1 vssd1 vccd1 vccd1 _10385_/C sky130_fd_sc_hd__nand3_4
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ _12122_/A _12122_/B _12309_/B _12122_/D vssd1 vssd1 vccd1 vccd1 _12122_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_184_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16930_ _16911_/Y _16917_/Y _16929_/X _17170_/B1 _14865_/B vssd1 vssd1 vccd1 vccd1
+ _17568_/D sky130_fd_sc_hd__a32oi_4
X_12053_ _12053_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _12053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11004_ _11157_/A _11002_/Y _10941_/Y _10946_/X vssd1 vssd1 vccd1 vccd1 _11055_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16861_ _16792_/A _16792_/B _16788_/Y vssd1 vssd1 vccd1 vccd1 _16863_/B sky130_fd_sc_hd__a21o_2
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout880 _17480_/Q vssd1 vssd1 vccd1 vccd1 _17302_/A1 sky130_fd_sc_hd__buf_6
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout891 _11506_/C vssd1 vssd1 vccd1 vccd1 _14794_/B sky130_fd_sc_hd__buf_4
X_15812_ _16015_/A _15898_/B _15811_/Y _15810_/X vssd1 vssd1 vccd1 vccd1 _15812_/X
+ sky130_fd_sc_hd__o31a_1
X_16792_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _16793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15743_ _15743_/A _15743_/B vssd1 vssd1 vccd1 vccd1 _15765_/A sky130_fd_sc_hd__xor2_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _12954_/B _12955_/B vssd1 vssd1 vccd1 vccd1 _12956_/B sky130_fd_sc_hd__nand2b_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _11906_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__xnor2_1
XFILLER_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15674_ _15675_/A _15675_/B vssd1 vssd1 vccd1 vccd1 _15674_/X sky130_fd_sc_hd__and2_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12886_/A _12886_/B _12886_/C vssd1 vssd1 vccd1 vccd1 _12899_/B sky130_fd_sc_hd__or3_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17413_/A _17419_/B vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__or2_1
XFILLER_178_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14625_ _14660_/B _14625_/B vssd1 vssd1 vccd1 vccd1 _14627_/C sky130_fd_sc_hd__nor2_1
X_11837_ _14912_/B _11837_/B vssd1 vssd1 vccd1 vccd1 _11837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14556_ _14557_/A _14557_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14558_/A sky130_fd_sc_hd__o21a_1
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _12567_/B _17354_/A2 _17343_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17501_/D
+ sky130_fd_sc_hd__o211a_1
X_11768_ _11768_/A _11768_/B vssd1 vssd1 vccd1 vccd1 _16921_/A sky130_fd_sc_hd__or2_1
XFILLER_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10719_ _10720_/A _10718_/Y _10962_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _11013_/A
+ sky130_fd_sc_hd__and4bb_4
X_13507_ _13619_/A _13507_/B vssd1 vssd1 vccd1 vccd1 _13514_/A sky130_fd_sc_hd__nand2_1
X_14487_ _14676_/A _14545_/C vssd1 vssd1 vccd1 vccd1 _14489_/B sky130_fd_sc_hd__nand2_1
X_17275_ _17459_/Q _17293_/A2 _17273_/X _17274_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17459_/D sky130_fd_sc_hd__o221a_1
XFILLER_186_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ _11586_/A _11586_/C _11620_/A vssd1 vssd1 vccd1 vccd1 _11700_/C sky130_fd_sc_hd__a21o_1
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16226_ _16880_/A _16226_/B _16226_/C _17119_/C vssd1 vssd1 vccd1 vccd1 _16227_/B
+ sky130_fd_sc_hd__and4_2
X_13438_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13439_/B sky130_fd_sc_hd__and2_1
X_16157_ _16157_/A _16157_/B vssd1 vssd1 vccd1 vccd1 _16158_/B sky130_fd_sc_hd__xnor2_4
X_13369_ _13369_/A _13369_/B _13369_/C vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__and3_2
XFILLER_170_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15108_ _15108_/A _15108_/B vssd1 vssd1 vccd1 vccd1 _15108_/Y sky130_fd_sc_hd__nand2_1
X_16088_ _16197_/B _16088_/B vssd1 vssd1 vccd1 vccd1 _16089_/B sky130_fd_sc_hd__or2_4
XFILLER_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15039_ _15038_/A _14956_/Y _15038_/Y _15097_/A vssd1 vssd1 vccd1 vccd1 _15039_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09600_ _09580_/X _09597_/B _09599_/Y _09480_/X vssd1 vssd1 vccd1 vccd1 _09629_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _09485_/X _09530_/X _09393_/X _09398_/Y vssd1 vssd1 vccd1 vccd1 _09531_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09462_ _09462_/A _09468_/A _09462_/C vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__or3_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09393_ _09395_/B _09393_/B _09393_/C _09393_/D vssd1 vssd1 vccd1 vccd1 _09393_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout132 _16152_/A vssd1 vssd1 vccd1 vccd1 _16760_/B sky130_fd_sc_hd__buf_6
Xfanout143 _15020_/X vssd1 vssd1 vccd1 vccd1 _15821_/A sky130_fd_sc_hd__buf_6
Xfanout154 _14890_/Y vssd1 vssd1 vccd1 vccd1 _16056_/A sky130_fd_sc_hd__buf_6
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout165 _17296_/Y vssd1 vssd1 vccd1 vccd1 _17360_/A2 sky130_fd_sc_hd__buf_4
Xfanout176 _15575_/Y vssd1 vssd1 vccd1 vccd1 _15774_/B sky130_fd_sc_hd__buf_4
XFILLER_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout187 _15327_/X vssd1 vssd1 vccd1 vccd1 _15752_/B sky130_fd_sc_hd__buf_6
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout198 _17164_/C vssd1 vssd1 vccd1 vccd1 _16582_/A sky130_fd_sc_hd__buf_4
XFILLER_75_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _11900_/B _10036_/D _10645_/C _12107_/A vssd1 vssd1 vccd1 vccd1 _09729_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12740_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12903_/B sky130_fd_sc_hd__and2b_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12671_ _12671_/A _12671_/B vssd1 vssd1 vccd1 vccd1 _12673_/B sky130_fd_sc_hd__xnor2_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14473_/A _14409_/C _14409_/A vssd1 vssd1 vccd1 vccd1 _14411_/B sky130_fd_sc_hd__a21o_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _11622_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _15614_/A sky130_fd_sc_hd__or2_1
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/A _15390_/B vssd1 vssd1 vccd1 vccd1 _15390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341_ _14340_/B _14340_/C _14340_/A vssd1 vssd1 vccd1 vccd1 _14342_/B sky130_fd_sc_hd__a21o_1
XFILLER_184_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ _11553_/A _11553_/B _14794_/B _11553_/D vssd1 vssd1 vccd1 vccd1 _11637_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17060_ _17060_/A _17060_/B vssd1 vssd1 vccd1 vccd1 _17062_/B sky130_fd_sc_hd__nor2_1
X_10504_ _10508_/C _10933_/D _10395_/A _10393_/Y vssd1 vssd1 vccd1 vccd1 _10505_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14272_ _14273_/A _14273_/B _14273_/C vssd1 vssd1 vccd1 vccd1 _14350_/B sky130_fd_sc_hd__a21oi_2
XFILLER_155_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11484_ _11484_/A _11484_/B _11522_/A vssd1 vssd1 vccd1 vccd1 _11485_/B sky130_fd_sc_hd__or3_1
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16011_ _16011_/A _16011_/B _16011_/C vssd1 vssd1 vccd1 vccd1 _16011_/X sky130_fd_sc_hd__or3_4
XFILLER_183_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13223_ _16649_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10435_ _10436_/B _10436_/A vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__and2b_1
XFILLER_137_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _13154_/A _13154_/B vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ _10366_/A _17467_/D _10709_/A vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__and3_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__xnor2_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13085_ _13085_/A _13085_/B _13085_/C vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__or3_1
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10297_ _10419_/A _10532_/B _10755_/D _10534_/D vssd1 vssd1 vccd1 vccd1 _10300_/A
+ sky130_fd_sc_hd__and4_1
X_16913_ _14865_/B _17134_/C _16913_/C vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__and3b_1
X_12036_ _12865_/S _12034_/X _12035_/X vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__o21ai_4
XFILLER_144_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16844_ _16906_/B _16844_/B vssd1 vssd1 vccd1 vccd1 _16846_/C sky130_fd_sc_hd__and2_1
XFILLER_66_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1006 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16775_ _16775_/A _16775_/B vssd1 vssd1 vccd1 vccd1 _16777_/C sky130_fd_sc_hd__xnor2_1
X_13987_ _13988_/A _13988_/B vssd1 vssd1 vccd1 vccd1 _14077_/A sky130_fd_sc_hd__nor2_4
XFILLER_46_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15726_ _15726_/A _15918_/A _16745_/B _15726_/D vssd1 vssd1 vccd1 vccd1 _15834_/A
+ sky130_fd_sc_hd__and4_4
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12938_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__and3_2
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _15703_/A _15658_/B vssd1 vssd1 vccd1 vccd1 _15749_/B sky130_fd_sc_hd__and2_4
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _17399_/A _13566_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__and3_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14608_ _14609_/A _14609_/B vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__nor2_2
X_15588_ _15588_/A _15588_/B vssd1 vssd1 vccd1 vccd1 _15590_/C sky130_fd_sc_hd__xnor2_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327_ input42/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17327_/X sky130_fd_sc_hd__or3_1
X_14539_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14585_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_179_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_978 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _17595_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17258_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16209_ _14859_/B _16209_/B _16209_/C vssd1 vssd1 vccd1 vccd1 _16210_/B sky130_fd_sc_hd__and3b_1
XFILLER_127_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17189_ input30/X input34/X input5/X input4/X vssd1 vssd1 vccd1 vccd1 _17191_/C sky130_fd_sc_hd__or4_1
XFILLER_161_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08962_ _08962_/A _08962_/B _08962_/C vssd1 vssd1 vccd1 vccd1 _08985_/B sky130_fd_sc_hd__and3_1
XFILLER_142_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08893_ _08893_/A _08893_/B vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__xnor2_4
XFILLER_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _11953_/A _09637_/B _09947_/B _10067_/B vssd1 vssd1 vccd1 vccd1 _09517_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_65_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _11900_/B _11867_/D _11859_/C _09584_/A vssd1 vssd1 vccd1 vccd1 _09445_/Y
+ sky130_fd_sc_hd__a22oi_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09376_ _09942_/A _09637_/B _09803_/B _09947_/B vssd1 vssd1 vccd1 vccd1 _09379_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _10219_/A _10342_/A vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__and2b_2
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__nor2_2
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _10209_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__nand2_2
XFILLER_102_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13910_ _14027_/B _13910_/B vssd1 vssd1 vccd1 vccd1 _13912_/B sky130_fd_sc_hd__or2_1
XFILLER_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14890_ _14881_/X _14889_/X _08723_/Y vssd1 vssd1 vccd1 vccd1 _14890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13841_ _13841_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _13841_/X sky130_fd_sc_hd__or2_1
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwb_buttons_leds_951 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_951/HI led_enb[4] sky130_fd_sc_hd__conb_1
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16560_ _16560_/A _16560_/B vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__nand2_2
X_13772_ _14153_/B _14141_/D _14050_/D _14153_/A vssd1 vssd1 vccd1 vccd1 _13774_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10984_ _10984_/A _10985_/A _10984_/C vssd1 vssd1 vccd1 vccd1 _11162_/A sky130_fd_sc_hd__or3_2
XFILLER_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15511_ _15512_/A _15512_/B vssd1 vssd1 vccd1 vccd1 _15511_/X sky130_fd_sc_hd__and2b_1
XFILLER_71_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ _12723_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _12725_/A sky130_fd_sc_hd__nor2_1
XFILLER_188_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16491_ _16735_/A _14127_/X _16582_/A _15104_/X vssd1 vssd1 vccd1 vccd1 _16492_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12655_/B sky130_fd_sc_hd__nand2_1
X_15442_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15442_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_188_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _15305_/C _11605_/B _11610_/B _11605_/D vssd1 vssd1 vccd1 vccd1 _11607_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_157_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12585_ _12585_/A _12585_/B _12585_/C vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__and3_1
X_15373_ _14896_/B _15373_/B _15373_/C vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__and3b_1
XFILLER_157_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17112_ _17164_/A _16582_/A _15252_/X _16653_/A _14705_/B vssd1 vssd1 vccd1 vccd1
+ _17113_/C sky130_fd_sc_hd__o32a_1
X_14324_ _14324_/A _14389_/B _14325_/B vssd1 vssd1 vccd1 vccd1 _14393_/A sky130_fd_sc_hd__or3_1
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _11532_/A _11532_/B _11574_/A vssd1 vssd1 vccd1 vccd1 _11537_/C sky130_fd_sc_hd__o21ba_2
XFILLER_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14255_ _14255_/A _14255_/B vssd1 vssd1 vccd1 vccd1 _14258_/B sky130_fd_sc_hd__xnor2_2
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17043_ _17119_/A _17043_/B _17043_/C vssd1 vssd1 vccd1 vccd1 _17085_/B sky130_fd_sc_hd__and3_1
XFILLER_99_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap118 _11949_/Y vssd1 vssd1 vccd1 vccd1 _11998_/A sky130_fd_sc_hd__buf_4
X_11467_ _11506_/A _11553_/A _15401_/A _11506_/C vssd1 vssd1 vccd1 vccd1 _11472_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_171_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _16644_/C _16651_/A vssd1 vssd1 vccd1 vccd1 _16649_/A sky130_fd_sc_hd__nand2_4
X_10418_ _10418_/A _10423_/A _10418_/C vssd1 vssd1 vccd1 vccd1 _10427_/B sky130_fd_sc_hd__or3_4
XFILLER_87_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ _14186_/A _14186_/B vssd1 vssd1 vccd1 vccd1 _14188_/C sky130_fd_sc_hd__or2_2
X_11398_ _11403_/A _11368_/Y _11384_/Y _11396_/X vssd1 vssd1 vccd1 vccd1 _11400_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13137_/A _13137_/B vssd1 vssd1 vccd1 vccd1 _13268_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__and2_1
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _12021_/A _15101_/A1 _14956_/A vssd1 vssd1 vccd1 vccd1 _12020_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16827_ _16827_/A _16827_/B _16827_/C _16827_/D vssd1 vssd1 vccd1 vccd1 _16828_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_94_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16758_ _16758_/A _16758_/B _16758_/C vssd1 vssd1 vccd1 vccd1 _16759_/B sky130_fd_sc_hd__and3_1
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15709_ _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15710_/C sky130_fd_sc_hd__nor2_1
X_16689_ _16690_/A _16690_/B vssd1 vssd1 vccd1 vccd1 _16770_/B sky130_fd_sc_hd__and2b_1
XFILLER_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09230_ _09230_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__xnor2_4
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09161_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09161_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09092_ _09092_/A vssd1 vssd1 vccd1 vccd1 _09093_/B sky130_fd_sc_hd__inv_2
XFILLER_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09994_ _09994_/A _16809_/B vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__xnor2_4
XFILLER_103_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08945_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__xnor2_2
XFILLER_192_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08876_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__xnor2_2
XFILLER_96_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ _10904_/B _09428_/B vssd1 vssd1 vccd1 vccd1 _16990_/B sky130_fd_sc_hd__nand2_4
XFILLER_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09359_ _09366_/A _09366_/B _09366_/C vssd1 vssd1 vccd1 vccd1 _09370_/B sky130_fd_sc_hd__a21o_1
XFILLER_166_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ _12370_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__xnor2_4
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _14790_/A _15175_/B vssd1 vssd1 vccd1 vccd1 _11321_/X sky130_fd_sc_hd__and2_1
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14040_ _13950_/A _13948_/C _13745_/D _13948_/A vssd1 vssd1 vccd1 vccd1 _14040_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11252_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__xnor2_4
XFILLER_181_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10203_ _10559_/A _10805_/C _10203_/C vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__and3_1
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _11182_/A _11182_/B _11182_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__o21a_2
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10134_ _10134_/A _10134_/B _10134_/C vssd1 vssd1 vccd1 vccd1 _10134_/Y sky130_fd_sc_hd__nand3_4
X_15991_ _15992_/A _15992_/B _15990_/Y vssd1 vssd1 vccd1 vccd1 _15991_/X sky130_fd_sc_hd__o21ba_2
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ _10198_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__and2_2
X_14942_ _14942_/A _15553_/A _15891_/B vssd1 vssd1 vccd1 vccd1 _14942_/X sky130_fd_sc_hd__or3_1
XFILLER_0_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14873_ _15069_/A _16317_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _14876_/D sky130_fd_sc_hd__or3b_2
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16612_ _16611_/B _16612_/B vssd1 vssd1 vccd1 vccd1 _16613_/B sky130_fd_sc_hd__and2b_1
X_13824_ _13824_/A _13824_/B vssd1 vssd1 vccd1 vccd1 _13827_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17592_ fanout944/X _17592_/D vssd1 vssd1 vccd1 vccd1 _17592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16543_ _16543_/A _16543_/B vssd1 vssd1 vccd1 vccd1 _16545_/B sky130_fd_sc_hd__xnor2_1
X_13755_ _13650_/B _13652_/B _13648_/X vssd1 vssd1 vccd1 vccd1 _13757_/B sky130_fd_sc_hd__a21oi_1
X_10967_ _10915_/A _10914_/B _10914_/A vssd1 vssd1 vccd1 vccd1 _10969_/B sky130_fd_sc_hd__o21ba_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12704_/X _12705_/X _13627_/S vssd1 vssd1 vccd1 vccd1 _12706_/X sky130_fd_sc_hd__mux2_1
X_16474_ _16563_/A _16384_/Y _16472_/X _15523_/A vssd1 vssd1 vccd1 vccd1 _16475_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13686_ _13686_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13687_/B sky130_fd_sc_hd__nand2_1
X_10898_ _14922_/S _10791_/C _10897_/C vssd1 vssd1 vccd1 vccd1 _10898_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15425_ _15426_/A _15426_/B vssd1 vssd1 vccd1 vccd1 _15514_/A sky130_fd_sc_hd__nand2_1
XFILLER_188_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12637_ _14769_/A _14770_/A _12637_/C _12637_/D vssd1 vssd1 vccd1 vccd1 _12792_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_141_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12568_ _12568_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__xnor2_4
X_15356_ _15356_/A _15356_/B vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__nand2_4
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14307_ _14225_/A _16970_/A _14225_/B vssd1 vssd1 vccd1 vccd1 _14309_/B sky130_fd_sc_hd__o21ba_1
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11519_ _11561_/B _11518_/C _11563_/D _11629_/A vssd1 vssd1 vccd1 vccd1 _11519_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_176_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12499_ _12499_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12501_/A sky130_fd_sc_hd__nor2_2
X_15287_ _15287_/A _15287_/B vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__xor2_4
XFILLER_171_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17026_ _11771_/Y _17025_/Y _16922_/A vssd1 vssd1 vccd1 vccd1 _17026_/Y sky130_fd_sc_hd__o21ai_1
X_14238_ _14237_/A _14237_/B _14236_/X vssd1 vssd1 vccd1 vccd1 _14239_/B sky130_fd_sc_hd__o21ba_1
XFILLER_176_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14169_ _14170_/A _14245_/A _14170_/C vssd1 vssd1 vccd1 vccd1 _14171_/A sky130_fd_sc_hd__o21a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout709 _13564_/D vssd1 vssd1 vccd1 vccd1 _14141_/D sky130_fd_sc_hd__buf_6
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ input70/X vssd1 vssd1 vccd1 vccd1 _08730_/Y sky130_fd_sc_hd__clkinv_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09213_ _09213_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09214_/C sky130_fd_sc_hd__xnor2_1
XFILLER_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09144_ _12176_/A _12129_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09147_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_108_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ _09076_/A _09076_/B _09076_/C vssd1 vssd1 vccd1 vccd1 _09115_/A sky130_fd_sc_hd__a21oi_4
XFILLER_190_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09977_ _10366_/A _10479_/B _09841_/A _09839_/Y vssd1 vssd1 vccd1 vccd1 _09983_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08928_ _08832_/Y _08875_/X _08905_/A _09051_/A vssd1 vssd1 vccd1 vccd1 _08930_/C
+ sky130_fd_sc_hd__o211a_4
XTAP_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08859_ _08859_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11870_ _12245_/A _11870_/B _11871_/A vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__and3_2
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _10822_/A _10820_/Y _14785_/A _10957_/D vssd1 vssd1 vccd1 vccd1 _11099_/A
+ sky130_fd_sc_hd__and4bb_4
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13540_ _13658_/A _13948_/C _13657_/B vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__and3_1
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _11629_/B _10993_/D vssd1 vssd1 vccd1 vccd1 _10897_/C sky130_fd_sc_hd__and2_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13471_ _13471_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__xnor2_2
XFILLER_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10683_ _10679_/X _10682_/Y _10575_/Y _10585_/X vssd1 vssd1 vccd1 vccd1 _10685_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15210_ _15203_/X _15208_/X _15238_/A vssd1 vssd1 vccd1 vccd1 _15932_/B sky130_fd_sc_hd__a21bo_4
XFILLER_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12422_ _12257_/A _12259_/B _12257_/B vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__o21ba_4
X_16190_ _16281_/A _16533_/B vssd1 vssd1 vccd1 vccd1 _16191_/B sky130_fd_sc_hd__nand2_2
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15141_ _15270_/A _15141_/B vssd1 vssd1 vccd1 vccd1 _15393_/B sky130_fd_sc_hd__or2_4
X_12353_ _12353_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _12354_/B sky130_fd_sc_hd__and2_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11304_ _11304_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__nor2_2
XFILLER_154_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15072_ _14887_/Y _15071_/Y _14791_/A vssd1 vssd1 vccd1 vccd1 _16127_/B sky130_fd_sc_hd__o21a_2
X_12284_ _12284_/A _12284_/B vssd1 vssd1 vccd1 vccd1 _12286_/C sky130_fd_sc_hd__or2_2
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14023_ _13809_/A _13809_/B _13923_/B _13922_/A vssd1 vssd1 vccd1 vccd1 _14025_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11235_ _11153_/B _11151_/C _11151_/B vssd1 vssd1 vccd1 vccd1 _11235_/X sky130_fd_sc_hd__o21a_2
XFILLER_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11166_ _11165_/A _11165_/B _11165_/C vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__o21ai_1
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _11026_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__nand2_4
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15974_ _15840_/Y _15864_/B _15839_/Y vssd1 vssd1 vccd1 vccd1 _15976_/B sky130_fd_sc_hd__a21oi_4
X_11097_ _11098_/A _11096_/Y _14785_/A _11097_/D vssd1 vssd1 vccd1 vccd1 _11242_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10048_ _10050_/B _10163_/A _10050_/A vssd1 vssd1 vccd1 vccd1 _10053_/A sky130_fd_sc_hd__a21o_2
X_14925_ _16012_/S _14926_/B vssd1 vssd1 vccd1 vccd1 _14925_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14856_ _15898_/A _15811_/A _15811_/B vssd1 vssd1 vccd1 vccd1 _16014_/B sky130_fd_sc_hd__and3_1
XFILLER_64_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _13688_/A _13688_/B _13706_/Y vssd1 vssd1 vccd1 vccd1 _13809_/B sky130_fd_sc_hd__a21boi_2
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17575_ fanout926/X _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/Q sky130_fd_sc_hd__dfxtp_1
X_14787_ _14787_/A _15381_/A vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__nor2_2
X_11999_ _11998_/A _11998_/B _12197_/B _11998_/D vssd1 vssd1 vccd1 vccd1 _11999_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_32_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16526_ _16527_/A _16527_/B _16527_/C vssd1 vssd1 vccd1 vccd1 _16630_/A sky130_fd_sc_hd__o21ai_4
XFILLER_188_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13738_ _13950_/A _13844_/D _13739_/A vssd1 vssd1 vccd1 vccd1 _13849_/B sky130_fd_sc_hd__and3_1
XFILLER_56_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16457_ _16457_/A _16457_/B vssd1 vssd1 vccd1 vccd1 _16459_/B sky130_fd_sc_hd__xnor2_1
X_13669_ _13778_/B _13669_/B vssd1 vssd1 vccd1 vccd1 _13671_/C sky130_fd_sc_hd__nor2_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ _15408_/A _15408_/B _15408_/C vssd1 vssd1 vccd1 vccd1 _15418_/B sky130_fd_sc_hd__or3_4
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16388_ _16387_/B _16387_/C _16387_/A vssd1 vssd1 vccd1 vccd1 _16389_/C sky130_fd_sc_hd__o21ai_4
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15339_ _15206_/X _15338_/Y _14896_/B vssd1 vssd1 vccd1 vccd1 _15755_/B sky130_fd_sc_hd__o21ai_4
XFILLER_184_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_929 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17009_ _17037_/A _17009_/B vssd1 vssd1 vccd1 vccd1 _17010_/B sky130_fd_sc_hd__nand2_2
X_09900_ _10171_/B _10543_/B _10657_/B _14789_/A vssd1 vssd1 vccd1 vccd1 _09900_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_132_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout506 _12592_/B vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__clkbuf_8
X_09831_ _09740_/A _09740_/B _09740_/C vssd1 vssd1 vccd1 vccd1 _09832_/B sky130_fd_sc_hd__a21oi_1
Xfanout517 _12442_/A vssd1 vssd1 vccd1 vccd1 _12104_/A sky130_fd_sc_hd__buf_6
XFILLER_101_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout528 _15457_/A vssd1 vssd1 vccd1 vccd1 _14667_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout539 _09470_/B vssd1 vssd1 vccd1 vccd1 _11930_/B sky130_fd_sc_hd__buf_6
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09762_ _09762_/A _09762_/B _09891_/A vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__nand3_2
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09693_ _10235_/A _10490_/C _10479_/B _10236_/A vssd1 vssd1 vccd1 vccd1 _09693_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_55_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_182_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09127_ _12174_/A _12174_/B _12127_/D _11920_/D vssd1 vssd1 vccd1 vccd1 _09139_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_163_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09058_ _12107_/A _11900_/B _13088_/B _11867_/C vssd1 vssd1 vccd1 vccd1 _09061_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_151_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_940 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11020_ _11020_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__xnor2_4
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12971_ _12971_/A _12971_/B vssd1 vssd1 vccd1 vccd1 _12974_/A sky130_fd_sc_hd__xor2_1
XTAP_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14719_/A _14710_/B _14710_/C vssd1 vssd1 vccd1 vccd1 _14744_/B sky130_fd_sc_hd__and3b_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _12772_/A _12127_/C vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _15690_/A _15690_/B _15690_/C vssd1 vssd1 vccd1 vccd1 _15779_/B sky130_fd_sc_hd__or3_4
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14641_ _14738_/A _14708_/B _14641_/C _14641_/D vssd1 vssd1 vccd1 vccd1 _14678_/A
+ sky130_fd_sc_hd__and4_2
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _14840_/A _13626_/B vssd1 vssd1 vccd1 vccd1 _11853_/Y sky130_fd_sc_hd__nand2_2
XFILLER_82_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17360_ _13947_/B _17360_/A2 _17359_/X _17426_/C1 vssd1 vssd1 vccd1 vccd1 _17509_/D
+ sky130_fd_sc_hd__o211a_1
X_10804_ _10962_/A _10912_/C vssd1 vssd1 vccd1 vccd1 _10808_/A sky130_fd_sc_hd__nand2_4
X_14572_ _14517_/Y _14519_/X _14621_/B _14571_/X vssd1 vssd1 vccd1 vccd1 _14624_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _14872_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__or2_1
XFILLER_186_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16311_ _14836_/A _16293_/Y _16301_/Y _17156_/B _16310_/X vssd1 vssd1 vccd1 vccd1
+ _16311_/X sky130_fd_sc_hd__o221a_1
X_13523_ _14775_/A _13523_/B vssd1 vssd1 vccd1 vccd1 _13523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17291_ _17606_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17291_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _10735_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _10750_/A sky130_fd_sc_hd__xnor2_2
XFILLER_186_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16242_ _16347_/A _16242_/B vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__nand2b_4
XFILLER_40_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13454_ _13454_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13455_/C sky130_fd_sc_hd__nor2_1
X_10666_ _10519_/Y _10588_/X _10632_/A _10632_/Y vssd1 vssd1 vccd1 vccd1 _10667_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_185_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ _17403_/A _17399_/A _13450_/D _13866_/D vssd1 vssd1 vccd1 vccd1 _12561_/A
+ sky130_fd_sc_hd__and4_1
X_16173_ _16171_/A _16814_/B _16066_/A _16064_/A vssd1 vssd1 vccd1 vccd1 _16174_/B
+ sky130_fd_sc_hd__a31o_4
X_13385_ _13509_/B _13385_/B vssd1 vssd1 vccd1 vccd1 _13508_/B sky130_fd_sc_hd__nor2_1
X_10597_ _10597_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10599_/B sky130_fd_sc_hd__xnor2_4
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_86_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15124_ _15709_/A _10013_/B _09712_/B _10897_/B _14942_/A _10993_/C vssd1 vssd1 vccd1
+ vccd1 _15125_/B sky130_fd_sc_hd__mux4_1
Xoutput109 _17437_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[3] sky130_fd_sc_hd__clkbuf_2
X_12336_ _12336_/A _12336_/B vssd1 vssd1 vccd1 vccd1 _12354_/A sky130_fd_sc_hd__nor2_4
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12267_ _12268_/A _12268_/B _12268_/C vssd1 vssd1 vccd1 vccd1 _12267_/Y sky130_fd_sc_hd__a21oi_4
X_15055_ _14790_/A _16735_/A _12063_/X _15054_/X vssd1 vssd1 vccd1 vccd1 _15055_/X
+ sky130_fd_sc_hd__o31a_1
X_14006_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14115_/A sky130_fd_sc_hd__nand2b_1
X_11218_ _11218_/A _11218_/B vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__nand2_4
XFILLER_141_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12198_ _12198_/A _12198_/B _12198_/C vssd1 vssd1 vccd1 vccd1 _12367_/B sky130_fd_sc_hd__or3_4
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput80 _17473_/Q vssd1 vssd1 vccd1 vccd1 leds[7] sky130_fd_sc_hd__clkbuf_2
Xoutput91 _17450_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_150_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11149_ _11154_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _11151_/B sky130_fd_sc_hd__nand2_2
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15957_ _16619_/A _16041_/A _16062_/C vssd1 vssd1 vccd1 vccd1 _15957_/X sky130_fd_sc_hd__o21ba_1
XFILLER_64_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ _15553_/A _15553_/B vssd1 vssd1 vccd1 vccd1 _15475_/A sky130_fd_sc_hd__nor2_8
XFILLER_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15888_ _15888_/A _15888_/B vssd1 vssd1 vccd1 vccd1 _15889_/B sky130_fd_sc_hd__nand2_2
XFILLER_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14839_ _14839_/A _14839_/B vssd1 vssd1 vccd1 vccd1 _14839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17558_ fanout939/X _17558_/D vssd1 vssd1 vccd1 vccd1 _17558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_189_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16509_ _16509_/A _16509_/B _16509_/C vssd1 vssd1 vccd1 vccd1 _16510_/B sky130_fd_sc_hd__and3_1
XFILLER_149_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17489_ fanout931/X _17489_/D vssd1 vssd1 vccd1 vccd1 _17489_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_177_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout303 _15175_/A vssd1 vssd1 vccd1 vccd1 _15806_/B1 sky130_fd_sc_hd__buf_4
Xfanout314 _17541_/Q vssd1 vssd1 vccd1 vccd1 _12618_/A sky130_fd_sc_hd__buf_4
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout325 _17134_/A vssd1 vssd1 vccd1 vccd1 _14050_/B sky130_fd_sc_hd__buf_6
Xfanout336 _12657_/A vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__buf_2
X_09814_ _09772_/X _09813_/X _09668_/Y _09683_/X vssd1 vssd1 vccd1 vccd1 _09814_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout347 _17537_/Q vssd1 vssd1 vccd1 vccd1 _14766_/A sky130_fd_sc_hd__buf_6
XFILLER_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout358 _12487_/A vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__buf_8
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout369 _17534_/Q vssd1 vssd1 vccd1 vccd1 _17411_/A sky130_fd_sc_hd__buf_6
XFILLER_101_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09745_ _09621_/X _09743_/Y _09740_/B _09724_/X vssd1 vssd1 vccd1 vccd1 _09745_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09678_/B _09681_/A _09678_/A vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10520_ _10519_/A _10519_/Y _10406_/B _10474_/Y vssd1 vssd1 vccd1 vccd1 _10555_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_168_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10451_ _10451_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10453_/C sky130_fd_sc_hd__or2_1
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13170_ _13170_/A _13170_/B vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__nor2_2
X_10382_ _10382_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__xnor2_2
XFILLER_151_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ _12122_/A _12122_/B _12309_/B _12122_/D vssd1 vssd1 vccd1 vccd1 _12121_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_124_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12052_ _12021_/A _09892_/D _10991_/C vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__a21o_1
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11003_ _10941_/Y _10946_/X _11157_/A _11002_/Y vssd1 vssd1 vccd1 vccd1 _11157_/B
+ sky130_fd_sc_hd__o211ai_4
X_16860_ _14383_/A _16859_/Y _16858_/Y vssd1 vssd1 vccd1 vccd1 _16863_/A sky130_fd_sc_hd__a21oi_4
Xfanout870 _10360_/D vssd1 vssd1 vccd1 vccd1 _17469_/D sky130_fd_sc_hd__buf_6
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15811_ _15811_/A _15811_/B vssd1 vssd1 vccd1 vccd1 _15811_/Y sky130_fd_sc_hd__nor2_1
Xfanout881 _10809_/D vssd1 vssd1 vccd1 vccd1 _17468_/D sky130_fd_sc_hd__buf_4
X_16791_ _16791_/A _16791_/B vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__nand2_1
Xfanout892 _15008_/A vssd1 vssd1 vccd1 vccd1 _11506_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15742_ _15742_/A _15742_/B _15743_/B vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__nor3_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _12955_/B _12954_/B vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__nand2b_2
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _11906_/B _11906_/A vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__and2b_2
X_15673_ _15673_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15675_/B sky130_fd_sc_hd__xnor2_2
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12886_/A _12886_/B _12886_/C vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__o21ai_4
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ input52/X _17422_/A2 _17411_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17534_/D
+ sky130_fd_sc_hd__o211a_1
X_14624_ _14624_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14625_/B sky130_fd_sc_hd__and2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _09712_/B _12659_/B _11839_/S vssd1 vssd1 vccd1 vccd1 _11837_/B sky130_fd_sc_hd__mux2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ input51/X _17355_/B _17355_/C vssd1 vssd1 vccd1 vccd1 _17343_/X sky130_fd_sc_hd__or3_1
X_14555_ _14555_/A _14555_/B vssd1 vssd1 vccd1 vccd1 _14557_/C sky130_fd_sc_hd__xnor2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11767_ _11768_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11767_/X sky130_fd_sc_hd__or2_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13506_ _13506_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13507_/B sky130_fd_sc_hd__or2_1
X_17274_ _17568_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17274_/X sky130_fd_sc_hd__and2_1
X_10718_ _10963_/B _10962_/B _10963_/C _10963_/A vssd1 vssd1 vccd1 vccd1 _10718_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_186_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14486_ _14486_/A _14557_/A vssd1 vssd1 vccd1 vccd1 _14489_/A sky130_fd_sc_hd__or2_1
XFILLER_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11698_ _11622_/B _15614_/B _11622_/A vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__o21bai_2
X_16225_ _16315_/B _16827_/C _16409_/B _15734_/A vssd1 vssd1 vccd1 vccd1 _16227_/A
+ sky130_fd_sc_hd__o22a_1
X_13437_ _13438_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__nor2_2
X_10649_ _10649_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _10735_/B sky130_fd_sc_hd__xnor2_4
XFILLER_139_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16156_ _16157_/B _16157_/A vssd1 vssd1 vccd1 vccd1 _16270_/B sky130_fd_sc_hd__and2b_1
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13369_/C sky130_fd_sc_hd__or2_2
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15107_ _11472_/B _14791_/X _14797_/X vssd1 vssd1 vccd1 vccd1 _15108_/B sky130_fd_sc_hd__a21o_1
X_12319_ _12487_/B _12659_/B _13194_/D _12487_/A vssd1 vssd1 vccd1 vccd1 _12323_/A
+ sky130_fd_sc_hd__a22oi_4
X_16087_ _16281_/A _16355_/B _16086_/C vssd1 vssd1 vccd1 vccd1 _16088_/B sky130_fd_sc_hd__a21oi_1
X_13299_ _13658_/A _13948_/D _13657_/B vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__a21boi_4
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15038_ _15038_/A _15038_/B vssd1 vssd1 vccd1 vccd1 _15038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16989_ _16989_/A _16989_/B vssd1 vssd1 vccd1 vccd1 _16991_/C sky130_fd_sc_hd__or2_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09530_ _09485_/X _09530_/B _09530_/C _09530_/D vssd1 vssd1 vccd1 vccd1 _09530_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _09335_/A _09459_/Y _09455_/B _09440_/X vssd1 vssd1 vccd1 vccd1 _09461_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_64_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09395_/B _09392_/B _09393_/C _09393_/D vssd1 vssd1 vccd1 vccd1 _09395_/C
+ sky130_fd_sc_hd__nor4_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout133 _15755_/B vssd1 vssd1 vccd1 vccd1 _16041_/A sky130_fd_sc_hd__buf_12
XFILLER_59_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout144 _16165_/A vssd1 vssd1 vccd1 vccd1 _15278_/A sky130_fd_sc_hd__buf_6
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout155 _17384_/A2 vssd1 vssd1 vccd1 vccd1 _17396_/A2 sky130_fd_sc_hd__buf_4
Xfanout166 _17296_/Y vssd1 vssd1 vccd1 vccd1 _17354_/A2 sky130_fd_sc_hd__buf_2
Xfanout177 _15552_/X vssd1 vssd1 vccd1 vccd1 _16827_/B sky130_fd_sc_hd__buf_4
Xfanout188 _15752_/A vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__buf_6
Xfanout199 _14926_/X vssd1 vssd1 vccd1 vccd1 _17164_/C sky130_fd_sc_hd__buf_6
XFILLER_170_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09728_ _12107_/A _11900_/B _10036_/D _10645_/C vssd1 vssd1 vccd1 vccd1 _09731_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09659_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__nor2_4
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__xor2_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11621_ _11620_/A _11620_/C _11624_/A vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__o21a_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14340_ _14340_/A _14340_/B _14340_/C vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__nand3_4
X_11552_ _11526_/A _11525_/C _11525_/B vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__a21o_1
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10503_ _10503_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10503_/Y sky130_fd_sc_hd__nand3_2
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14271_ _14350_/A _14271_/B vssd1 vssd1 vccd1 vccd1 _14273_/C sky130_fd_sc_hd__or2_1
X_11483_ _11484_/B _11522_/A _11484_/A vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__o21ai_2
XFILLER_184_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16010_ _15034_/Y _15037_/X _15039_/X _15057_/X _15035_/S _15458_/A vssd1 vssd1 vccd1
+ vccd1 _16010_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10434_ _10434_/A _10547_/A vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__nor2_4
X_13222_ _16649_/A _13223_/B vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__or2_2
XFILLER_136_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13153_ _13154_/B _13154_/A vssd1 vssd1 vccd1 vccd1 _13295_/A sky130_fd_sc_hd__nand2b_2
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _10236_/X _10365_/B vssd1 vssd1 vccd1 vccd1 _10370_/C sky130_fd_sc_hd__and2b_4
XFILLER_151_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12104_/A _12270_/C vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13084_ _13084_/A _13213_/B vssd1 vssd1 vccd1 vccd1 _13085_/C sky130_fd_sc_hd__nor2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10296_/A _10301_/A _10296_/C vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__or3_4
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_33_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16912_ _16913_/C _17134_/C _14865_/B vssd1 vssd1 vccd1 vccd1 _16914_/A sky130_fd_sc_hd__a21boi_2
X_12035_ _16011_/B _12390_/S _12035_/C vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__or3_2
XFILLER_111_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16843_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16844_/B sky130_fd_sc_hd__or2_1
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_1018 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16774_ _16774_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16775_/B sky130_fd_sc_hd__xnor2_2
X_13986_ _13986_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13988_/B sky130_fd_sc_hd__nor2_2
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ _16136_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _15820_/C sky130_fd_sc_hd__nand2_2
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _12985_/A vssd1 vssd1 vccd1 vccd1 _13125_/A sky130_fd_sc_hd__inv_2
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15656_ _15656_/A _15656_/B vssd1 vssd1 vccd1 vccd1 _15679_/A sky130_fd_sc_hd__xnor2_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ _17399_/A _13566_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__a21oi_2
XFILLER_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14558_/B _14560_/B _14558_/A vssd1 vssd1 vccd1 vccd1 _14609_/B sky130_fd_sc_hd__o21ba_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11819_ _17367_/A _12546_/B _12546_/C _11818_/Y vssd1 vssd1 vccd1 vccd1 _11820_/A
+ sky130_fd_sc_hd__a31o_4
X_15587_ _15685_/B _15587_/B vssd1 vssd1 vccd1 vccd1 _15588_/B sky130_fd_sc_hd__xnor2_4
XFILLER_61_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _12799_/A _12799_/B vssd1 vssd1 vccd1 vccd1 _12801_/A sky130_fd_sc_hd__nor2_4
XFILLER_105_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17326_ _13551_/D _17328_/A2 _17325_/X _17402_/C1 vssd1 vssd1 vccd1 vccd1 _17492_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14538_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14538_/X sky130_fd_sc_hd__or2_1
XFILLER_105_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17257_ _17453_/Q _17293_/A2 _17255_/X _17256_/X _17358_/C1 vssd1 vssd1 vccd1 vccd1
+ _17453_/D sky130_fd_sc_hd__o221a_1
X_14469_ _14469_/A _14469_/B vssd1 vssd1 vccd1 vccd1 _14471_/B sky130_fd_sc_hd__xnor2_1
XFILLER_190_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16208_ _16209_/C _16209_/B _14859_/B vssd1 vssd1 vccd1 vccd1 _16300_/A sky130_fd_sc_hd__a21boi_4
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ input15/X input20/X input22/X input21/X vssd1 vssd1 vccd1 vccd1 _17191_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_190_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16139_ _16140_/A _16140_/B vssd1 vssd1 vccd1 vccd1 _16250_/B sky130_fd_sc_hd__and2b_1
XFILLER_143_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ _08962_/B _08962_/C _08962_/A vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__a21oi_2
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08892_ _16315_/A _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__o21ba_4
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09513_ _09513_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__nor2_1
XFILLER_65_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09584_/A _12595_/B _12795_/B _11859_/C vssd1 vssd1 vccd1 vccd1 _09447_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_52_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _09375_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10150_ _10970_/A _10755_/D _10039_/A _10037_/Y vssd1 vssd1 vccd1 vccd1 _10151_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _10081_/A _10081_/B vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__and2_1
XFILLER_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13840_ _12862_/X _12866_/B _17369_/A vssd1 vssd1 vccd1 vccd1 _14839_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwb_buttons_leds_952 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_952/HI led_enb[5] sky130_fd_sc_hd__conb_1
XFILLER_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13771_ _13921_/A _13771_/B vssd1 vssd1 vccd1 vccd1 _13812_/A sky130_fd_sc_hd__nand2_2
X_10983_ _10984_/A _10984_/C vssd1 vssd1 vccd1 vccd1 _10985_/B sky130_fd_sc_hd__nor2_2
XFILLER_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15510_ _15510_/A _15510_/B vssd1 vssd1 vccd1 vccd1 _15512_/B sky130_fd_sc_hd__xor2_4
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12722_ _17397_/A _17395_/A _14215_/B _13566_/B vssd1 vssd1 vccd1 vccd1 _12723_/B
+ sky130_fd_sc_hd__and4_1
X_16490_ _12560_/A _17163_/A2 _16489_/X vssd1 vssd1 vccd1 vccd1 _16492_/B sky130_fd_sc_hd__o21ba_1
XFILLER_130_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15441_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__and2b_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12653_ _12654_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _12655_/A sky130_fd_sc_hd__or2_4
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11603_/A _11603_/C _11603_/B vssd1 vssd1 vccd1 vccd1 _11605_/D sky130_fd_sc_hd__o21ai_1
XFILLER_129_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15372_ _17377_/A _15796_/B _14896_/B vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__o21a_1
X_12584_ _12585_/A _12585_/B _12585_/C vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__a21oi_1
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17111_ _14596_/Y _17163_/A2 _17110_/X _16977_/A vssd1 vssd1 vccd1 vccd1 _17113_/B
+ sky130_fd_sc_hd__o211a_1
X_14323_ _14242_/A _14244_/B _14242_/B vssd1 vssd1 vccd1 vccd1 _14325_/B sky130_fd_sc_hd__o21ba_1
X_11535_ _11541_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11537_/B sky130_fd_sc_hd__nand2_2
XFILLER_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17042_ _17119_/A _17043_/B _17043_/C vssd1 vssd1 vccd1 vccd1 _17044_/A sky130_fd_sc_hd__a21oi_1
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14254_ _14254_/A _14554_/B vssd1 vssd1 vccd1 vccd1 _14255_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ _11444_/A _11444_/C _11444_/B vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__a21o_1
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap119 _12631_/A vssd1 vssd1 vccd1 vccd1 _12784_/B1 sky130_fd_sc_hd__clkbuf_2
X_13205_ _13201_/Y _13203_/A _13075_/A _13075_/Y vssd1 vssd1 vccd1 vccd1 _13249_/B
+ sky130_fd_sc_hd__o211ai_4
X_10417_ _10418_/A _10418_/C vssd1 vssd1 vccd1 vccd1 _10423_/B sky130_fd_sc_hd__nor2_2
X_14185_ _14185_/A _14185_/B vssd1 vssd1 vccd1 vccd1 _14186_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11397_ _11384_/Y _11396_/X _11403_/A _11368_/Y vssd1 vssd1 vccd1 vccd1 _11403_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_140_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _13136_/A vssd1 vssd1 vccd1 vccd1 _13137_/B sky130_fd_sc_hd__inv_2
XFILLER_98_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10348_ _10348_/A _10348_/B _10348_/C vssd1 vssd1 vccd1 vccd1 _11775_/B sky130_fd_sc_hd__or3_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _10387_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__and2_2
XFILLER_97_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13067_ _17425_/A _17423_/A _13067_/C _13067_/D vssd1 vssd1 vccd1 vccd1 _13068_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_94_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _12374_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12018_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _16683_/A _16758_/B _16695_/B _16604_/B vssd1 vssd1 vccd1 vccd1 _16828_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ _16758_/A _16758_/B _16758_/C vssd1 vssd1 vccd1 vccd1 _16759_/A sky130_fd_sc_hd__a21oi_1
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13969_ _13969_/A _13969_/B vssd1 vssd1 vccd1 vccd1 _13971_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15708_ _15707_/A _15707_/B _15707_/C vssd1 vssd1 vccd1 vccd1 _15708_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16688_ _16688_/A _16688_/B vssd1 vssd1 vccd1 vccd1 _16690_/B sky130_fd_sc_hd__xor2_2
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15639_ _17038_/C _15639_/B vssd1 vssd1 vccd1 vccd1 _16499_/B sky130_fd_sc_hd__or2_4
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _09926_/A _12597_/B _14948_/B vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__and3_2
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17309_ input64/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17309_/X sky130_fd_sc_hd__or3_1
X_09091_ _09091_/A _09091_/B _09318_/A vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__and3_2
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_960 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09986_/A _09988_/B _09986_/B vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__o21ba_4
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08944_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08875_ _08832_/A _08832_/C _08832_/B vssd1 vssd1 vccd1 vccd1 _08875_/X sky130_fd_sc_hd__o21a_2
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09427_ _17119_/B _16933_/A vssd1 vssd1 vccd1 vccd1 _09427_/Y sky130_fd_sc_hd__nor2_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ _09358_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _09366_/C sky130_fd_sc_hd__or2_1
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__xnor2_2
XFILLER_166_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11320_ _11320_/A _11320_/B _11320_/C vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__or3_4
XFILLER_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11251_ _11347_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11348_/A sky130_fd_sc_hd__or2_4
XFILLER_162_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10202_ _10202_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10203_/C sky130_fd_sc_hd__xnor2_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11182_ _11182_/A _11182_/B _11182_/C vssd1 vssd1 vccd1 vccd1 _11182_/Y sky130_fd_sc_hd__nor3_4
XFILLER_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ _10133_/A _10133_/B _10133_/C vssd1 vssd1 vccd1 vccd1 _10134_/C sky130_fd_sc_hd__nand3_4
X_15990_ _16096_/B _15990_/B vssd1 vssd1 vccd1 vccd1 _15990_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_76_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10064_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14941_ _11841_/A _15373_/B _10560_/D vssd1 vssd1 vccd1 vccd1 _14941_/X sky130_fd_sc_hd__a21o_1
XFILLER_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14872_ _14872_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _16977_/A sky130_fd_sc_hd__or2_4
X_16611_ _16612_/B _16611_/B vssd1 vssd1 vccd1 vccd1 _16697_/B sky130_fd_sc_hd__and2b_1
X_13823_ _13823_/A _13823_/B vssd1 vssd1 vccd1 vccd1 _13827_/A sky130_fd_sc_hd__xor2_4
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17591_ fanout938/X _17591_/D vssd1 vssd1 vccd1 vccd1 _17591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16542_ _16542_/A _16542_/B vssd1 vssd1 vccd1 vccd1 _16543_/B sky130_fd_sc_hd__nor2_2
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13754_ _13754_/A _13754_/B vssd1 vssd1 vccd1 vccd1 _13756_/B sky130_fd_sc_hd__xnor2_1
XFILLER_188_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10966_ _10966_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__xnor2_4
X_12705_ _12044_/Y _12046_/Y _12049_/Y _12051_/Y _15038_/A _15312_/S vssd1 vssd1 vccd1
+ vccd1 _12705_/X sky130_fd_sc_hd__mux4_2
X_16473_ _16563_/A _16384_/Y _16472_/X vssd1 vssd1 vccd1 vccd1 _16475_/A sky130_fd_sc_hd__a21oi_1
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13685_ _13686_/A _13686_/B vssd1 vssd1 vccd1 vccd1 _13787_/A sky130_fd_sc_hd__or2_2
X_10897_ _14922_/S _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__and3_1
XFILLER_176_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15424_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15426_/B sky130_fd_sc_hd__xor2_4
X_12636_ _14770_/A _12637_/C _12637_/D _14769_/A vssd1 vssd1 vccd1 vccd1 _12640_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_54_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15355_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _15356_/B sky130_fd_sc_hd__or2_2
XFILLER_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12567_ _17393_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__nand2_4
XFILLER_157_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14306_ _14306_/A _14306_/B vssd1 vssd1 vccd1 vccd1 _14309_/A sky130_fd_sc_hd__xnor2_2
XFILLER_129_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ _11629_/A _11561_/B _11518_/C _11563_/D vssd1 vssd1 vccd1 vccd1 _11521_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_171_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15286_ _15287_/A _15287_/B vssd1 vssd1 vccd1 vccd1 _15286_/Y sky130_fd_sc_hd__nor2_1
X_12498_ _12498_/A _12498_/B _12498_/C vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__and3_1
XFILLER_176_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ _16972_/A _16972_/B _10583_/A vssd1 vssd1 vccd1 vccd1 _17025_/Y sky130_fd_sc_hd__a21boi_1
X_14237_ _14237_/A _14237_/B _14236_/X vssd1 vssd1 vccd1 vccd1 _14239_/A sky130_fd_sc_hd__nor3b_4
X_11449_ _11453_/B _11449_/B _11449_/C vssd1 vssd1 vccd1 vccd1 _11495_/A sky130_fd_sc_hd__and3_4
XFILLER_125_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14168_ _14168_/A _14641_/D vssd1 vssd1 vccd1 vccd1 _14170_/C sky130_fd_sc_hd__nand2_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13120_/B _13120_/A vssd1 vssd1 vccd1 vccd1 _13119_/Y sky130_fd_sc_hd__nand2b_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _14188_/B _14101_/B vssd1 vssd1 vccd1 vccd1 _14194_/A sky130_fd_sc_hd__nand2_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16809_ _16809_/A _16809_/B _16809_/C vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__and3_1
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09212_ _09212_/A _09212_/B vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__nor2_1
XFILLER_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09143_ _09143_/A _09231_/A vssd1 vssd1 vccd1 vccd1 _09145_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09074_ _09074_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _09076_/C sky130_fd_sc_hd__nand2_2
XFILLER_148_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__xnor2_4
XFILLER_162_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08927_ _08927_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__nand2_4
XFILLER_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ _12275_/A _12107_/B _12090_/B _12088_/C vssd1 vssd1 vccd1 vccd1 _08859_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _12088_/B _11881_/D _11870_/B _12088_/A vssd1 vssd1 vccd1 vccd1 _08792_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _11240_/A _11097_/D _11423_/C _11095_/A vssd1 vssd1 vccd1 vccd1 _10820_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10751_ _10993_/C _10659_/D _10660_/A _10658_/Y vssd1 vssd1 vccd1 vccd1 _10757_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_186_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _17415_/A _13866_/C vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__nand2_2
XFILLER_186_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10682_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10682_/Y sky130_fd_sc_hd__nor2_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12421_ _12421_/A _12421_/B _12421_/C vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__nand3_2
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15140_ _15270_/A _15141_/B vssd1 vssd1 vccd1 vccd1 _15140_/Y sky130_fd_sc_hd__nor2_2
XFILLER_127_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _12351_/A _12351_/B _12350_/X vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__o21bai_1
XFILLER_153_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11303_ _11260_/C _11563_/D _11261_/A _11259_/Y vssd1 vssd1 vccd1 vccd1 _11304_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_15071_ _15071_/A _15071_/B vssd1 vssd1 vccd1 vccd1 _15071_/Y sky130_fd_sc_hd__nor2_2
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12283_ _12283_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__nor2_1
X_14022_ _14113_/B _14022_/B vssd1 vssd1 vccd1 vccd1 _14025_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11234_ _11234_/A _11234_/B vssd1 vssd1 vccd1 vccd1 _11711_/A sky130_fd_sc_hd__or2_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _11165_/A _11165_/B _11165_/C vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__or3_1
XFILLER_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__nor2_2
XFILLER_49_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15973_ _16080_/B _15973_/B vssd1 vssd1 vccd1 vccd1 _15976_/A sky130_fd_sc_hd__nor2_4
X_11096_ _11240_/A _11423_/C _11605_/B _11095_/A vssd1 vssd1 vccd1 vccd1 _11096_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_110_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10047_ _10162_/A _10170_/A _10162_/C vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__o21ai_4
X_14924_ _14924_/A _14929_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _14926_/B sky130_fd_sc_hd__or3_4
XFILLER_36_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14855_ _15811_/A _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15898_/B sky130_fd_sc_hd__and3_1
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13806_ _13915_/B _13806_/B vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__or2_2
X_17574_ fanout938/X _17574_/D vssd1 vssd1 vccd1 vccd1 _17574_/Q sky130_fd_sc_hd__dfxtp_1
X_14786_ _14786_/A _15463_/A vssd1 vssd1 vccd1 vccd1 _14805_/B sky130_fd_sc_hd__or2_1
X_11998_ _11998_/A _11998_/B _12197_/B _11998_/D vssd1 vssd1 vccd1 vccd1 _11998_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16525_ _16616_/B _16525_/B vssd1 vssd1 vccd1 vccd1 _16527_/C sky130_fd_sc_hd__nor2_2
X_13737_ _14775_/A _13844_/D vssd1 vssd1 vccd1 vccd1 _13739_/B sky130_fd_sc_hd__nand2_1
X_10949_ _10946_/X _10947_/Y _10927_/X _11059_/A vssd1 vssd1 vccd1 vccd1 _10949_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16456_ _16457_/B _16457_/A vssd1 vssd1 vccd1 vccd1 _16456_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_177_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13668_ _13668_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13669_/B sky130_fd_sc_hd__and2_1
XFILLER_188_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15407_ _15408_/A _15408_/B _15408_/C vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__o21a_2
X_12619_ _12619_/A _12619_/B vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__nor2_2
X_16387_ _16387_/A _16387_/B _16387_/C vssd1 vssd1 vccd1 vccd1 _16389_/B sky130_fd_sc_hd__or3_2
X_13599_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__nor2_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15338_ _16935_/A _15147_/A _15393_/B vssd1 vssd1 vccd1 vccd1 _15338_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15269_ _15204_/A _16880_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _15270_/C sky130_fd_sc_hd__o21a_1
X_17008_ _17008_/A _17012_/B vssd1 vssd1 vccd1 vccd1 _17009_/B sky130_fd_sc_hd__or2_2
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09830_ _09769_/B _09776_/B _09769_/D _09769_/A vssd1 vssd1 vccd1 vccd1 _09830_/X
+ sky130_fd_sc_hd__a22o_2
Xfanout507 _17517_/Q vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__buf_6
XFILLER_141_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout518 _10640_/C vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__buf_6
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout529 _08718_/A vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__buf_6
XFILLER_141_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09761_ _09761_/A vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__inv_2
XFILLER_101_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09692_ _10236_/A _10235_/A _10490_/C _10479_/B vssd1 vssd1 vccd1 vccd1 _09695_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_187_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ _09128_/D vssd1 vssd1 vccd1 vccd1 _09126_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__nor2_1
XFILLER_151_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_952 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _09960_/A _09960_/B _09960_/C vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__and3_2
XTAP_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12970_ _12971_/B _12971_/A vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__and2b_1
XTAP_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _11921_/A _12179_/A vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__or2_1
XTAP_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14738_/A _14867_/A vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__nand2_4
XFILLER_61_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11852_ _15095_/B _11852_/B vssd1 vssd1 vccd1 vccd1 _11854_/C sky130_fd_sc_hd__or2_2
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10803_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10816_/A sky130_fd_sc_hd__xnor2_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14621_/A _14570_/C _14570_/A vssd1 vssd1 vccd1 vccd1 _14571_/X sky130_fd_sc_hd__a21o_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _14872_/A _14924_/C vssd1 vssd1 vccd1 vccd1 _15011_/B sky130_fd_sc_hd__nor2_4
X_16310_ _16310_/A _16310_/B _16310_/C _16310_/D vssd1 vssd1 vccd1 vccd1 _16310_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_186_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13522_ _13844_/A _13844_/B _14002_/B _13897_/B vssd1 vssd1 vccd1 vccd1 _13637_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_159_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17290_ _17464_/Q _17290_/A2 _17288_/X _17289_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17464_/D sky130_fd_sc_hd__o221a_1
X_10734_ _10662_/X _10732_/Y _10728_/B _10714_/X vssd1 vssd1 vccd1 vccd1 _10734_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_159_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16241_ _16241_/A _16241_/B _16239_/Y vssd1 vssd1 vccd1 vccd1 _16242_/B sky130_fd_sc_hd__or3b_4
X_13453_ _14387_/A _13564_/C _13453_/C vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__and3_1
XFILLER_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10665_ _10670_/B _10665_/B vssd1 vssd1 vccd1 vccd1 _10667_/B sky130_fd_sc_hd__nand2_2
XFILLER_167_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12404_ _14776_/A _13450_/D _13866_/D _17403_/A vssd1 vssd1 vccd1 vccd1 _12406_/A
+ sky130_fd_sc_hd__a22oi_1
X_16172_ _16172_/A _16172_/B vssd1 vssd1 vccd1 vccd1 _16174_/A sky130_fd_sc_hd__xor2_4
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13384_ _13261_/A _13263_/A _13504_/B _13382_/X vssd1 vssd1 vccd1 vccd1 _13385_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ _10709_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__or2_4
XFILLER_12_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15123_ _15126_/B vssd1 vssd1 vccd1 vccd1 _15123_/Y sky130_fd_sc_hd__inv_2
X_12335_ _12500_/A _12638_/B _12334_/C vssd1 vssd1 vccd1 vccd1 _12336_/B sky130_fd_sc_hd__a21oi_2
XFILLER_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ _16207_/B _15053_/X _15051_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _15054_/X
+ sky130_fd_sc_hd__o211a_1
X_12266_ _12266_/A _12437_/B vssd1 vssd1 vccd1 vccd1 _12268_/C sky130_fd_sc_hd__nand2_2
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14005_ _13904_/A _13904_/B _13902_/B vssd1 vssd1 vccd1 vccd1 _14007_/B sky130_fd_sc_hd__o21ai_4
X_11217_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__xnor2_4
X_12197_ _12197_/A _12197_/B vssd1 vssd1 vccd1 vccd1 _12198_/C sky130_fd_sc_hd__nor2_2
Xoutput81 _17474_/Q vssd1 vssd1 vccd1 vccd1 leds[8] sky130_fd_sc_hd__clkbuf_2
Xoutput92 _17451_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[17] sky130_fd_sc_hd__clkbuf_2
X_11148_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11149_/B sky130_fd_sc_hd__nand2_1
XFILLER_163_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15956_ _16446_/A _15956_/B vssd1 vssd1 vccd1 vccd1 _16062_/C sky130_fd_sc_hd__nor2_1
X_11079_ _11077_/A _11077_/C _11110_/A vssd1 vssd1 vccd1 vccd1 _11080_/D sky130_fd_sc_hd__o21ai_4
XFILLER_110_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14907_ _14899_/C _14906_/X _14905_/X _14903_/X vssd1 vssd1 vccd1 vccd1 _15553_/B
+ sky130_fd_sc_hd__o211a_4
X_15887_ _15884_/Y _15885_/Y _15886_/Y vssd1 vssd1 vccd1 vccd1 _15887_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14838_ _12016_/B _11781_/B _14837_/Y vssd1 vssd1 vccd1 vccd1 _14838_/X sky130_fd_sc_hd__o21a_2
XTAP_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17557_ fanout939/X _17557_/D vssd1 vssd1 vccd1 vccd1 _17557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14769_ _14769_/A _14769_/B vssd1 vssd1 vccd1 vccd1 _16918_/B sky130_fd_sc_hd__or2_2
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16508_ _16509_/A _16509_/B _16509_/C vssd1 vssd1 vccd1 vccd1 _16616_/A sky130_fd_sc_hd__a21oi_4
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17488_ fanout931/X _17488_/D vssd1 vssd1 vccd1 vccd1 _17488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16439_ _16439_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__xor2_2
XFILLER_20_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout304 _08719_/Y vssd1 vssd1 vccd1 vccd1 _15175_/A sky130_fd_sc_hd__buf_8
XFILLER_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout315 _14832_/A vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__buf_6
Xfanout326 _17134_/A vssd1 vssd1 vccd1 vccd1 _14213_/B sky130_fd_sc_hd__buf_4
XFILLER_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09813_/A _09813_/B _09813_/C vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__and3_2
Xfanout337 _17538_/Q vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__buf_8
Xfanout348 _13977_/B vssd1 vssd1 vccd1 vccd1 _14153_/B sky130_fd_sc_hd__buf_6
Xfanout359 _17535_/Q vssd1 vssd1 vccd1 vccd1 _12487_/A sky130_fd_sc_hd__buf_12
X_09744_ _09724_/X _09740_/B _09743_/Y _09621_/X vssd1 vssd1 vccd1 vccd1 _09776_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_74_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09675_ _09678_/B _09675_/B _09675_/C vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__nor3_2
XFILLER_54_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _10450_/A _10450_/B vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09109_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__and2_1
XFILLER_184_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10381_ _10382_/B _10382_/A vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__nand2b_2
XFILLER_191_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12120_ _12309_/A _12118_/Y _11905_/X _11909_/A vssd1 vssd1 vccd1 vccd1 _12122_/D
+ sky130_fd_sc_hd__a211o_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _14911_/B _12051_/B vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__nand2_1
XFILLER_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_974 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11002_ _10999_/X _11000_/Y _10977_/X _11051_/A vssd1 vssd1 vccd1 vccd1 _11002_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout860 _10805_/C vssd1 vssd1 vccd1 vccd1 _11005_/B sky130_fd_sc_hd__buf_8
Xfanout871 _10805_/D vssd1 vssd1 vccd1 vccd1 _10360_/D sky130_fd_sc_hd__buf_6
X_15810_ _14924_/A _12401_/A _13390_/X _15804_/Y _15809_/Y vssd1 vssd1 vccd1 vccd1
+ _15810_/X sky130_fd_sc_hd__o311a_1
X_16790_ _14168_/A _16789_/Y _16788_/Y vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__a21oi_2
Xfanout882 _10809_/D vssd1 vssd1 vccd1 vccd1 _11097_/D sky130_fd_sc_hd__buf_6
XFILLER_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout893 _11370_/C vssd1 vssd1 vccd1 vccd1 _15008_/A sky130_fd_sc_hd__buf_2
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15741_ _15741_/A _15741_/B vssd1 vssd1 vccd1 vccd1 _15743_/B sky130_fd_sc_hd__xnor2_2
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ _12795_/A _12795_/B _12796_/A _12794_/B vssd1 vssd1 vccd1 vccd1 _12954_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11904_ _08859_/A _08861_/B _08859_/B vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__o21ba_1
X_15672_ _15673_/A _15673_/B vssd1 vssd1 vccd1 vccd1 _15764_/B sky130_fd_sc_hd__nand2_2
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12884_/A _12884_/B vssd1 vssd1 vccd1 vccd1 _12886_/C sky130_fd_sc_hd__xnor2_4
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14624_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14660_/B sky130_fd_sc_hd__nor2_2
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17411_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17411_/X sky130_fd_sc_hd__or2_1
X_11835_ _12031_/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11835_/Y sky130_fd_sc_hd__nand2_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _12565_/C _17360_/A2 _17341_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17500_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14554_ _16965_/C _14554_/B vssd1 vssd1 vccd1 vccd1 _14555_/B sky130_fd_sc_hd__nand2_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _16866_/A _16866_/B vssd1 vssd1 vccd1 vccd1 _11766_/X sky130_fd_sc_hd__or2_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13505_ _13506_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__nand2_1
XFILLER_187_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17273_ _17600_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__a21o_1
X_10717_ _10963_/A _10963_/B _10962_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _10720_/A
+ sky130_fd_sc_hd__and4_2
X_14485_ _14593_/A _14593_/B _14545_/D _14485_/D vssd1 vssd1 vccd1 vccd1 _14557_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11697_ _15614_/A _15614_/B vssd1 vssd1 vccd1 vccd1 _15615_/A sky130_fd_sc_hd__nor2_1
X_16224_ _16224_/A vssd1 vssd1 vccd1 vccd1 _17559_/D sky130_fd_sc_hd__inv_2
X_13436_ _17421_/A _13664_/D vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__nand2_1
X_10648_ _10648_/A _10742_/A vssd1 vssd1 vccd1 vccd1 _10735_/A sky130_fd_sc_hd__or2_2
XFILLER_127_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16155_ _16155_/A _16155_/B vssd1 vssd1 vccd1 vccd1 _16157_/B sky130_fd_sc_hd__xnor2_4
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13367_ _13368_/A _13368_/B vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__nand2_4
XFILLER_115_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10579_ _10579_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _10582_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15106_ _15106_/A _15106_/B vssd1 vssd1 vccd1 vccd1 _15106_/Y sky130_fd_sc_hd__nand2_1
XFILLER_114_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12318_ _12150_/A _12149_/B _12149_/A vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__o21ba_4
X_16086_ _16281_/A _16355_/B _16086_/C vssd1 vssd1 vccd1 vccd1 _16197_/B sky130_fd_sc_hd__and3_1
XFILLER_181_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _13298_/A _13745_/D vssd1 vssd1 vccd1 vccd1 _13657_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _15097_/A _15037_/B vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__or2_2
X_12249_ _12250_/A _12250_/B vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__nand2b_2
XFILLER_123_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16988_ _16989_/A _16989_/B vssd1 vssd1 vccd1 vccd1 _17049_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _15939_/A _15939_/B vssd1 vssd1 vccd1 vccd1 _15940_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09460_ _09440_/X _09455_/B _09459_/Y _09335_/A vssd1 vssd1 vccd1 vccd1 _09460_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17609_ fanout925/X _17609_/D vssd1 vssd1 vccd1 vccd1 _17609_/Q sky130_fd_sc_hd__dfxtp_4
X_09391_ _09391_/A _09391_/B _09391_/C vssd1 vssd1 vccd1 vccd1 _09393_/D sky130_fd_sc_hd__and3_4
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout123 _17229_/B vssd1 vssd1 vccd1 vccd1 _17232_/B sky130_fd_sc_hd__buf_4
Xfanout134 _15755_/B vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout145 _16165_/A vssd1 vssd1 vccd1 vccd1 _15662_/A sky130_fd_sc_hd__buf_6
Xfanout156 _17384_/A2 vssd1 vssd1 vccd1 vccd1 _17422_/A2 sky130_fd_sc_hd__buf_4
Xfanout167 _16409_/B vssd1 vssd1 vccd1 vccd1 _16938_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout178 _15552_/X vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__buf_4
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ _09727_/A _09727_/B vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__nor2_1
XFILLER_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09658_ _09658_/A _09658_/B vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__or2_2
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A _09589_/B vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__xnor2_1
XFILLER_163_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11620_/A _11624_/A _11620_/C vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__nor3_1
XFILLER_179_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11551_ _11538_/A _11537_/C _11537_/B vssd1 vssd1 vccd1 vccd1 _11551_/X sky130_fd_sc_hd__o21a_2
XFILLER_184_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10502_ _10503_/A _10503_/B _10503_/C vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__a21o_4
X_14270_ _14270_/A _14270_/B _14270_/C vssd1 vssd1 vccd1 vccd1 _14271_/B sky130_fd_sc_hd__and3_1
X_11482_ _11484_/B _11481_/Y _11520_/C _11518_/C vssd1 vssd1 vccd1 vccd1 _11522_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_183_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13221_ _13221_/A _13221_/B vssd1 vssd1 vccd1 vccd1 _13223_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10433_ _10434_/A _10432_/Y _10993_/C _10543_/B vssd1 vssd1 vccd1 vccd1 _10547_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ _13019_/A _13021_/B _13019_/B vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__o21ba_1
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__xor2_4
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ _12103_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__nor2_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _13083_/A _13213_/A _13083_/C vssd1 vssd1 vccd1 vccd1 _13213_/B sky130_fd_sc_hd__nor3_2
X_10295_ _10296_/A _10296_/C vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nor2_2
X_16911_ _16911_/A _16911_/B vssd1 vssd1 vccd1 vccd1 _16911_/Y sky130_fd_sc_hd__nand2_2
X_12034_ _12031_/Y _12033_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__mux2_2
XFILLER_105_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16842_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16906_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout690 _12021_/B vssd1 vssd1 vccd1 vccd1 _14863_/B sky130_fd_sc_hd__buf_6
XFILLER_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16773_ _16774_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__and2b_1
X_13985_ _13985_/A _13985_/B vssd1 vssd1 vccd1 vccd1 _13988_/A sky130_fd_sc_hd__xor2_4
XFILLER_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15724_ _16136_/A _16020_/B vssd1 vssd1 vccd1 vccd1 _15726_/D sky130_fd_sc_hd__and2_4
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12936_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__a21oi_4
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15655_ _15655_/A _15655_/B _15656_/B vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__and3_1
XFILLER_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _14421_/S _12864_/Y _12866_/Y _13516_/S _08718_/A vssd1 vssd1 vccd1 vccd1
+ _12867_/X sky130_fd_sc_hd__a221o_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14606_ _14606_/A _14606_/B vssd1 vssd1 vccd1 vccd1 _14609_/A sky130_fd_sc_hd__xor2_2
XFILLER_159_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11818_ _17367_/A _11818_/B vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__nor2_1
X_15586_ _15685_/B _15587_/B vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__and2b_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _12798_/A _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12799_/B sky130_fd_sc_hd__and3_1
XFILLER_187_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _13939_/A _14281_/Y _14534_/Y _14535_/Y _14536_/X vssd1 vssd1 vccd1 vccd1
+ _14629_/B sky130_fd_sc_hd__o311ai_4
X_17325_ input41/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17325_/X sky130_fd_sc_hd__or3_1
X_11749_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__xnor2_4
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468_ _14469_/A _14469_/B vssd1 vssd1 vccd1 vccd1 _14531_/A sky130_fd_sc_hd__nor2_1
X_17256_ _17562_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__and2_1
XFILLER_146_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13419_ _13420_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13419_/Y sky130_fd_sc_hd__nand2b_2
X_16207_ _16294_/B _16207_/B _16207_/C vssd1 vssd1 vccd1 vccd1 _16207_/X sky130_fd_sc_hd__or3_4
X_17187_ input28/X _17362_/B _17429_/B vssd1 vssd1 vccd1 vccd1 _17187_/Y sky130_fd_sc_hd__nor3_1
X_14399_ _14466_/A _14400_/C _14400_/A vssd1 vssd1 vccd1 vccd1 _14399_/X sky130_fd_sc_hd__a21o_1
XFILLER_127_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16138_ _16410_/A _16499_/B vssd1 vssd1 vccd1 vccd1 _16140_/B sky130_fd_sc_hd__nor2_2
XFILLER_115_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16069_ _16070_/A _16070_/B vssd1 vssd1 vccd1 vccd1 _16069_/Y sky130_fd_sc_hd__nand2b_1
X_08960_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _08962_/C sky130_fd_sc_hd__nand2_1
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08891_ _08904_/B _08904_/C _08904_/A vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__a21o_4
XFILLER_97_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1007 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09512_ _10062_/A _09937_/B _09379_/A _09377_/Y vssd1 vssd1 vccd1 vccd1 _09513_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09443_ _09443_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__nor2_1
XFILLER_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09374_ _10062_/A _09791_/B _09206_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _09375_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_178_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10080_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__or2_1
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwb_buttons_leds_953 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_953/HI led_enb[6] sky130_fd_sc_hd__conb_1
X_13770_ _13770_/A _13770_/B _13770_/C vssd1 vssd1 vccd1 vccd1 _13771_/B sky130_fd_sc_hd__or3_1
X_10982_ _10647_/C _10745_/D _10746_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _10984_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12721_ _13405_/B _14215_/B _13566_/B _14777_/A vssd1 vssd1 vccd1 vccd1 _12723_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_167_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _15363_/A _15363_/B _15361_/Y vssd1 vssd1 vccd1 vccd1 _15442_/B sky130_fd_sc_hd__a21bo_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ _12800_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _11603_/A _11603_/B _11603_/C vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__or3_2
X_15371_ _15303_/A _15370_/X _15794_/A _11691_/Y vssd1 vssd1 vccd1 vccd1 _15390_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12583_ _12583_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12585_/C sky130_fd_sc_hd__xnor2_2
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _14324_/A _14389_/B vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__nor2_1
XFILLER_90_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17110_ _14867_/A _16974_/B _14929_/X _14827_/Y vssd1 vssd1 vccd1 vccd1 _17110_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11534_ _11534_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11535_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17041_ _16982_/A _17119_/B _17039_/X _17085_/A vssd1 vssd1 vccd1 vccd1 _17043_/C
+ sky130_fd_sc_hd__a211oi_2
X_14253_ _14253_/A _14253_/B vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__nor2_4
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _11465_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _15997_/A sky130_fd_sc_hd__xor2_4
XFILLER_165_980 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13204_ _13075_/A _13075_/Y _13201_/Y _13203_/A vssd1 vssd1 vccd1 vccd1 _13249_/A
+ sky130_fd_sc_hd__a211o_4
X_10416_ _10299_/C _10659_/D _10300_/A _10298_/Y vssd1 vssd1 vccd1 vccd1 _10418_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14184_ _14185_/A _14273_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _14186_/A sky130_fd_sc_hd__and3_1
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11396_ _11396_/A _11396_/B _11396_/C vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__and3_4
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13135_ _13264_/B _13132_/X _12993_/X _12999_/A vssd1 vssd1 vccd1 vccd1 _13136_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10347_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__or2_1
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _17423_/A _13067_/C _13067_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _13068_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_140_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10278_ _10278_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10387_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _11780_/Y _12377_/A _12015_/Y vssd1 vssd1 vccd1 vccd1 _12018_/B sky130_fd_sc_hd__o21ai_2
XFILLER_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16825_ _16938_/A _16935_/B _16746_/A _16744_/B vssd1 vssd1 vccd1 vccd1 _16829_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_48_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16756_ _16827_/A _16827_/C vssd1 vssd1 vccd1 vccd1 _16758_/C sky130_fd_sc_hd__nor2_2
X_13968_ _14215_/A _14141_/D vssd1 vssd1 vccd1 vccd1 _13969_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _15707_/A _15707_/B _15707_/C vssd1 vssd1 vccd1 vccd1 _15707_/Y sky130_fd_sc_hd__nand3_1
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _12919_/A _13065_/B vssd1 vssd1 vccd1 vccd1 _12920_/C sky130_fd_sc_hd__nand2_2
X_16687_ _16685_/X _16687_/B vssd1 vssd1 vccd1 vccd1 _16688_/B sky130_fd_sc_hd__and2b_1
X_13899_ _13790_/A _13792_/B _13790_/B vssd1 vssd1 vccd1 vccd1 _13900_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15638_ _17038_/C _15639_/B vssd1 vssd1 vccd1 vccd1 _15638_/Y sky130_fd_sc_hd__nor2_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15569_ _16262_/A _16410_/A vssd1 vssd1 vccd1 vccd1 _15570_/B sky130_fd_sc_hd__nor2_4
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17308_ _12295_/D _17328_/A2 _17307_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17483_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09090_ _09091_/B _09318_/A _09091_/A vssd1 vssd1 vccd1 vccd1 _09093_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17239_ _17447_/Q _17290_/A2 _17237_/X _17238_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17447_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_972 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09992_ _10004_/B _10004_/C _10004_/A vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__a21o_2
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _08943_/A _08943_/B vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__xnor2_4
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08874_ _08874_/A _08874_/B _08873_/C _08873_/D vssd1 vssd1 vccd1 vccd1 _08874_/X
+ sky130_fd_sc_hd__or4bb_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ _09566_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _17038_/B sky130_fd_sc_hd__nand2_8
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09357_ _09357_/A _09364_/A _09357_/C vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__nor3_1
XFILLER_138_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09288_ _09289_/B _09289_/A vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__nand2b_2
XFILLER_176_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11255_/B _11250_/B vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__nand2_1
XFILLER_180_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10201_ _10202_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10469_/A sky130_fd_sc_hd__and2b_1
XFILLER_192_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11181_ _11181_/A _11181_/B vssd1 vssd1 vccd1 vccd1 _11182_/C sky130_fd_sc_hd__xnor2_4
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_161_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__xnor2_4
XFILLER_95_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _10062_/A _09944_/D _09945_/A _09943_/Y vssd1 vssd1 vccd1 vccd1 _10064_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_88_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14940_ _17607_/Q _17477_/D _17476_/D _17608_/Q vssd1 vssd1 vccd1 vccd1 _16391_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_121_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14871_ _14872_/A _14933_/B vssd1 vssd1 vccd1 vccd1 _14871_/Y sky130_fd_sc_hd__nor2_4
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16610_ _16697_/A _16610_/B vssd1 vssd1 vccd1 vccd1 _16612_/B sky130_fd_sc_hd__or2_1
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13822_ _13823_/A _13823_/B vssd1 vssd1 vccd1 vccd1 _13930_/B sky130_fd_sc_hd__and2b_1
X_17590_ fanout939/X _17590_/D vssd1 vssd1 vccd1 vccd1 _17590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _16541_/A _16541_/B vssd1 vssd1 vccd1 vccd1 _16542_/B sky130_fd_sc_hd__nor2_1
X_13753_ _13754_/B _13754_/A vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__nand2b_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _10965_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__nor2_2
X_12704_ _12020_/Y _12022_/Y _12053_/Y _12055_/Y _12390_/S _15254_/S vssd1 vssd1 vccd1
+ vccd1 _12704_/X sky130_fd_sc_hd__mux4_2
XFILLER_44_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16472_ _16563_/B _16564_/A vssd1 vssd1 vccd1 vccd1 _16472_/X sky130_fd_sc_hd__or2_1
X_13684_ _13587_/B _13589_/B _13587_/A vssd1 vssd1 vccd1 vccd1 _13686_/B sky130_fd_sc_hd__o21ba_1
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10896_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__or2_4
XFILLER_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12635_ _12478_/A _12478_/B _12477_/A vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__a21oi_2
X_15423_ _15424_/A _15424_/B vssd1 vssd1 vccd1 vccd1 _15505_/A sky130_fd_sc_hd__nor2_4
XFILLER_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15354_ _15355_/A _15355_/B vssd1 vssd1 vccd1 vccd1 _15356_/A sky130_fd_sc_hd__nand2_2
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12566_ _12566_/A _12566_/B vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__nor2_2
XFILLER_180_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14305_ _14306_/A _14306_/B vssd1 vssd1 vccd1 vccd1 _14378_/A sky130_fd_sc_hd__nand2b_2
XFILLER_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11517_ _11651_/A _15175_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__nand2_4
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ _15285_/A _15285_/B vssd1 vssd1 vccd1 vccd1 _15287_/B sky130_fd_sc_hd__xnor2_4
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12498_/A _12498_/B _12498_/C vssd1 vssd1 vccd1 vccd1 _12499_/A sky130_fd_sc_hd__a21oi_1
X_14236_ _14315_/A _14236_/B vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__and2_1
XFILLER_172_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17024_ _17024_/A _17024_/B vssd1 vssd1 vccd1 vccd1 _17024_/X sky130_fd_sc_hd__xor2_1
XFILLER_116_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11448_ _11448_/A _11448_/B vssd1 vssd1 vccd1 vccd1 _11449_/C sky130_fd_sc_hd__and2_2
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14167_ _14450_/A _14318_/B _14545_/C _14545_/D vssd1 vssd1 vccd1 vccd1 _14245_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_113_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ _11553_/A _11377_/C _11377_/D _11506_/A vssd1 vssd1 vccd1 vccd1 _11380_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_124_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _13118_/A _13118_/B vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand2_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14098_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14101_/B sky130_fd_sc_hd__nand2_1
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13049_/A _13049_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13061_/B sky130_fd_sc_hd__nand3_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1034 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16808_ _16809_/A _16809_/C _16743_/C _16938_/A vssd1 vssd1 vccd1 vccd1 _16808_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16739_ _16917_/A _16791_/B _16725_/X _16738_/X vssd1 vssd1 vccd1 vccd1 _16739_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ _09211_/A _09211_/B _09373_/A vssd1 vssd1 vccd1 vccd1 _09212_/B sky130_fd_sc_hd__nor3_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09142_ _12174_/A _12174_/B _12127_/C _12127_/D vssd1 vssd1 vccd1 vccd1 _09231_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09073_ _08985_/A _08985_/B _08985_/C vssd1 vssd1 vccd1 vccd1 _09074_/B sky130_fd_sc_hd__o21ai_1
XFILLER_147_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_950 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_162_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09975_ _09865_/A _09864_/C _09864_/B vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08926_ _08917_/X _09053_/A _09012_/A _08910_/Y vssd1 vssd1 vccd1 vccd1 _09012_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08857_ _12107_/B _12090_/B _12088_/C _12275_/A vssd1 vssd1 vccd1 vccd1 _08859_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _12245_/A _11867_/D _08779_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08796_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10750_ _10750_/A _10750_/B _10750_/C vssd1 vssd1 vccd1 vccd1 _10760_/B sky130_fd_sc_hd__nand3_2
XFILLER_111_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _09410_/A _09408_/Y _09409_/C _09791_/B vssd1 vssd1 vccd1 vccd1 _09548_/A
+ sky130_fd_sc_hd__and4bb_2
X_10681_ _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__xnor2_4
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12421_/A _12421_/B _12421_/C vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__a21o_4
XFILLER_138_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _12351_/A _12351_/B _12350_/X vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__or3b_1
XFILLER_154_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _11302_/A _11302_/B vssd1 vssd1 vccd1 vccd1 _16295_/A sky130_fd_sc_hd__xor2_2
XFILLER_193_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15070_ _14888_/C _14876_/D _14877_/Y _15069_/X vssd1 vssd1 vccd1 vccd1 _15071_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _12283_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__and2_2
XFILLER_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _14021_/A _14021_/B vssd1 vssd1 vccd1 vccd1 _14022_/B sky130_fd_sc_hd__or2_1
XFILLER_141_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11233_ _11155_/A _11154_/C _11154_/A vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__o21a_1
XFILLER_84_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_994 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11165_/C sky130_fd_sc_hd__nor2_1
XFILLER_161_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10115_ _10115_/A _10241_/B _10490_/C _10490_/D vssd1 vssd1 vccd1 vccd1 _10116_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15972_ _15972_/A _15972_/B vssd1 vssd1 vccd1 vccd1 _15973_/B sky130_fd_sc_hd__and2_1
X_11095_ _11095_/A _11240_/A _11423_/C _11605_/B vssd1 vssd1 vccd1 vccd1 _11098_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_96_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10162_/C sky130_fd_sc_hd__xnor2_2
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14923_ _15131_/A _14922_/X _10647_/C vssd1 vssd1 vccd1 vccd1 _14923_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14854_ _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15811_/B sky130_fd_sc_hd__and2_1
XFILLER_36_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _13805_/A _13805_/B vssd1 vssd1 vccd1 vccd1 _13806_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17573_ fanout939/X _17573_/D vssd1 vssd1 vccd1 vccd1 _17573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11997_ _11998_/A _11998_/B _12197_/B _11998_/D vssd1 vssd1 vccd1 vccd1 _11997_/Y
+ sky130_fd_sc_hd__nor4_4
X_14785_ _14785_/A _15541_/A vssd1 vssd1 vccd1 vccd1 _14785_/X sky130_fd_sc_hd__or2_2
X_16524_ _16524_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16525_/B sky130_fd_sc_hd__and2_1
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13736_ _13736_/A _13849_/A vssd1 vssd1 vccd1 vccd1 _13739_/A sky130_fd_sc_hd__nor2_2
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10948_ _10927_/X _11059_/A _10946_/X _10947_/Y vssd1 vssd1 vccd1 vccd1 _10951_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_32_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16455_ _16455_/A _16455_/B vssd1 vssd1 vccd1 vccd1 _16457_/B sky130_fd_sc_hd__xnor2_1
X_13667_ _13668_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13778_/B sky130_fd_sc_hd__nor2_2
X_10879_ _10879_/A _10879_/B vssd1 vssd1 vccd1 vccd1 _11114_/B sky130_fd_sc_hd__xnor2_4
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15406_/A _15406_/B vssd1 vssd1 vccd1 vccd1 _15408_/C sky130_fd_sc_hd__xor2_1
X_12618_ _12618_/A _12770_/B _12770_/D _12618_/D vssd1 vssd1 vccd1 vccd1 _12619_/B
+ sky130_fd_sc_hd__and4_1
X_16386_ _17131_/A _16386_/B vssd1 vssd1 vccd1 vccd1 _16386_/Y sky130_fd_sc_hd__nand2_2
X_13598_ _13598_/A _13598_/B vssd1 vssd1 vccd1 vccd1 _13600_/B sky130_fd_sc_hd__or2_1
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15337_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15346_/A sky130_fd_sc_hd__xnor2_4
X_12549_ _13516_/S _12547_/X _12548_/Y vssd1 vssd1 vccd1 vccd1 _12549_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _17490_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15268_ _15337_/A _15268_/B vssd1 vssd1 vccd1 vccd1 _15281_/A sky130_fd_sc_hd__nand2_4
XFILLER_144_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17007_ _17007_/A _17007_/B vssd1 vssd1 vccd1 vccd1 _17037_/B sky130_fd_sc_hd__xnor2_4
X_14219_ _14297_/A _14219_/B vssd1 vssd1 vccd1 vccd1 _14221_/C sky130_fd_sc_hd__and2_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15199_ _14887_/B _15198_/X _14924_/A vssd1 vssd1 vccd1 vccd1 _15199_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_141_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout508 _17517_/Q vssd1 vssd1 vccd1 vccd1 _09748_/B sky130_fd_sc_hd__buf_6
XFILLER_140_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout519 _14788_/A vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__buf_4
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _09762_/B _09891_/A _09762_/A vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__a21oi_4
XFILLER_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__nor2_2
XFILLER_55_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09125_ _12174_/B _12127_/D _11920_/D _12174_/A vssd1 vssd1 vccd1 vccd1 _09128_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09056_ _17381_/A _12565_/D _08916_/A _08914_/Y vssd1 vssd1 vccd1 vccd1 _09057_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_191_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_190_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09958_ _09770_/Y _09830_/X _09915_/A _10059_/A vssd1 vssd1 vccd1 vccd1 _09960_/C
+ sky130_fd_sc_hd__a211o_4
XTAP_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _08910_/A _08910_/B _08910_/C vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__a21o_2
XFILLER_44_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09765_/X _09887_/Y _09885_/A _09869_/X vssd1 vssd1 vccd1 vccd1 _09912_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11920_ _12770_/A _11920_/B _12127_/D _11920_/D vssd1 vssd1 vccd1 vccd1 _12179_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _12700_/D _11851_/B vssd1 vssd1 vccd1 vccd1 _11852_/B sky130_fd_sc_hd__nand2_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10802_ _10802_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__nor2_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14570_/A _14621_/A _14570_/C vssd1 vssd1 vccd1 vccd1 _14621_/B sky130_fd_sc_hd__nand3_4
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _17476_/D _17477_/D vssd1 vssd1 vccd1 vccd1 _14924_/C sky130_fd_sc_hd__nand2b_4
XFILLER_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _13844_/B _14002_/B _14155_/B _13844_/A vssd1 vssd1 vccd1 vccd1 _13524_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _10714_/X _10728_/B _10732_/Y _10662_/X vssd1 vssd1 vccd1 vccd1 _10771_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_41_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16240_ _16241_/A _16241_/B _16239_/Y vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__o21ba_1
X_13452_ _14387_/A _14052_/B _13453_/C vssd1 vssd1 vccd1 vccd1 _13454_/A sky130_fd_sc_hd__a21oi_1
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10664_ _10670_/A _10636_/Y _10651_/Y _10662_/X vssd1 vssd1 vccd1 vccd1 _10665_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_186_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12403_ _12403_/A _12403_/B vssd1 vssd1 vccd1 vccd1 _17579_/D sky130_fd_sc_hd__nand2_1
XFILLER_173_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16171_ _16171_/A _16352_/B vssd1 vssd1 vccd1 vccd1 _16172_/B sky130_fd_sc_hd__nand2_4
XFILLER_154_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ _13504_/B _13382_/X _13261_/A _13263_/A vssd1 vssd1 vccd1 vccd1 _13509_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_167_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10595_ _10595_/A _10595_/B vssd1 vssd1 vccd1 vccd1 _10709_/B sky130_fd_sc_hd__xnor2_4
XFILLER_127_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12334_ _12500_/A _12638_/B _12334_/C vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__and3_2
X_15122_ _15056_/A _10543_/C _11841_/X _15131_/A _15121_/X vssd1 vssd1 vccd1 vccd1
+ _15126_/B sky130_fd_sc_hd__o311a_1
XFILLER_154_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15053_ _11650_/X _11675_/C _11655_/A _15052_/Y vssd1 vssd1 vccd1 vccd1 _15053_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12265_ _12437_/A _12265_/B _12265_/C vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__nand3_4
XFILLER_135_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _14092_/B _14004_/B vssd1 vssd1 vccd1 vccd1 _14007_/A sky130_fd_sc_hd__nand2_2
X_11216_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__xor2_4
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12196_ _12360_/B _12194_/X _11949_/Y _11997_/Y vssd1 vssd1 vccd1 vccd1 _12198_/B
+ sky130_fd_sc_hd__a211oi_4
Xoutput71 _17466_/Q vssd1 vssd1 vccd1 vccd1 leds[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput82 _17475_/Q vssd1 vssd1 vccd1 vccd1 leds[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput93 _17452_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[18] sky130_fd_sc_hd__clkbuf_2
X_11147_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11154_/A sky130_fd_sc_hd__or2_4
XFILLER_150_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15955_ _16619_/A _15956_/B vssd1 vssd1 vccd1 vccd1 _15955_/Y sky130_fd_sc_hd__nor2_2
X_11078_ _10895_/A _10864_/Y _10881_/Y _11112_/A vssd1 vssd1 vccd1 vccd1 _11080_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14906_ _14906_/A _14906_/B _15175_/B vssd1 vssd1 vccd1 vccd1 _14906_/X sky130_fd_sc_hd__or3_1
X_10029_ _10029_/A _10029_/B _10029_/C vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__or3_2
X_15886_ _15884_/Y _15885_/Y _15523_/A vssd1 vssd1 vccd1 vccd1 _15886_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14837_ _14837_/A _17070_/B vssd1 vssd1 vccd1 vccd1 _14837_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17556_ fanout939/X _17556_/D vssd1 vssd1 vccd1 vccd1 _17556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_189_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14768_ _17415_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _16970_/B sky130_fd_sc_hd__or2_1
X_16507_ _16507_/A _16507_/B vssd1 vssd1 vccd1 vccd1 _16509_/C sky130_fd_sc_hd__xnor2_2
XFILLER_60_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ _13720_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13824_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17487_ fanout931/X _17487_/D vssd1 vssd1 vccd1 vccd1 _17487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14699_ _14699_/A _14699_/B vssd1 vssd1 vccd1 vccd1 _14701_/B sky130_fd_sc_hd__xor2_2
XFILLER_176_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16438_ _16439_/A _16439_/B vssd1 vssd1 vccd1 vccd1 _16527_/B sky130_fd_sc_hd__nor2_2
XFILLER_191_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16369_ _16369_/A _16369_/B vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__xor2_4
XFILLER_158_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _17613_/Q vssd1 vssd1 vccd1 vccd1 _15147_/A sky130_fd_sc_hd__clkbuf_8
Xfanout316 _14832_/A vssd1 vssd1 vccd1 vccd1 _14050_/A sky130_fd_sc_hd__buf_6
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout327 _14708_/B vssd1 vssd1 vccd1 vccd1 _14593_/B sky130_fd_sc_hd__buf_6
X_09812_ _09812_/A _09812_/B _09812_/C vssd1 vssd1 vccd1 vccd1 _09813_/C sky130_fd_sc_hd__or3_2
XFILLER_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout338 _14765_/A vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__buf_6
Xfanout349 _13977_/B vssd1 vssd1 vccd1 vccd1 _14599_/B sky130_fd_sc_hd__buf_8
X_09743_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09743_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09674_ _09674_/A _09674_/B _09819_/A vssd1 vssd1 vccd1 vccd1 _09675_/C sky130_fd_sc_hd__nor3_2
XFILLER_55_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09108_ _09108_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09110_/B sky130_fd_sc_hd__xnor2_1
XFILLER_108_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10380_ _10487_/A _10379_/B _10379_/A vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__o21ba_1
XFILLER_184_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09039_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__xnor2_4
XFILLER_108_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ _16014_/A _15898_/A _12060_/S vssd1 vssd1 vccd1 vccd1 _12051_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11001_ _10977_/X _11051_/A _10999_/X _11000_/Y vssd1 vssd1 vccd1 vccd1 _11157_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout850 _10912_/C vssd1 vssd1 vccd1 vccd1 _10490_/D sky130_fd_sc_hd__buf_6
Xfanout861 _17306_/A1 vssd1 vssd1 vccd1 vccd1 _10805_/C sky130_fd_sc_hd__buf_8
Xfanout872 _10805_/D vssd1 vssd1 vccd1 vccd1 _10957_/D sky130_fd_sc_hd__buf_6
XFILLER_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout883 _17480_/Q vssd1 vssd1 vccd1 vccd1 _10809_/D sky130_fd_sc_hd__buf_8
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout894 _11370_/C vssd1 vssd1 vccd1 vccd1 _11423_/C sky130_fd_sc_hd__buf_6
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15740_ _15740_/A _15740_/B vssd1 vssd1 vccd1 vccd1 _15741_/B sky130_fd_sc_hd__xor2_4
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12952_ _13092_/B _12952_/B vssd1 vssd1 vccd1 vccd1 _12955_/B sky130_fd_sc_hd__nand2_1
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11903_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11906_/A sky130_fd_sc_hd__xnor2_2
X_15671_ _15671_/A _15671_/B vssd1 vssd1 vccd1 vccd1 _15673_/B sky130_fd_sc_hd__xor2_4
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12884_/A _12884_/B vssd1 vssd1 vccd1 vccd1 _13033_/B sky130_fd_sc_hd__nand2b_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17410_ input51/X _17422_/A2 _17409_/X _17414_/C1 vssd1 vssd1 vccd1 vccd1 _17533_/D
+ sky130_fd_sc_hd__o211a_1
X_14622_ _14661_/A _14622_/B vssd1 vssd1 vccd1 vccd1 _14624_/B sky130_fd_sc_hd__or2_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _13067_/C _10839_/D _11839_/S vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__mux2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ input50/X _17359_/B _17359_/C vssd1 vssd1 vccd1 vccd1 _17341_/X sky130_fd_sc_hd__or3_1
X_14553_ _14553_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14555_/A sky130_fd_sc_hd__nor2_1
X_11765_ _16568_/A _11760_/X _11764_/X vssd1 vssd1 vccd1 vccd1 _16866_/B sky130_fd_sc_hd__a21oi_4
XFILLER_159_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10716_ _10716_/A _10716_/B vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__xnor2_4
X_13504_ _13504_/A _13504_/B vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__or2_1
X_17272_ _17458_/Q _17293_/A2 _17270_/X _17271_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17458_/D sky130_fd_sc_hd__o221a_1
X_14484_ _14593_/B _14428_/B _14485_/D _14593_/A vssd1 vssd1 vccd1 vccd1 _14486_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_158_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11696_ _15525_/A _15447_/A _11672_/Y _11624_/Y vssd1 vssd1 vccd1 vccd1 _15614_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_187_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16223_ _16205_/X _16207_/X _16222_/Y _16806_/A2 _14859_/B vssd1 vssd1 vccd1 vccd1
+ _16224_/A sky130_fd_sc_hd__a32o_2
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13435_ _13435_/A _13586_/A vssd1 vssd1 vccd1 vccd1 _13438_/A sky130_fd_sc_hd__or2_1
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _10648_/A _10646_/Y _10647_/C _10647_/D vssd1 vssd1 vccd1 vccd1 _10742_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_139_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16154_ _16155_/A _16155_/B vssd1 vssd1 vccd1 vccd1 _16270_/A sky130_fd_sc_hd__nor2_1
X_13366_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__xnor2_2
XFILLER_177_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10578_ _10325_/A _10329_/B _10579_/A _10577_/X vssd1 vssd1 vccd1 vccd1 _10579_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15105_ _11679_/A _11679_/B _16389_/A vssd1 vssd1 vccd1 vccd1 _15106_/B sky130_fd_sc_hd__o21a_1
XFILLER_155_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12317_ _12186_/A _12186_/B _12189_/A vssd1 vssd1 vccd1 vccd1 _12357_/A sky130_fd_sc_hd__o21ai_4
XFILLER_177_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16085_ _16197_/A _16085_/B vssd1 vssd1 vccd1 vccd1 _16086_/C sky130_fd_sc_hd__and2b_1
X_13297_ _13643_/A _13908_/B _13159_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13304_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_142_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12248_ _12429_/B _12248_/B vssd1 vssd1 vccd1 vccd1 _12250_/B sky130_fd_sc_hd__and2b_4
X_15036_ _14949_/Y _14952_/Y _15038_/A vssd1 vssd1 vccd1 vccd1 _15037_/B sky130_fd_sc_hd__mux2_1
XFILLER_123_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12179_ _12179_/A _12179_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12180_/B sky130_fd_sc_hd__nor3_2
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16987_ _17119_/A _17043_/B vssd1 vssd1 vccd1 vccd1 _16989_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15938_ _15939_/A _15939_/B vssd1 vssd1 vccd1 vccd1 _16072_/B sky130_fd_sc_hd__and2_2
XFILLER_149_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15869_ _15414_/B _15746_/X _15750_/X vssd1 vssd1 vccd1 vccd1 _15871_/B sky130_fd_sc_hd__o21ba_1
XFILLER_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17608_ fanout925/X _17608_/D vssd1 vssd1 vccd1 vccd1 _17608_/Q sky130_fd_sc_hd__dfxtp_4
X_09390_ _09343_/X _09344_/Y _09387_/A _09388_/Y vssd1 vssd1 vccd1 vccd1 _09393_/C
+ sky130_fd_sc_hd__o211a_4
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17539_ fanout944/X _17539_/D vssd1 vssd1 vccd1 vccd1 _17539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout124 _17229_/B vssd1 vssd1 vccd1 vccd1 _17292_/B sky130_fd_sc_hd__clkbuf_4
Xfanout135 _15199_/Y vssd1 vssd1 vccd1 vccd1 _16536_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_945 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout146 _15749_/A vssd1 vssd1 vccd1 vccd1 _16165_/A sky130_fd_sc_hd__buf_6
XFILLER_87_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout157 _17384_/A2 vssd1 vssd1 vccd1 vccd1 _17426_/A2 sky130_fd_sc_hd__buf_2
Xfanout168 _16030_/B vssd1 vssd1 vccd1 vccd1 _16662_/D sky130_fd_sc_hd__buf_4
XFILLER_102_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout179 _15551_/Y vssd1 vssd1 vccd1 vccd1 _16758_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09726_ _11902_/A _09892_/C _09587_/A _09585_/Y vssd1 vssd1 vccd1 vccd1 _09727_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ _09786_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09658_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09589_/B _09589_/A vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__and2b_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ _11542_/A _11541_/C _11541_/A vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__o21a_2
XFILLER_156_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10501_ _10501_/A _10501_/B vssd1 vssd1 vccd1 vccd1 _10503_/C sky130_fd_sc_hd__xnor2_2
XFILLER_184_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11481_ _11561_/B _11480_/C _11561_/C _11480_/A vssd1 vssd1 vccd1 vccd1 _11481_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_183_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13220_ _13220_/A _13220_/B _13220_/C vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__nand3_1
XFILLER_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10432_ _10431_/A _10545_/D _10180_/C vssd1 vssd1 vccd1 vccd1 _10432_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13151_ _13151_/A _13151_/B vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__xnor2_2
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__nor2_2
XFILLER_88_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12102_ _17379_/A _12270_/B _12270_/D _12102_/D vssd1 vssd1 vccd1 vccd1 _12103_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13082_ _13083_/A _13213_/A _13083_/C vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__o21a_1
XFILLER_3_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10294_ _15711_/A _10657_/B _10288_/A _10172_/Y vssd1 vssd1 vccd1 vccd1 _10296_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16910_ _16910_/A _16910_/B vssd1 vssd1 vccd1 vccd1 _16911_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _08969_/C _12032_/Y _12700_/D vssd1 vssd1 vccd1 vccd1 _12033_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16841_ _16841_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16843_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout680 _14863_/A vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__buf_4
XFILLER_59_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout691 _17500_/Q vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__buf_6
X_16772_ _16688_/A _16687_/B _16685_/X vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__a21o_1
X_13984_ _13985_/B _13985_/A vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15723_ _15816_/A _16747_/A vssd1 vssd1 vccd1 vccd1 _15730_/A sky130_fd_sc_hd__nor2_4
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12935_ _12935_/A _12935_/B vssd1 vssd1 vccd1 vccd1 _12938_/C sky130_fd_sc_hd__or2_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15654_ _15743_/A _15654_/B vssd1 vssd1 vccd1 vccd1 _15656_/B sky130_fd_sc_hd__nor2_2
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _14421_/S _12866_/B vssd1 vssd1 vccd1 vccd1 _12866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _14606_/B _14606_/A vssd1 vssd1 vccd1 vccd1 _14646_/B sky130_fd_sc_hd__nand2b_2
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _11814_/Y _11816_/Y _17365_/A vssd1 vssd1 vccd1 vccd1 _11818_/B sky130_fd_sc_hd__mux2_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _15499_/A _15499_/B _15488_/Y vssd1 vssd1 vccd1 vccd1 _15587_/B sky130_fd_sc_hd__o21ai_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12798_/A _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12799_/A sky130_fd_sc_hd__a21oi_4
XFILLER_14_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _13434_/D _17328_/A2 _17323_/X _17392_/C1 vssd1 vssd1 vccd1 vccd1 _17491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14536_ _14415_/X _14534_/B _14534_/Y _14280_/X vssd1 vssd1 vccd1 vccd1 _14536_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11748_ _16794_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _16727_/B sky130_fd_sc_hd__and2_2
XFILLER_159_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_186_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17255_ _17594_/Q _17291_/A2 _17291_/B1 vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__a21o_1
X_14467_ _14524_/A _14524_/B vssd1 vssd1 vccd1 vccd1 _14469_/B sky130_fd_sc_hd__xnor2_2
XFILLER_147_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11679_ _11679_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _15106_/A sky130_fd_sc_hd__nand2_1
X_16206_ _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16207_/C sky130_fd_sc_hd__nor2_1
X_13418_ _13418_/A _13418_/B vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__and2_2
X_17186_ input29/X wire217/X vssd1 vssd1 vccd1 vccd1 _17429_/B sky130_fd_sc_hd__nand2_1
X_14398_ _14395_/Y _14396_/X _14316_/A _14332_/X vssd1 vssd1 vccd1 vccd1 _14400_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_161_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16137_ _16137_/A _16250_/A vssd1 vssd1 vccd1 vccd1 _16140_/A sky130_fd_sc_hd__or2_2
XFILLER_142_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _13349_/A _13349_/B vssd1 vssd1 vccd1 vccd1 _13368_/A sky130_fd_sc_hd__xnor2_4
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16068_ _16068_/A _16068_/B vssd1 vssd1 vccd1 vccd1 _16070_/B sky130_fd_sc_hd__xor2_2
XFILLER_69_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ _14906_/A _14899_/C _15018_/X _15143_/A vssd1 vssd1 vccd1 vccd1 _15402_/B
+ sky130_fd_sc_hd__o22ai_4
X_08890_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _08904_/C sky130_fd_sc_hd__nand2_1
XFILLER_69_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_97_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_1035 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1019 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09511_ _09511_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _11902_/A _11870_/B _09302_/A _09300_/Y vssd1 vssd1 vccd1 vccd1 _09443_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09373_/A _09373_/B vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__nor2_4
XFILLER_52_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _09709_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__xnor2_4
Xwb_buttons_leds_954 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_954/HI led_enb[7] sky130_fd_sc_hd__conb_1
X_10981_ _10974_/A _10973_/B _10973_/A vssd1 vssd1 vccd1 vccd1 _10985_/A sky130_fd_sc_hd__o21ba_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12720_ _12720_/A _12720_/B vssd1 vssd1 vccd1 vccd1 _12727_/A sky130_fd_sc_hd__xor2_1
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12651_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11602_ _11568_/A _11568_/C _11568_/B vssd1 vssd1 vccd1 vccd1 _11603_/C sky130_fd_sc_hd__a21oi_1
XFILLER_168_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12582_ _12583_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12761_/B sky130_fd_sc_hd__and2b_1
X_15370_ _11692_/B _11691_/B _11693_/Y vssd1 vssd1 vccd1 vccd1 _15370_/X sky130_fd_sc_hd__a21o_1
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14321_ _14387_/A _14599_/D _14321_/C vssd1 vssd1 vccd1 vccd1 _14389_/B sky130_fd_sc_hd__and3_1
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ _11534_/A _11534_/B vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__or2_4
XFILLER_168_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _17040_/A _17040_/B vssd1 vssd1 vccd1 vccd1 _17085_/A sky130_fd_sc_hd__nor2_2
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ _14252_/A _14252_/B _14252_/C vssd1 vssd1 vccd1 vccd1 _14253_/B sky130_fd_sc_hd__and3_1
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11464_ _11708_/A _11464_/B vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__or2_4
XFILLER_183_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10415_ _10415_/A _10513_/A vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__nor2_4
XFILLER_99_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13203_ _13203_/A vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__inv_2
X_14183_ _14273_/B _14184_/C vssd1 vssd1 vccd1 vccd1 _14185_/B sky130_fd_sc_hd__and2_1
X_11395_ _11395_/A _11395_/B _11435_/A vssd1 vssd1 vccd1 vccd1 _11396_/C sky130_fd_sc_hd__nand3_2
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _17105_/A sky130_fd_sc_hd__nor2_1
X_13134_ _13137_/A vssd1 vssd1 vccd1 vccd1 _13134_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13065_ _13065_/A _13065_/B _13065_/C vssd1 vssd1 vccd1 vccd1 _13075_/B sky130_fd_sc_hd__nand3_2
X_10277_ _14788_/A _10534_/D _10167_/A _10165_/Y vssd1 vssd1 vccd1 vccd1 _10278_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_105_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ _12016_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__nand2_1
XFILLER_94_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16824_ _16935_/A _16760_/B _16761_/A _16759_/B vssd1 vssd1 vccd1 vccd1 _16830_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_78_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _16661_/X _16665_/B _16663_/B vssd1 vssd1 vccd1 vccd1 _16762_/A sky130_fd_sc_hd__o21ai_2
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13967_ _13967_/A _13967_/B vssd1 vssd1 vccd1 vccd1 _13969_/A sky130_fd_sc_hd__nor2_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15706_ _15705_/A _15705_/B _15705_/C vssd1 vssd1 vccd1 vccd1 _15706_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12918_ _13065_/A _12918_/B _12918_/C vssd1 vssd1 vccd1 vccd1 _13065_/B sky130_fd_sc_hd__nand3_4
X_16686_ _16686_/A _16686_/B _16684_/Y vssd1 vssd1 vccd1 vccd1 _16687_/B sky130_fd_sc_hd__or3b_1
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13898_ _13898_/A _13898_/B vssd1 vssd1 vccd1 vccd1 _13901_/B sky130_fd_sc_hd__xnor2_2
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15637_ _16108_/C _15071_/A _15262_/A vssd1 vssd1 vccd1 vccd1 _15639_/B sky130_fd_sc_hd__a21bo_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _13838_/S _12849_/B vssd1 vssd1 vccd1 vccd1 _12849_/X sky130_fd_sc_hd__or2_1
XFILLER_15_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15568_ _15568_/A _15568_/B vssd1 vssd1 vccd1 vccd1 _15570_/A sky130_fd_sc_hd__and2_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17307_ input63/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17307_/X sky130_fd_sc_hd__or3_1
X_14519_ _14519_/A _14519_/B _14519_/C vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__and3_4
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15499_ _15499_/A _15499_/B vssd1 vssd1 vccd1 vccd1 _15501_/C sky130_fd_sc_hd__xor2_2
XFILLER_175_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17238_ _17556_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__and2_1
XFILLER_128_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_115_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17169_ _17169_/A1 _17167_/X _17168_/Y _17166_/X vssd1 vssd1 vccd1 vccd1 _17169_/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09991_ _10004_/B _10004_/C _10004_/A vssd1 vssd1 vccd1 vccd1 _09991_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_142_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08942_ _11932_/A _12270_/C vssd1 vssd1 vccd1 vccd1 _08943_/B sky130_fd_sc_hd__nand2_2
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08873_ _08874_/A _08874_/B _08873_/C _08873_/D vssd1 vssd1 vccd1 vccd1 _08873_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09425_ _11791_/C _09712_/B vssd1 vssd1 vccd1 vccd1 _16933_/A sky130_fd_sc_hd__nand2_8
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09366_/B sky130_fd_sc_hd__nand2b_2
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09287_ _09421_/A _09285_/X _17081_/B _16990_/A vssd1 vssd1 vccd1 vccd1 _09289_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_107_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__nor2_2
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11180_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11181_/B sky130_fd_sc_hd__xor2_4
XFILLER_122_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ _10132_/B _10132_/A vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__nand2b_2
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10062_ _10062_/A _10062_/B _10062_/C vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__and3_4
XFILLER_48_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14870_ _14831_/Y _17151_/B _16485_/A _14869_/X vssd1 vssd1 vccd1 vccd1 _17575_/D
+ sky130_fd_sc_hd__a31o_2
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13821_ _14254_/A _14865_/B _13705_/A _13703_/A vssd1 vssd1 vccd1 vccd1 _13823_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ _16627_/A vssd1 vssd1 vccd1 vccd1 _16542_/A sky130_fd_sc_hd__inv_2
X_13752_ _13642_/A _13644_/B _13642_/B vssd1 vssd1 vccd1 vccd1 _13754_/B sky130_fd_sc_hd__o21ba_1
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10964_ _10963_/B _10911_/B _10963_/D _10963_/A vssd1 vssd1 vccd1 vccd1 _10965_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ _12701_/Y _12702_/X _13627_/S vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__mux2_1
X_16471_ _16470_/A _16470_/B _16470_/C vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__a21oi_2
X_13683_ _13683_/A _13683_/B vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__xor2_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10895_ _10895_/A _11080_/A vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__and2_2
XFILLER_71_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15422_ _15422_/A _15422_/B vssd1 vssd1 vccd1 vccd1 _15424_/B sky130_fd_sc_hd__xor2_4
X_12634_ _12518_/A _12518_/B _12516_/Y vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__a21bo_2
XFILLER_70_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15353_ _15278_/A _15397_/A _15279_/A _15276_/Y vssd1 vssd1 vccd1 vccd1 _15355_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_184_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12565_ _17397_/A _17395_/A _12565_/C _12565_/D vssd1 vssd1 vccd1 vccd1 _12566_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14304_ _14304_/A _14304_/B vssd1 vssd1 vccd1 vccd1 _14306_/B sky130_fd_sc_hd__xnor2_4
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11523_/A sky130_fd_sc_hd__nor2_2
XFILLER_102_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15284_ _15285_/A _15285_/B vssd1 vssd1 vccd1 vccd1 _15352_/A sky130_fd_sc_hd__or2_4
XFILLER_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12496_ _12496_/A _12496_/B vssd1 vssd1 vccd1 vccd1 _12498_/C sky130_fd_sc_hd__xor2_1
XFILLER_144_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17023_ _17023_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _17024_/B sky130_fd_sc_hd__nand2_1
X_14235_ _14235_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14236_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ _11447_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__nand2_1
XFILLER_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14166_ _14318_/B _14545_/C _14545_/D _14450_/A vssd1 vssd1 vccd1 vccd1 _14170_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11378_ _11553_/B _14906_/B vssd1 vssd1 vccd1 vccd1 _11380_/B sky130_fd_sc_hd__nand2_1
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10450_/A _10329_/B _10329_/C vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__and3_4
X_13117_ _13117_/A _13117_/B _13117_/C vssd1 vssd1 vccd1 vccd1 _13118_/B sky130_fd_sc_hd__nand3_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14098_/A _14098_/B vssd1 vssd1 vccd1 vccd1 _14188_/B sky130_fd_sc_hd__or2_4
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13048_ _13049_/A _13049_/B _13049_/C vssd1 vssd1 vccd1 vccd1 _13061_/A sky130_fd_sc_hd__a21o_4
XFILLER_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1046 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_935 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16807_ _16807_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16811_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14999_ _15100_/A _14999_/B vssd1 vssd1 vccd1 vccd1 _14999_/Y sky130_fd_sc_hd__nand2_1
X_16738_ _16389_/A _16794_/B _16728_/Y _16737_/X vssd1 vssd1 vccd1 vccd1 _16738_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_62_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16669_ _16667_/A _16938_/D _16670_/A _16814_/A _16813_/B vssd1 vssd1 vccd1 vccd1
+ _16671_/B sky130_fd_sc_hd__o32a_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09210_ _09211_/B _09373_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__o21a_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09141_ _12174_/B _12127_/C _12127_/D _12174_/A vssd1 vssd1 vccd1 vccd1 _09143_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_147_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _09071_/A _09259_/A _08930_/X _09018_/Y vssd1 vssd1 vccd1 vccd1 _09119_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_190_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _09885_/A _09885_/B _09885_/C vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__a21oi_2
X_08925_ _09012_/A _08910_/Y _08917_/X _09053_/A vssd1 vssd1 vccd1 vccd1 _08927_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_58_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08856_ _08856_/A _08856_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08787_ _08798_/A _08787_/B _12258_/A _11881_/D vssd1 vssd1 vccd1 vccd1 _08821_/A
+ sky130_fd_sc_hd__and4b_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09408_ _09407_/B _09647_/B _09937_/B _09838_/A vssd1 vssd1 vccd1 vccd1 _09408_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10673_/A _10673_/B _10674_/Y vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__a21oi_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09339_ _09339_/A _09344_/B _09339_/C vssd1 vssd1 vccd1 vccd1 _09391_/C sky130_fd_sc_hd__or3_4
XFILLER_178_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12350_ _12517_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__and2_1
XFILLER_193_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11301_ _11711_/A _11711_/B vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__and2b_1
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12281_ _12281_/A _12281_/B vssd1 vssd1 vccd1 vccd1 _12283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14020_ _14021_/A _14021_/B vssd1 vssd1 vccd1 vccd1 _14113_/B sky130_fd_sc_hd__nand2_1
X_11232_ _11232_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__xnor2_4
XFILLER_49_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _14794_/A _09892_/C _10756_/A _10754_/Y vssd1 vssd1 vccd1 vccd1 _11165_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10114_ _10241_/B _10490_/C _10490_/D _10694_/A vssd1 vssd1 vccd1 vccd1 _10116_/A
+ sky130_fd_sc_hd__a22oi_4
X_15971_ _15972_/A _15972_/B vssd1 vssd1 vccd1 vccd1 _16080_/B sky130_fd_sc_hd__nor2_4
X_11094_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10045_ _10162_/A _10044_/Y _15711_/A _10543_/B vssd1 vssd1 vccd1 vccd1 _10170_/A
+ sky130_fd_sc_hd__and4bb_4
XFILLER_49_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14922_ _14920_/X _14921_/X _14922_/S vssd1 vssd1 vccd1 vccd1 _14922_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14853_ _15624_/A _15541_/A _15541_/B vssd1 vssd1 vccd1 vccd1 _15709_/B sky130_fd_sc_hd__and3_2
XFILLER_17_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13804_ _13805_/A _13805_/B vssd1 vssd1 vccd1 vccd1 _13915_/B sky130_fd_sc_hd__and2_1
XFILLER_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17572_ fanout945/X _17572_/D vssd1 vssd1 vccd1 vccd1 _17572_/Q sky130_fd_sc_hd__dfxtp_1
X_14784_ _14784_/A _15624_/A vssd1 vssd1 vccd1 vccd1 _15622_/B sky130_fd_sc_hd__or2_2
X_11996_ _12197_/A _11994_/X _09248_/B _09248_/Y vssd1 vssd1 vccd1 vccd1 _11998_/D
+ sky130_fd_sc_hd__o211a_4
XFILLER_1_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16523_ _16524_/A _16524_/B vssd1 vssd1 vccd1 vccd1 _16616_/B sky130_fd_sc_hd__nor2_2
X_13735_ _13844_/A _13844_/B _13948_/D _14002_/B vssd1 vssd1 vccd1 vccd1 _13849_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10947_ _10946_/A _10946_/B _10946_/C vssd1 vssd1 vccd1 vccd1 _10947_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16454_ _16454_/A _16454_/B vssd1 vssd1 vccd1 vccd1 _16455_/B sky130_fd_sc_hd__xor2_2
XFILLER_182_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13666_ _14215_/A _13764_/C vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__nand2_1
X_10878_ _10878_/A _11121_/A vssd1 vssd1 vccd1 vccd1 _11114_/A sky130_fd_sc_hd__or2_4
XFILLER_188_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15405_ _16315_/C _16262_/A vssd1 vssd1 vccd1 vccd1 _15406_/B sky130_fd_sc_hd__nor2_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12770_/B _12465_/B _12618_/D _12618_/A vssd1 vssd1 vccd1 vccd1 _12619_/A
+ sky130_fd_sc_hd__a22oi_4
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _16385_/A _16385_/B vssd1 vssd1 vccd1 vccd1 _16386_/B sky130_fd_sc_hd__xor2_4
X_13597_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _13598_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15336_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15336_/Y sky130_fd_sc_hd__nand2_1
X_12548_ _13516_/S _12548_/B vssd1 vssd1 vccd1 vccd1 _12548_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_185_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15267_ _15918_/A _16536_/A _16533_/A _15726_/A vssd1 vssd1 vccd1 vccd1 _15268_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_2 _16103_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12481_/A _12481_/B _12481_/C vssd1 vssd1 vccd1 vccd1 _12479_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17006_ _17007_/A _17007_/B vssd1 vssd1 vccd1 vccd1 _17093_/A sky130_fd_sc_hd__or2_1
X_14218_ _14218_/A _14218_/B _14218_/C vssd1 vssd1 vccd1 vccd1 _14219_/B sky130_fd_sc_hd__or3_1
XFILLER_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15198_ _15147_/A _11789_/X _15393_/B vssd1 vssd1 vccd1 vccd1 _15198_/X sky130_fd_sc_hd__a21o_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_153_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14149_ _14150_/A _14150_/B _14150_/C vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__o21a_1
Xfanout509 _10036_/B vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_63_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09690_ _10366_/A _10490_/C _09552_/A _09550_/Y vssd1 vssd1 vccd1 vccd1 _09696_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_187_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09124_ _11920_/B _12772_/A _09172_/B _17466_/D vssd1 vssd1 vccd1 vccd1 _09167_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_109_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09055_ _09055_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _09055_/Y sky130_fd_sc_hd__nand3_2
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1008 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_135_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__and2_2
XFILLER_106_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ _08908_/A _08908_/B vssd1 vssd1 vccd1 vccd1 _08910_/C sky130_fd_sc_hd__or2_2
XTAP_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09869_/X _09885_/A _09887_/Y _09765_/X vssd1 vssd1 vccd1 vccd1 _09912_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08862_/B _08839_/B vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__nor2_1
XFILLER_45_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11651_/A _11675_/B _11675_/C vssd1 vssd1 vccd1 vccd1 _11851_/B sky130_fd_sc_hd__o21ai_4
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ _11314_/A _10911_/B _10800_/C vssd1 vssd1 vccd1 vccd1 _10802_/B sky130_fd_sc_hd__a21oi_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _12016_/B _11781_/B vssd1 vssd1 vccd1 vccd1 _14837_/A sky130_fd_sc_hd__and2_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13520_ _14840_/A _14637_/A1 _12548_/B _13519_/Y _08718_/A vssd1 vssd1 vccd1 vccd1
+ _13520_/X sky130_fd_sc_hd__a311o_1
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10732_ _10662_/A _10662_/B _10662_/C vssd1 vssd1 vccd1 vccd1 _10732_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13451_ _13451_/A _13569_/A vssd1 vssd1 vccd1 vccd1 _13453_/C sky130_fd_sc_hd__nor2_1
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10663_ _10651_/Y _10662_/X _10670_/A _10636_/Y vssd1 vssd1 vccd1 vccd1 _10670_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_139_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _11849_/A _12396_/X _12401_/X _16653_/A vssd1 vssd1 vccd1 vccd1 _12403_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16170_ _16170_/A _16170_/B vssd1 vssd1 vccd1 vccd1 _16172_/A sky130_fd_sc_hd__nand2_4
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10594_ _11027_/B _17469_/D vssd1 vssd1 vccd1 vccd1 _10595_/B sky130_fd_sc_hd__nand2_2
X_13382_ _13504_/A _13380_/X _13221_/A _13224_/A vssd1 vssd1 vccd1 vccd1 _13382_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15121_ _11841_/A _10899_/D _10897_/C _10993_/C vssd1 vssd1 vccd1 vccd1 _15121_/X
+ sky130_fd_sc_hd__a211o_1
X_12333_ _12333_/A _12333_/B vssd1 vssd1 vccd1 vccd1 _12334_/C sky130_fd_sc_hd__xnor2_1
XFILLER_103_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15052_ _11675_/C _11655_/A _11676_/A vssd1 vssd1 vccd1 vccd1 _15052_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _12437_/A _12265_/B _12265_/C vssd1 vssd1 vccd1 vccd1 _12266_/A sky130_fd_sc_hd__a21o_1
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14003_ _14326_/A _14593_/D _14002_/C vssd1 vssd1 vccd1 vccd1 _14004_/B sky130_fd_sc_hd__a21o_1
XFILLER_123_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11215_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11215_/Y sky130_fd_sc_hd__nor2_1
X_12195_ _11998_/A _11997_/Y _12360_/B _12194_/X vssd1 vssd1 vccd1 vccd1 _12198_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_150_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput72 _17476_/Q vssd1 vssd1 vccd1 vccd1 leds[10] sky130_fd_sc_hd__clkbuf_2
Xoutput83 _17542_/Q vssd1 vssd1 vccd1 vccd1 o_wb_ack sky130_fd_sc_hd__clkbuf_2
X_11146_ _11146_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _11148_/B sky130_fd_sc_hd__and2_1
XFILLER_122_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput94 _17453_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[19] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_62_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15954_ _15954_/A _15954_/B vssd1 vssd1 vccd1 vccd1 _15964_/A sky130_fd_sc_hd__and2_2
X_11077_ _11077_/A _11110_/A _11077_/C vssd1 vssd1 vccd1 vccd1 _11080_/B sky130_fd_sc_hd__or3_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14905_ _15208_/C _15208_/D _14905_/C _14905_/D vssd1 vssd1 vccd1 vccd1 _14905_/X
+ sky130_fd_sc_hd__or4_1
X_10028_ _10028_/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/C sky130_fd_sc_hd__nor2_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15885_ _15788_/Y _15790_/X _15787_/X vssd1 vssd1 vccd1 vccd1 _15885_/Y sky130_fd_sc_hd__a21boi_4
XFILLER_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14836_ _14836_/A _14836_/B _14933_/B vssd1 vssd1 vccd1 vccd1 _16007_/A sky130_fd_sc_hd__nand3_2
XTAP_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ fanout935/X _17555_/D vssd1 vssd1 vccd1 vccd1 _17555_/Q sky130_fd_sc_hd__dfxtp_1
X_14767_ _17415_/A _16974_/A vssd1 vssd1 vccd1 vccd1 _14767_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11979_ _12176_/A _12338_/D vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__nand2_2
XFILLER_147_1040 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16506_ _16503_/A _16670_/A _16504_/Y _16505_/X vssd1 vssd1 vccd1 vccd1 _16507_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_108_1002 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13718_ _13718_/A _13718_/B vssd1 vssd1 vccd1 vccd1 _13720_/B sky130_fd_sc_hd__nand2_2
X_17486_ fanout927/X _17486_/D vssd1 vssd1 vccd1 vccd1 _17486_/Q sky130_fd_sc_hd__dfxtp_1
X_14698_ _14698_/A _14698_/B vssd1 vssd1 vccd1 vccd1 _14699_/B sky130_fd_sc_hd__nand2_1
XFILLER_176_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16437_ _16437_/A _16437_/B vssd1 vssd1 vccd1 vccd1 _16439_/B sky130_fd_sc_hd__xnor2_4
XFILLER_176_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _13749_/B _13648_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13650_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16368_ _16273_/A _16273_/B _16256_/X vssd1 vssd1 vccd1 vccd1 _16369_/B sky130_fd_sc_hd__a21o_2
XFILLER_30_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15319_ _15039_/X _15057_/X _15059_/Y _15061_/Y _15130_/S _15901_/S vssd1 vssd1 vccd1
+ vccd1 _15319_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16299_ _16394_/A _16299_/B vssd1 vssd1 vccd1 vccd1 _16301_/A sky130_fd_sc_hd__nand2_1
XFILLER_173_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout306 _17612_/Q vssd1 vssd1 vccd1 vccd1 _15147_/C sky130_fd_sc_hd__buf_6
XFILLER_193_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout317 _14832_/A vssd1 vssd1 vccd1 vccd1 _14213_/A sky130_fd_sc_hd__buf_4
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__xor2_4
Xfanout328 _17134_/A vssd1 vssd1 vccd1 vccd1 _14708_/B sky130_fd_sc_hd__buf_6
XFILLER_115_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout339 _17538_/Q vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__buf_6
XFILLER_143_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _09812_/B vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__inv_2
XFILLER_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09673_ _10560_/B _09555_/C _09386_/B _09384_/X vssd1 vssd1 vccd1 vccd1 _09675_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_39_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_176_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_164_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09107_ _12772_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09038_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__nand2b_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11000_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _11000_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_46_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout840 _10911_/B vssd1 vssd1 vccd1 vccd1 _10490_/C sky130_fd_sc_hd__buf_6
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout851 _10963_/D vssd1 vssd1 vccd1 vccd1 _10912_/C sky130_fd_sc_hd__buf_12
Xfanout862 _15175_/B vssd1 vssd1 vccd1 vccd1 _14848_/B sky130_fd_sc_hd__buf_4
Xfanout873 _17481_/Q vssd1 vssd1 vccd1 vccd1 _10805_/D sky130_fd_sc_hd__buf_6
Xfanout884 _15401_/A vssd1 vssd1 vccd1 vccd1 _14792_/B sky130_fd_sc_hd__clkbuf_8
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout895 _17479_/Q vssd1 vssd1 vccd1 vccd1 _11370_/C sky130_fd_sc_hd__buf_8
X_12951_ _17407_/A _12950_/B _12950_/C vssd1 vssd1 vccd1 vccd1 _12952_/B sky130_fd_sc_hd__a21o_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11902_/A _12734_/D vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__nand2_2
X_15670_ _15671_/A _15671_/B vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__nand2_2
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _13040_/B _12882_/B vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__and2b_4
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14621_/A _14621_/B _14621_/C vssd1 vssd1 vccd1 vccd1 _14622_/B sky130_fd_sc_hd__and3_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11827_/X _11832_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _11833_/X sky130_fd_sc_hd__mux2_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _12565_/D _17360_/A2 _17339_/X _17406_/C1 vssd1 vssd1 vccd1 vccd1 _17499_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14599_/A _14599_/B _14708_/D _14641_/C vssd1 vssd1 vccd1 vccd1 _14553_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _16727_/B _16795_/A _11762_/X _11763_/Y vssd1 vssd1 vccd1 vccd1 _11764_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13503_/A _13503_/B vssd1 vssd1 vccd1 vccd1 _13506_/A sky130_fd_sc_hd__xnor2_1
X_17271_ _17567_/Q _17286_/B vssd1 vssd1 vccd1 vccd1 _17271_/X sky130_fd_sc_hd__and2_1
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10715_ _10715_/A _10715_/B _10715_/C vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__nand3_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14483_ _08718_/A _14481_/X _14482_/X vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_41_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11695_ _11691_/Y _11693_/Y _11694_/X _11672_/Y vssd1 vssd1 vccd1 vccd1 _15447_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_158_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16222_ _16212_/Y _16213_/X _16221_/X vssd1 vssd1 vccd1 vccd1 _16222_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13434_ _14050_/A _14050_/B _13434_/C _13434_/D vssd1 vssd1 vccd1 vccd1 _13586_/A
+ sky130_fd_sc_hd__and4_1
X_10646_ _10933_/B _10645_/C _10743_/C _10933_/A vssd1 vssd1 vccd1 vccd1 _10646_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16153_ _16153_/A _16153_/B vssd1 vssd1 vccd1 vccd1 _16155_/B sky130_fd_sc_hd__xor2_4
XFILLER_158_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _13366_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13365_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10577_ _10463_/B _10471_/X _10573_/X _10575_/Y vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_177_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15104_ _15715_/B _15103_/X _15901_/S vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _12316_/A _12316_/B _12316_/C vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__nand3_2
X_16084_ _16084_/A _16084_/B _16082_/X vssd1 vssd1 vccd1 vccd1 _16085_/B sky130_fd_sc_hd__or3b_1
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _13170_/A _13172_/B _13170_/B vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__o21ba_4
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ _16011_/C _15034_/Y _15035_/S vssd1 vssd1 vccd1 vccd1 _15627_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12247_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12248_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12178_ _12179_/A _12179_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__o21a_1
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11129_ _11130_/B _11130_/C _11130_/A vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__a21o_1
X_16986_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16991_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15937_ _15937_/A _15937_/B vssd1 vssd1 vccd1 vccd1 _15939_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15868_ _15868_/A _15868_/B vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__or2_1
XFILLER_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17607_ fanout925/X _17607_/D vssd1 vssd1 vccd1 vccd1 _17607_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14819_ _16649_/B _16649_/C _16649_/A vssd1 vssd1 vccd1 vccd1 _16730_/A sky130_fd_sc_hd__a21bo_1
XFILLER_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15799_ _15797_/Y _15798_/Y _15309_/B vssd1 vssd1 vccd1 vccd1 _15799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17538_ fanout937/X _17538_/D vssd1 vssd1 vccd1 vccd1 _17538_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_189_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17469_ fanout928/X _17469_/D vssd1 vssd1 vccd1 vccd1 _17469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout125 _17229_/B vssd1 vssd1 vccd1 vccd1 _17286_/B sky130_fd_sc_hd__clkbuf_4
Xfanout136 _15199_/Y vssd1 vssd1 vccd1 vccd1 _16171_/A sky130_fd_sc_hd__clkbuf_8
Xfanout147 _14969_/Y vssd1 vssd1 vccd1 vccd1 _15918_/A sky130_fd_sc_hd__buf_4
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout158 _17384_/A2 vssd1 vssd1 vccd1 vccd1 _17377_/B sky130_fd_sc_hd__buf_4
XFILLER_102_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout169 _15817_/X vssd1 vssd1 vccd1 vccd1 _17043_/B sky130_fd_sc_hd__buf_4
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09725_ _09725_/A _09725_/B _09725_/C vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__nand3_4
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09656_ _09656_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__or3_4
XFILLER_83_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09587_/A _09727_/A vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__nor2_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _10485_/X _10499_/A _10384_/X _10475_/Y vssd1 vssd1 vccd1 vccd1 _10500_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11480_ _11480_/A _11561_/B _11480_/C _11561_/C vssd1 vssd1 vccd1 vccd1 _11484_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_184_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10431_ _10431_/A _10431_/B _14956_/A vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__and3_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _13950_/A _14215_/B vssd1 vssd1 vccd1 vccd1 _13151_/B sky130_fd_sc_hd__nand2_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10362_ _10374_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__or2_4
XFILLER_109_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12101_ _12270_/B _12270_/D _12102_/D _17379_/A vssd1 vssd1 vccd1 vccd1 _12103_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_3_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10293_ _10293_/A _10399_/A vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__nor2_4
X_13081_ _14771_/A _13966_/D vssd1 vssd1 vccd1 vccd1 _13083_/C sky130_fd_sc_hd__nand2_1
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_105_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _12060_/S _17134_/B vssd1 vssd1 vccd1 vccd1 _12032_/Y sky130_fd_sc_hd__nor2_2
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _16841_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__nand2b_1
Xfanout670 _14864_/A vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__buf_4
Xfanout681 fanout686/X vssd1 vssd1 vccd1 vccd1 _14863_/A sky130_fd_sc_hd__buf_4
X_16771_ _16771_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16775_/A sky130_fd_sc_hd__and2_1
Xfanout692 _13566_/B vssd1 vssd1 vccd1 vccd1 _14213_/C sky130_fd_sc_hd__buf_8
X_13983_ _13878_/A _13880_/B _13878_/B vssd1 vssd1 vccd1 vccd1 _13985_/B sky130_fd_sc_hd__o21ba_4
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15722_ _15206_/A _16977_/A _15721_/X vssd1 vssd1 vccd1 vccd1 _17554_/D sky130_fd_sc_hd__o21a_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12934_ _12933_/A _12933_/B _12933_/C vssd1 vssd1 vccd1 vccd1 _12935_/B sky130_fd_sc_hd__o21a_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15653_ _15742_/A _15742_/B vssd1 vssd1 vccd1 vccd1 _15654_/B sky130_fd_sc_hd__and2_1
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _12390_/X _12393_/B _12865_/S vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__mux2_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14553_/A _14555_/B _14553_/B vssd1 vssd1 vccd1 vccd1 _14606_/B sky130_fd_sc_hd__o21ba_1
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _14981_/A _14978_/B _14912_/B vssd1 vssd1 vccd1 vccd1 _11816_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15584_ _15584_/A _15584_/B vssd1 vssd1 vccd1 vccd1 _15685_/B sky130_fd_sc_hd__xnor2_4
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12796_/A _12796_/B vssd1 vssd1 vccd1 vccd1 _12798_/C sky130_fd_sc_hd__xor2_4
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ input40/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17323_/X sky130_fd_sc_hd__or3_1
XFILLER_186_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14535_ _14414_/A _14475_/A _14533_/B vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11758_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__or2_1
XFILLER_187_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17254_ _17452_/Q _17293_/A2 _17252_/X _17253_/X _17293_/C1 vssd1 vssd1 vccd1 vccd1
+ _17452_/D sky130_fd_sc_hd__o221a_1
X_14466_ _14466_/A _14466_/B vssd1 vssd1 vccd1 vccd1 _14524_/B sky130_fd_sc_hd__and2_2
XFILLER_175_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11678_/A _11678_/B vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__and2_1
XFILLER_174_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _16292_/B _16205_/B vssd1 vssd1 vccd1 vccd1 _16205_/X sky130_fd_sc_hd__or2_4
XFILLER_174_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13417_ _13417_/A _13417_/B _13417_/C vssd1 vssd1 vccd1 vccd1 _13418_/B sky130_fd_sc_hd__or3_1
X_10629_ _10614_/X _10615_/Y _10623_/X _10627_/X vssd1 vssd1 vccd1 vccd1 _10632_/C
+ sky130_fd_sc_hd__a211o_2
X_17185_ input25/X _17362_/A input1/X _17428_/C vssd1 vssd1 vccd1 vccd1 _17185_/X
+ sky130_fd_sc_hd__and4_1
X_14397_ _14316_/A _14332_/X _14395_/Y _14396_/X vssd1 vssd1 vccd1 vccd1 _14466_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _16136_/A _16136_/B _16136_/C vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__and3_1
X_13348_ _17405_/A _13566_/B vssd1 vssd1 vccd1 vccd1 _13349_/B sky130_fd_sc_hd__nand2_4
XFILLER_182_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16067_ _15853_/B _15955_/Y _15960_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _16068_/B
+ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_170_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13279_ _13948_/A _13948_/B _14155_/B _14063_/C vssd1 vssd1 vccd1 vccd1 _13280_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15018_ _11334_/C _14967_/C _14967_/D _14900_/X _14877_/Y vssd1 vssd1 vccd1 vccd1
+ _15018_/X sky130_fd_sc_hd__o32a_2
XFILLER_64_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16969_ _16969_/A _16969_/B vssd1 vssd1 vccd1 vccd1 _16969_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _10067_/A _12770_/D _09382_/C vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__a21oi_1
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09441_ _09441_/A _09441_/B _09441_/C vssd1 vssd1 vccd1 vccd1 _09441_/Y sky130_fd_sc_hd__nand3_2
XFILLER_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09372_ _12166_/A _09509_/B _09209_/C vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__a21oi_2
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_192_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_145_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_99_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_88_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _09709_/A _09709_/B vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__nand2b_2
X_10980_ _11124_/C _10932_/B _10936_/B _10935_/A vssd1 vssd1 vccd1 vccd1 _10987_/A
+ sky130_fd_sc_hd__a31o_4
Xwb_buttons_leds_955 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_955/HI led_enb[8] sky130_fd_sc_hd__conb_1
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09639_ _09640_/A _09638_/Y _10321_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09795_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_43_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _12649_/B _12650_/B vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__nand2b_1
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__nand2_1
X_12581_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12583_/B sky130_fd_sc_hd__xnor2_2
XFILLER_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14320_ _14387_/A _14599_/D _14321_/C vssd1 vssd1 vccd1 vccd1 _14324_/A sky130_fd_sc_hd__a21oi_1
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11532_ _11532_/A _11532_/B _11574_/A vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__nor3b_4
XFILLER_183_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_184_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14251_ _14252_/A _14252_/B _14252_/C vssd1 vssd1 vccd1 vccd1 _14253_/A sky130_fd_sc_hd__a21oi_4
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11463_ _11416_/B _11413_/B _11413_/C vssd1 vssd1 vccd1 vccd1 _11464_/B sky130_fd_sc_hd__o21a_1
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13332_/A _13202_/B _13202_/C vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__and3_4
XFILLER_183_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10414_ _10415_/A _10413_/Y _10970_/A _10745_/D vssd1 vssd1 vccd1 vccd1 _10513_/A
+ sky130_fd_sc_hd__and4bb_2
X_14182_ _14254_/A _14181_/B _14181_/C vssd1 vssd1 vccd1 vccd1 _14184_/C sky130_fd_sc_hd__a21o_1
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_178_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11394_ _11453_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__and2_2
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13133_ _12993_/X _12999_/A _13264_/B _13132_/X vssd1 vssd1 vccd1 vccd1 _13137_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10345_ _10345_/A _10581_/A vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__nor2_2
XFILLER_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_155_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13065_/A _13065_/B _13065_/C vssd1 vssd1 vccd1 vccd1 _13075_/A sky130_fd_sc_hd__a21o_4
XFILLER_155_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10276_ _10276_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__xor2_1
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12015_ _09679_/A _09826_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _12015_/Y sky130_fd_sc_hd__o21bai_4
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16823_ _16897_/A _16823_/B vssd1 vssd1 vccd1 vccd1 _16832_/A sky130_fd_sc_hd__or2_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13966_ _14050_/A _14050_/B _14050_/D _13966_/D vssd1 vssd1 vccd1 vccd1 _13967_/B
+ sky130_fd_sc_hd__and4_1
X_16754_ _16680_/X _16684_/B _16682_/B vssd1 vssd1 vccd1 vccd1 _16764_/B sky130_fd_sc_hd__o21a_1
XFILLER_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15705_ _15705_/A _15705_/B _15705_/C vssd1 vssd1 vccd1 vccd1 _15705_/Y sky130_fd_sc_hd__nand3_1
X_12917_ _13065_/A _12918_/B _12918_/C vssd1 vssd1 vccd1 vccd1 _12919_/A sky130_fd_sc_hd__a21o_1
X_16685_ _16686_/A _16686_/B _16684_/Y vssd1 vssd1 vccd1 vccd1 _16685_/X sky130_fd_sc_hd__o21ba_1
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13897_ _17409_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _13898_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1048 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12848_ _12212_/X _12217_/B _17367_/A vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__mux2_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15636_ _15636_/A vssd1 vssd1 vccd1 vccd1 _17553_/D sky130_fd_sc_hd__clkinv_2
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15567_ _15567_/A _15666_/A vssd1 vssd1 vccd1 vccd1 _15568_/B sky130_fd_sc_hd__nand2_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12779_/A _12779_/B vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__nor2_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14518_ _14518_/A _14518_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14519_/C sky130_fd_sc_hd__nand3_1
X_17306_ _17306_/A1 _17328_/A2 _17305_/X _17380_/C1 vssd1 vssd1 vccd1 vccd1 _17482_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15498_ _15498_/A _15498_/B vssd1 vssd1 vccd1 vccd1 _15499_/B sky130_fd_sc_hd__xor2_4
XFILLER_30_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14449_ _16913_/C _14708_/C vssd1 vssd1 vccd1 vccd1 _14509_/B sky130_fd_sc_hd__nand2_1
X_17237_ _17588_/Q _17288_/A2 _17288_/B1 vssd1 vssd1 vccd1 vccd1 _17237_/X sky130_fd_sc_hd__a21o_1
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ _17167_/A _17167_/B _17167_/C vssd1 vssd1 vccd1 vccd1 _17168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_190_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_66_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16119_ _16112_/B _17162_/A2 _16733_/B1 _17119_/A _16218_/C1 vssd1 vssd1 vccd1 vccd1
+ _16119_/X sky130_fd_sc_hd__a221o_1
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17099_ _17099_/A vssd1 vssd1 vccd1 vccd1 _17099_/Y sky130_fd_sc_hd__inv_2
X_09990_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10004_/C sky130_fd_sc_hd__nand2_2
XFILLER_170_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08943_/A sky130_fd_sc_hd__nor2_4
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08872_ _08874_/A _08874_/B _08873_/C _08873_/D vssd1 vssd1 vccd1 vccd1 _08872_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_97_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09424_ _16809_/A _16758_/A vssd1 vssd1 vccd1 vccd1 _09424_/X sky130_fd_sc_hd__and2_4
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09355_ _09355_/A _09355_/B vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__xnor2_4
XFILLER_166_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09286_ _17081_/B _16990_/A _09285_/X vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__o21ai_4
XFILLER_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10130_ _10128_/B _10251_/B _10128_/A vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__o21ba_2
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__xnor2_2
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _13820_/A _13820_/B vssd1 vssd1 vccd1 vccd1 _13823_/A sky130_fd_sc_hd__xor2_4
XFILLER_56_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _13751_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__xnor2_2
X_10963_ _10963_/A _10963_/B _10963_/C _10963_/D vssd1 vssd1 vccd1 vccd1 _10965_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _12027_/X _12034_/X _12865_/S vssd1 vssd1 vccd1 vccd1 _12702_/X sky130_fd_sc_hd__mux2_1
X_16470_ _16470_/A _16470_/B _16470_/C vssd1 vssd1 vccd1 vccd1 _16563_/B sky130_fd_sc_hd__and3_1
X_13682_ _13582_/A _13584_/B _13582_/B vssd1 vssd1 vccd1 vccd1 _13683_/B sky130_fd_sc_hd__o21ba_1
XFILLER_188_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _10881_/Y _11112_/A _10895_/A _10864_/Y vssd1 vssd1 vccd1 vccd1 _11080_/A
+ sky130_fd_sc_hd__o211ai_4
X_15421_ _15422_/A _15422_/B vssd1 vssd1 vccd1 vccd1 _15507_/A sky130_fd_sc_hd__and2b_2
X_12633_ _12630_/X _12631_/Y _12481_/A _12481_/Y vssd1 vssd1 vccd1 vccd1 _12676_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_188_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15352_ _15352_/A _15352_/B vssd1 vssd1 vccd1 vccd1 _15359_/A sky130_fd_sc_hd__xnor2_4
X_12564_ _17395_/A _12565_/C _12565_/D _17397_/A vssd1 vssd1 vccd1 vccd1 _12566_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_180_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _16965_/C _14545_/C vssd1 vssd1 vccd1 vccd1 _14304_/B sky130_fd_sc_hd__nand2_4
Xwire120 wire120/A vssd1 vssd1 vccd1 vccd1 wire120/X sky130_fd_sc_hd__buf_4
XFILLER_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11515_ _11520_/C _11518_/C _11484_/B _11481_/Y vssd1 vssd1 vccd1 vccd1 _11522_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_102_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15283_ _15283_/A _15283_/B vssd1 vssd1 vccd1 vccd1 _15285_/B sky130_fd_sc_hd__xnor2_4
X_12495_ _12795_/A _12638_/B vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__nand2_1
XFILLER_144_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17022_ _17018_/A _17066_/A _17066_/B _17156_/B vssd1 vssd1 vccd1 vccd1 _17022_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14234_ _14235_/A _14235_/B vssd1 vssd1 vccd1 vccd1 _14315_/A sky130_fd_sc_hd__or2_1
XFILLER_109_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11446_ _11396_/X _11421_/Y _11444_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _11449_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_137_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ _14165_/A _14165_/B vssd1 vssd1 vccd1 vccd1 _14185_/A sky130_fd_sc_hd__xnor2_1
XFILLER_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11377_ _11506_/A _11377_/B _11377_/C _11377_/D vssd1 vssd1 vccd1 vccd1 _11380_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_153_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_996 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ _13117_/A _13117_/B _13117_/C vssd1 vssd1 vccd1 vccd1 _13118_/A sky130_fd_sc_hd__a21o_1
XFILLER_152_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10329_/B _10329_/C vssd1 vssd1 vccd1 vccd1 _10450_/B sky130_fd_sc_hd__and2_1
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14096_ _14200_/B _14096_/B vssd1 vssd1 vccd1 vccd1 _14098_/B sky130_fd_sc_hd__or2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13047_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13049_/C sky130_fd_sc_hd__nand2_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10260_/B _10260_/A vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__nand2b_2
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _13789_/C _16806_/A2 _16805_/X vssd1 vssd1 vccd1 vccd1 _17566_/D sky130_fd_sc_hd__a21oi_1
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14998_ _15100_/A _14998_/B vssd1 vssd1 vccd1 vccd1 _14998_/Y sky130_fd_sc_hd__nand2_1
X_16737_ _16485_/A _16730_/Y _16732_/X _16736_/X vssd1 vssd1 vccd1 vccd1 _16737_/X
+ sky130_fd_sc_hd__a211o_2
X_13949_ _13949_/A _13949_/B vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__nor2_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16668_ _16670_/A _16670_/B _16670_/C vssd1 vssd1 vccd1 vccd1 _16671_/A sky130_fd_sc_hd__a21oi_1
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15619_ _15453_/B _15453_/C _15529_/Y _15449_/Y vssd1 vssd1 vccd1 vccd1 _15620_/B
+ sky130_fd_sc_hd__a211o_1
X_16599_ _16600_/A _16600_/B vssd1 vssd1 vccd1 vccd1 _16601_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09140_ _09106_/A _09108_/B _09106_/B vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__o21ba_4
XFILLER_188_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09071_ _09071_/A _09071_/B _09071_/C vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__nor3_4
XFILLER_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_163_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09973_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__and2_2
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08924_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__and2_2
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_85_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08855_ _17375_/A _12102_/D vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__nand2_1
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08786_ _08787_/B vssd1 vssd1 vccd1 vccd1 _08786_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _09838_/A _09407_/B _09647_/B _09937_/B vssd1 vssd1 vccd1 vccd1 _09410_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09338_ _09338_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09339_/C sky130_fd_sc_hd__xnor2_2
XFILLER_178_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _09269_/A _09269_/B _09275_/B vssd1 vssd1 vccd1 vccd1 _09290_/B sky130_fd_sc_hd__or3_1
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ _11299_/B _11415_/A vssd1 vssd1 vccd1 vccd1 _11711_/B sky130_fd_sc_hd__nand2b_2
X_12280_ _12281_/B _12281_/A vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__and2b_2
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ _11229_/A _11199_/X _11229_/B vssd1 vssd1 vccd1 vccd1 _11231_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11162_ _11162_/A _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__and3_2
XFILLER_136_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_96_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10113_/A _10113_/B _10119_/B vssd1 vssd1 vccd1 vccd1 _10133_/B sky130_fd_sc_hd__or3_4
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15970_ _16084_/B _15970_/B vssd1 vssd1 vccd1 vccd1 _15972_/B sky130_fd_sc_hd__or2_2
X_11093_ _14785_/A _10957_/D _10822_/A _10820_/Y vssd1 vssd1 vccd1 vccd1 _11099_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10044_ _10171_/B _10657_/B _10659_/D _14789_/A vssd1 vssd1 vccd1 vccd1 _10044_/Y
+ sky130_fd_sc_hd__a22oi_2
X_14921_ _14848_/B _14848_/A _15314_/A _15381_/A _14942_/A _14958_/A vssd1 vssd1 vccd1
+ vccd1 _14921_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14852_ _15541_/A _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15624_/B sky130_fd_sc_hd__and3_1
XFILLER_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13803_ _13803_/A _13803_/B vssd1 vssd1 vccd1 vccd1 _13805_/B sky130_fd_sc_hd__xnor2_1
XFILLER_17_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17571_ fanout945/X _17571_/D vssd1 vssd1 vccd1 vccd1 _17571_/Q sky130_fd_sc_hd__dfxtp_1
X_14783_ _15262_/A _15709_/A vssd1 vssd1 vccd1 vccd1 _15707_/B sky130_fd_sc_hd__or2_2
XFILLER_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11995_ _09248_/B _09248_/Y _12197_/A _11994_/X vssd1 vssd1 vccd1 vccd1 _12197_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13734_ _13844_/B _14175_/B _14002_/B _13844_/A vssd1 vssd1 vccd1 vccd1 _13736_/A
+ sky130_fd_sc_hd__a22oi_2
X_16522_ _16522_/A _16522_/B vssd1 vssd1 vccd1 vccd1 _16524_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10946_ _10946_/A _10946_/B _10946_/C vssd1 vssd1 vccd1 vccd1 _10946_/X sky130_fd_sc_hd__and3_4
XFILLER_95_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16453_ _16453_/A _16453_/B vssd1 vssd1 vccd1 vccd1 _16454_/B sky130_fd_sc_hd__xnor2_2
X_13665_ _13665_/A _13778_/A vssd1 vssd1 vccd1 vccd1 _13668_/A sky130_fd_sc_hd__or2_1
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10877_ _10878_/A _10876_/Y _11553_/B _10971_/B vssd1 vssd1 vccd1 vccd1 _11121_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__xnor2_2
X_12616_ _12616_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__or2_2
XFILLER_188_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16384_ _16385_/A _16385_/B vssd1 vssd1 vccd1 vccd1 _16384_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13597_/A _13597_/B vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__and2_2
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15335_ _15337_/A _15337_/B vssd1 vssd1 vccd1 vccd1 _15335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12547_ _11810_/X _11818_/B _17367_/A vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15820_/A _16262_/A _15331_/A vssd1 vssd1 vccd1 vccd1 _15337_/A sky130_fd_sc_hd__or3_4
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12478_ _12478_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _12481_/C sky130_fd_sc_hd__xor2_4
XFILLER_138_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_3 _16478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14217_ _14218_/A _14218_/B _14218_/C vssd1 vssd1 vccd1 vccd1 _14297_/A sky130_fd_sc_hd__o21ai_4
XFILLER_172_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17005_ _16955_/A _16955_/B _16953_/A vssd1 vssd1 vccd1 vccd1 _17007_/B sky130_fd_sc_hd__a21oi_4
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11429_ _11553_/A _11561_/D _15402_/A _11506_/A vssd1 vssd1 vccd1 vccd1 _11430_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15197_ _15821_/A _16226_/C vssd1 vssd1 vccd1 vccd1 _15220_/A sky130_fd_sc_hd__nand2_4
XFILLER_126_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _14148_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14150_/C sky130_fd_sc_hd__xnor2_1
XFILLER_125_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14079_ _14318_/B _14545_/D _14080_/C vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__a21oi_1
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09123_ _12772_/A _17466_/D vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__nand2_4
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09054_ _09055_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__a21o_4
XFILLER_190_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _09956_/A _09956_/B vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__or2_1
XFILLER_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09765_/A _09765_/B _09765_/C vssd1 vssd1 vccd1 vccd1 _09887_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_58_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _17381_/A _12090_/B _08835_/Y _08862_/A vssd1 vssd1 vccd1 vccd1 _08839_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_58_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _09023_/A _09023_/B _12166_/B _12158_/C vssd1 vssd1 vccd1 vccd1 _08773_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _11314_/A _10911_/B _10800_/C vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__and3_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11781_/B vssd1 vssd1 vccd1 vccd1 _11780_/Y sky130_fd_sc_hd__inv_2
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10731_ _10712_/X _10730_/Y _10631_/X _10693_/Y vssd1 vssd1 vccd1 vccd1 _10766_/C
+ sky130_fd_sc_hd__a211o_4
XFILLER_80_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_158_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _13895_/A _14383_/A _13564_/D _13450_/D vssd1 vssd1 vccd1 vccd1 _13569_/A
+ sky130_fd_sc_hd__and4_1
X_10662_ _10662_/A _10662_/B _10662_/C vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__and3_4
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _12401_/A _12401_/B vssd1 vssd1 vccd1 vccd1 _12401_/X sky130_fd_sc_hd__or2_1
X_13381_ _13221_/A _13224_/A _13504_/A _13380_/X vssd1 vssd1 vccd1 vccd1 _13504_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_166_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10593_ _10593_/A _10593_/B vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__nand2_2
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15120_ _15119_/A _15119_/B _15309_/B vssd1 vssd1 vccd1 vccd1 _15120_/X sky130_fd_sc_hd__a21o_1
X_12332_ _12166_/A _12166_/B _12167_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12333_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_154_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15051_/A _16304_/A _15050_/X vssd1 vssd1 vccd1 vccd1 _15051_/X sky130_fd_sc_hd__or3b_1
X_12263_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12265_/C sky130_fd_sc_hd__xnor2_4
XFILLER_108_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ _14326_/A _14002_/B _14002_/C vssd1 vssd1 vccd1 vccd1 _14092_/B sky130_fd_sc_hd__nand3_2
XFILLER_181_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11214_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12194_ _12360_/A _12193_/B _12193_/C vssd1 vssd1 vccd1 vccd1 _12194_/X sky130_fd_sc_hd__a21o_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_966 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_150_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput73 _17477_/Q vssd1 vssd1 vccd1 vccd1 leds[11] sky130_fd_sc_hd__clkbuf_2
X_11145_ _11145_/A _11145_/B _11145_/C vssd1 vssd1 vccd1 vccd1 _11153_/B sky130_fd_sc_hd__and3_4
Xoutput84 _17434_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_49_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput95 _17435_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[1] sky130_fd_sc_hd__clkbuf_2
X_15953_ _15953_/A _15953_/B vssd1 vssd1 vccd1 vccd1 _15954_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11076_ _11059_/A _11059_/B _11059_/C vssd1 vssd1 vccd1 vccd1 _11077_/C sky130_fd_sc_hd__a21oi_4
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14904_ _08731_/A _15147_/A vssd1 vssd1 vccd1 vccd1 _14905_/D sky130_fd_sc_hd__nand2b_1
X_10027_ _10028_/A _10027_/B _10027_/C _10027_/D vssd1 vssd1 vccd1 vccd1 _10028_/B
+ sky130_fd_sc_hd__and4b_4
XFILLER_76_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15884_ _15884_/A _15884_/B vssd1 vssd1 vccd1 vccd1 _15884_/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14835_ _14836_/A _14836_/B _14933_/B vssd1 vssd1 vccd1 vccd1 _15108_/A sky130_fd_sc_hd__and3_4
XTAP_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ fanout946/X _17554_/D vssd1 vssd1 vccd1 vccd1 _17554_/Q sky130_fd_sc_hd__dfxtp_2
X_14766_ _14766_/A _17028_/A vssd1 vssd1 vccd1 vccd1 _17023_/B sky130_fd_sc_hd__or2_2
X_11978_ _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11980_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16505_ _16505_/A _16505_/B vssd1 vssd1 vccd1 vccd1 _16505_/X sky130_fd_sc_hd__or2_1
XFILLER_147_1052 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13717_ _13818_/B _13717_/B vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__and2_2
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ _11057_/A _11057_/B _11057_/C vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__a21o_4
XFILLER_177_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14697_ _14698_/B _14699_/A vssd1 vssd1 vccd1 vccd1 _14729_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17485_ fanout927/X _17485_/D vssd1 vssd1 vccd1 vccd1 _17485_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_108_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16436_ _16436_/A _16436_/B vssd1 vssd1 vccd1 vccd1 _16437_/B sky130_fd_sc_hd__xnor2_4
X_13648_ _13749_/B _13648_/B _13648_/C vssd1 vssd1 vccd1 vccd1 _13648_/X sky130_fd_sc_hd__and3_1
XFILLER_158_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16367_ _16367_/A _16367_/B vssd1 vssd1 vccd1 vccd1 _16369_/A sky130_fd_sc_hd__xor2_4
X_13579_ _13579_/A _13579_/B vssd1 vssd1 vccd1 vccd1 _13597_/A sky130_fd_sc_hd__xnor2_2
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15318_ _14790_/A _16735_/A _12710_/B _15315_/X _15317_/X vssd1 vssd1 vccd1 vccd1
+ _15321_/C sky130_fd_sc_hd__o311a_1
X_16298_ _16298_/A _16391_/B _14777_/A vssd1 vssd1 vccd1 vccd1 _16299_/B sky130_fd_sc_hd__or3b_2
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15249_ _15244_/B _14929_/X _15713_/B1 _14848_/A vssd1 vssd1 vccd1 vccd1 _15249_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_172_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09810_ _09789_/A _09933_/A _09789_/B _09920_/A vssd1 vssd1 vccd1 vccd1 _09811_/B
+ sky130_fd_sc_hd__o31ai_4
Xfanout307 _08731_/A vssd1 vssd1 vccd1 vccd1 _15071_/A sky130_fd_sc_hd__buf_8
Xfanout318 _14290_/A vssd1 vssd1 vccd1 vccd1 _14593_/A sky130_fd_sc_hd__buf_6
XFILLER_119_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout329 _17540_/Q vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__buf_8
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1029 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09741_ _09768_/B _09832_/A _09768_/A vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09672_ _09674_/B _09819_/A _09674_/A vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__o21a_2
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09106_ _09106_/A _09106_/B vssd1 vssd1 vccd1 vccd1 _09108_/A sky130_fd_sc_hd__nor2_1
XFILLER_182_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09037_ _09037_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__xnor2_4
XFILLER_164_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_191_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout830 _17485_/Q vssd1 vssd1 vccd1 vccd1 _12618_/D sky130_fd_sc_hd__buf_12
Xfanout841 _10963_/C vssd1 vssd1 vccd1 vccd1 _10911_/B sky130_fd_sc_hd__buf_12
Xfanout852 _10963_/D vssd1 vssd1 vccd1 vccd1 _14848_/A sky130_fd_sc_hd__buf_6
XFILLER_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout863 _11377_/C vssd1 vssd1 vccd1 vccd1 _15175_/B sky130_fd_sc_hd__clkbuf_16
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout874 _11629_/C vssd1 vssd1 vccd1 vccd1 _15116_/B sky130_fd_sc_hd__clkbuf_8
Xfanout885 _15402_/A vssd1 vssd1 vccd1 vccd1 _15401_/A sky130_fd_sc_hd__buf_6
Xfanout896 _10560_/D vssd1 vssd1 vccd1 vccd1 _17466_/D sky130_fd_sc_hd__buf_8
XFILLER_58_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12950_ _17407_/A _12950_/B _12950_/C vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__nand3_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11901_ _11901_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__nor2_1
XFILLER_73_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12881_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _12882_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _14621_/A _14621_/B _14621_/C vssd1 vssd1 vccd1 vccd1 _14661_/A sky130_fd_sc_hd__a21oi_2
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _11829_/Y _11831_/Y _12390_/S vssd1 vssd1 vccd1 vccd1 _11832_/X sky130_fd_sc_hd__mux2_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14680_/A _14641_/C _14679_/B vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__a21boi_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11750_/A _16794_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10715_/A _10715_/B _10715_/C vssd1 vssd1 vccd1 vccd1 _10714_/X sky130_fd_sc_hd__a21o_4
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13347_/B _13349_/B _13347_/A vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__o21ba_1
X_17270_ _17599_/Q _17270_/A2 _17270_/B1 vssd1 vssd1 vccd1 vccd1 _17270_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _13838_/S _12866_/B _14210_/B _14758_/A vssd1 vssd1 vccd1 vccd1 _14482_/X
+ sky130_fd_sc_hd__o31a_1
X_11694_ _11672_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11694_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13433_ _17423_/A _13434_/C _13434_/D _17425_/A vssd1 vssd1 vccd1 vccd1 _13435_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16221_ _16221_/A _16221_/B _16215_/X vssd1 vssd1 vccd1 vccd1 _16221_/X sky130_fd_sc_hd__or3b_2
X_10645_ _10933_/A _10933_/B _10645_/C _10743_/C vssd1 vssd1 vccd1 vccd1 _10648_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_155_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16152_ _16152_/A _16812_/A vssd1 vssd1 vccd1 vccd1 _16153_/B sky130_fd_sc_hd__nand2_4
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13364_ _13482_/A _13364_/B vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__nor2_2
XFILLER_177_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10576_ _10573_/X _10575_/Y _10463_/B _10471_/X vssd1 vssd1 vccd1 vccd1 _10579_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _12316_/A _12316_/B _12316_/C vssd1 vssd1 vccd1 vccd1 _12526_/A sky130_fd_sc_hd__a21o_4
X_15103_ _15100_/Y _15102_/Y _15130_/S vssd1 vssd1 vccd1 vccd1 _15103_/X sky130_fd_sc_hd__mux2_1
X_16083_ _16084_/A _16084_/B _16082_/X vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__o21ba_1
XFILLER_177_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13295_ _13295_/A _13295_/B _13295_/C vssd1 vssd1 vccd1 vccd1 _13308_/B sky130_fd_sc_hd__nand3_2
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15034_ _15100_/A _15034_/B vssd1 vssd1 vccd1 vccd1 _15034_/Y sky130_fd_sc_hd__nand2_1
X_12246_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__nor2_1
XFILLER_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_170_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ _12177_/A _12177_/B vssd1 vssd1 vccd1 vccd1 _12179_/C sky130_fd_sc_hd__xnor2_2
XFILLER_3_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11128_ _11130_/B _11130_/C _11130_/A vssd1 vssd1 vccd1 vccd1 _11128_/Y sky130_fd_sc_hd__a21oi_4
X_16985_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _17046_/A sky130_fd_sc_hd__and2b_1
XFILLER_84_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15936_ _15937_/A _15937_/B vssd1 vssd1 vccd1 vccd1 _16072_/A sky130_fd_sc_hd__and2_1
XFILLER_37_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11059_ _11059_/A _11059_/B _11059_/C vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__and3_4
XFILLER_114_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_188_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15867_ _15867_/A _15867_/B vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__and2_1
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ fanout940/X _17606_/D vssd1 vssd1 vccd1 vccd1 _17606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14818_ _16576_/B _16577_/A _12869_/C vssd1 vssd1 vccd1 vccd1 _16649_/C sky130_fd_sc_hd__a21o_1
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _15705_/B _15705_/C _15705_/A vssd1 vssd1 vccd1 vccd1 _15798_/Y sky130_fd_sc_hd__a21boi_4
X_17537_ fanout933/X _17537_/D vssd1 vssd1 vccd1 vccd1 _17537_/Q sky130_fd_sc_hd__dfxtp_4
X_14749_ _14750_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__or2_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_177_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17468_ fanout928/X _17468_/D vssd1 vssd1 vccd1 vccd1 _17468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16419_ _16419_/A _16419_/B vssd1 vssd1 vccd1 vccd1 _16420_/A sky130_fd_sc_hd__xnor2_1
X_17399_ _17399_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17399_/X sky130_fd_sc_hd__or2_1
XFILLER_164_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_173_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_156_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_160_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout126 _17198_/X vssd1 vssd1 vccd1 vccd1 _17229_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout137 _15734_/B vssd1 vssd1 vccd1 vccd1 _16315_/C sky130_fd_sc_hd__buf_6
Xfanout148 _14969_/Y vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__buf_2
Xfanout159 _17362_/X vssd1 vssd1 vccd1 vccd1 _17384_/A2 sky130_fd_sc_hd__buf_6
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _09725_/A _09725_/B _09725_/C vssd1 vssd1 vccd1 vccd1 _09724_/X sky130_fd_sc_hd__a21o_4
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09655_ _09655_/A _09784_/A vssd1 vssd1 vccd1 vccd1 _09656_/C sky130_fd_sc_hd__nor2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_41_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09587_/A _09585_/Y _11902_/A _09892_/C vssd1 vssd1 vccd1 vccd1 _09727_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10430_ _10430_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__and2_2
XFILLER_183_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_100_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10361_ _10694_/B _10479_/B _10360_/D _10694_/A vssd1 vssd1 vccd1 vccd1 _10362_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_109_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _12097_/X _12268_/B _11891_/A _11891_/Y vssd1 vssd1 vccd1 vccd1 _12122_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _14769_/A _14770_/A _13866_/D _13229_/B vssd1 vssd1 vccd1 vccd1 _13213_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ _10293_/A _10291_/Y _14788_/A _10899_/D vssd1 vssd1 vccd1 vccd1 _10399_/A
+ sky130_fd_sc_hd__and4bb_2
XFILLER_152_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_151_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ _12031_/A _12031_/B vssd1 vssd1 vccd1 vccd1 _12031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout660 _09654_/D vssd1 vssd1 vccd1 vccd1 _12576_/C sky130_fd_sc_hd__buf_4
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout671 fanout676/X vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__buf_6
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _16770_/A _16770_/B _16770_/C vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__or3_1
Xfanout682 fanout686/X vssd1 vssd1 vccd1 vccd1 _14215_/B sky130_fd_sc_hd__buf_8
X_13982_ _13982_/A _13982_/B vssd1 vssd1 vccd1 vccd1 _13985_/A sky130_fd_sc_hd__xnor2_4
XFILLER_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout693 _16722_/A vssd1 vssd1 vccd1 vccd1 _13566_/B sky130_fd_sc_hd__buf_12
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15721_ _16911_/A _15700_/Y _15720_/X vssd1 vssd1 vccd1 vccd1 _15721_/X sky130_fd_sc_hd__a21o_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12933_ _12933_/A _12933_/B _12933_/C vssd1 vssd1 vccd1 vccd1 _12935_/A sky130_fd_sc_hd__nor3_4
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15652_ _15742_/A _15742_/B vssd1 vssd1 vccd1 vccd1 _15743_/A sky130_fd_sc_hd__nor2_2
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A vssd1 vssd1 vccd1 vccd1 _12864_/Y sky130_fd_sc_hd__inv_2
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14603_/A _14646_/A vssd1 vssd1 vccd1 vccd1 _14606_/A sky130_fd_sc_hd__and2_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11815_ _17363_/A _12597_/B vssd1 vssd1 vccd1 vccd1 _14978_/B sky130_fd_sc_hd__and2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _15584_/A _15584_/B vssd1 vssd1 vccd1 vccd1 _15583_/Y sky130_fd_sc_hd__nand2_2
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12795_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12796_/B sky130_fd_sc_hd__nand2_2
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _12659_/B _17322_/A2 _17321_/X _17322_/C1 vssd1 vssd1 vccd1 vccd1 _17490_/D
+ sky130_fd_sc_hd__o211a_1
X_14534_ _14534_/A _14534_/B vssd1 vssd1 vccd1 vccd1 _14534_/Y sky130_fd_sc_hd__nand2_2
XFILLER_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_42_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11746_ _11758_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _16794_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17253_ _17561_/Q _17292_/B vssd1 vssd1 vccd1 vccd1 _17253_/X sky130_fd_sc_hd__and2_1
X_14465_ _14465_/A _14465_/B vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__nand2_2
XFILLER_159_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11677_ _14791_/A _15008_/B _11681_/A _11658_/D vssd1 vssd1 vccd1 vccd1 _11678_/B
+ sky130_fd_sc_hd__a22o_1
X_16204_ _16098_/A _16101_/Y _16203_/B _15523_/A vssd1 vssd1 vccd1 vccd1 _16205_/B
+ sky130_fd_sc_hd__a31o_1
X_13416_ _13417_/A _13417_/B _13417_/C vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__o21ai_4
XFILLER_128_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10628_ _10623_/X _10627_/X _10614_/X _10615_/Y vssd1 vssd1 vccd1 vccd1 _10632_/B
+ sky130_fd_sc_hd__o211ai_4
X_14396_ _14396_/A _14396_/B vssd1 vssd1 vccd1 vccd1 _14396_/X sky130_fd_sc_hd__and2_1
X_17184_ input25/X _17428_/C vssd1 vssd1 vccd1 vccd1 _17362_/B sky130_fd_sc_hd__nand2_2
XFILLER_10_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16135_ _16315_/C _16030_/B _16234_/C vssd1 vssd1 vccd1 vccd1 _16137_/A sky130_fd_sc_hd__o21a_1
X_13347_ _13347_/A _13347_/B vssd1 vssd1 vccd1 vccd1 _13349_/A sky130_fd_sc_hd__nor2_2
XFILLER_154_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10559_ _10559_/A _10559_/B vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ _16066_/A _16066_/B vssd1 vssd1 vccd1 vccd1 _16068_/A sky130_fd_sc_hd__xnor2_4
X_13278_ _13948_/B _14155_/B _14063_/C _13948_/A vssd1 vssd1 vccd1 vccd1 _13280_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_64_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12229_ _13627_/S _16011_/B _12229_/C vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__or3_4
X_15017_ _14977_/X _15014_/Y _15016_/Y _16977_/A _11675_/B vssd1 vssd1 vccd1 vccd1
+ _17544_/D sky130_fd_sc_hd__o32a_1
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16968_ _16863_/A _16863_/B _16916_/A _16967_/X vssd1 vssd1 vccd1 vccd1 _16969_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15919_ _16025_/A _15820_/C _15917_/Y _15916_/X vssd1 vssd1 vccd1 vccd1 _15921_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16899_ _16829_/A _16828_/A _16828_/B _16830_/B _16830_/A vssd1 vssd1 vccd1 vccd1
+ _16900_/C sky130_fd_sc_hd__a32o_2
X_09440_ _09441_/A _09441_/B _09441_/C vssd1 vssd1 vccd1 vccd1 _09440_/X sky130_fd_sc_hd__a21o_4
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_80_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09371_ _12800_/A _09555_/C vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__nand2_2
XFILLER_80_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_159_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_181_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_146_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09707_ _16989_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09709_/B sky130_fd_sc_hd__xnor2_4
Xwb_buttons_leds_956 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_956/HI led_enb[9] sky130_fd_sc_hd__conb_1
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09638_ _09637_/B _11920_/D _09944_/D _09942_/A vssd1 vssd1 vccd1 vccd1 _09638_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _16933_/A _16982_/B vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__nand2_2
XFILLER_169_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11600_ _11558_/B _11600_/B vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__and2b_2
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12761_/A sky130_fd_sc_hd__and2b_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ _11496_/B _11493_/B _11493_/C vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__a21oi_4
XFILLER_184_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14250_ _14330_/B _14250_/B vssd1 vssd1 vccd1 vccd1 _14252_/C sky130_fd_sc_hd__nand2_2
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ _11703_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11465_/A sky130_fd_sc_hd__or2_4
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_183_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _13332_/A _13202_/B _13202_/C vssd1 vssd1 vccd1 vccd1 _13201_/Y sky130_fd_sc_hd__a21oi_4
X_10413_ _10971_/A _10412_/C _10640_/D _10525_/A vssd1 vssd1 vccd1 vccd1 _10413_/Y
+ sky130_fd_sc_hd__a22oi_2
X_14181_ _14254_/A _14181_/B _14181_/C vssd1 vssd1 vccd1 vccd1 _14273_/B sky130_fd_sc_hd__nand3_2
XFILLER_171_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11393_ _11393_/A _11393_/B _11393_/C vssd1 vssd1 vccd1 vccd1 _11394_/B sky130_fd_sc_hd__or3_1
XFILLER_152_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _13264_/A _13130_/Y _12956_/A _12960_/A vssd1 vssd1 vccd1 vccd1 _13132_/X
+ sky130_fd_sc_hd__o211a_1
X_10344_ _10070_/A _10072_/Y _10345_/A _10343_/Y vssd1 vssd1 vccd1 vccd1 _10581_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_3_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _13063_/A _13063_/B vssd1 vssd1 vccd1 vccd1 _13065_/C sky130_fd_sc_hd__nand2_2
XFILLER_152_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10275_ _10276_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__and2_2
XFILLER_151_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12014_ _12375_/A _12014_/B vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__nor2_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_24_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16822_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16823_/B sky130_fd_sc_hd__and2_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout490 _11902_/A vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__buf_6
XFILLER_47_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16753_ _16753_/A _16835_/A vssd1 vssd1 vccd1 vccd1 _16767_/A sky130_fd_sc_hd__or2_1
XFILLER_24_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13965_ _14213_/B _14050_/D _13866_/C _14213_/A vssd1 vssd1 vccd1 vccd1 _13967_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_19_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15704_ _15620_/A _15618_/B _15620_/B _15616_/Y vssd1 vssd1 vccd1 vccd1 _15705_/C
+ sky130_fd_sc_hd__a31o_2
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12916_ _13072_/B _12916_/B vssd1 vssd1 vccd1 vccd1 _12918_/C sky130_fd_sc_hd__nor2_2
XFILLER_185_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16684_ _16684_/A _16684_/B vssd1 vssd1 vccd1 vccd1 _16684_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_74_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13896_ _13896_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _13898_/A sky130_fd_sc_hd__nor2_2
XFILLER_46_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _15617_/A _16218_/C1 _15615_/X _15634_/Y vssd1 vssd1 vccd1 vccd1 _15636_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12847_/A _12847_/B vssd1 vssd1 vccd1 vccd1 _12847_/X sky130_fd_sc_hd__and2_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15566_ _15932_/A _15752_/B vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__nor2_4
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12778_/A _12778_/B _12778_/C vssd1 vssd1 vccd1 vccd1 _12779_/B sky130_fd_sc_hd__and3_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17305_ input62/X _17327_/B _17327_/C vssd1 vssd1 vccd1 vccd1 _17305_/X sky130_fd_sc_hd__or3_1
X_14517_ _14519_/B vssd1 vssd1 vccd1 vccd1 _14517_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_30_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _11731_/B _11729_/B _11729_/C vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__nor3_4
XFILLER_187_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_174_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15497_ _15662_/A _15497_/B vssd1 vssd1 vccd1 vccd1 _15498_/B sky130_fd_sc_hd__nand2_2
XFILLER_147_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _17446_/Q _17290_/A2 _17234_/X _17235_/X _17290_/C1 vssd1 vssd1 vccd1 vccd1
+ _17446_/D sky130_fd_sc_hd__o221a_1
X_14448_ _13895_/B _14554_/B _14708_/D _16913_/C vssd1 vssd1 vccd1 vccd1 _14451_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_30_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17167_ _17167_/A _17167_/B _17167_/C vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__and3_1
X_14379_ _14446_/A _14379_/B vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16118_ _15175_/A _16116_/X _16117_/X _15808_/A vssd1 vssd1 vccd1 vccd1 _16122_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17098_ _17421_/A _17134_/C _14867_/A vssd1 vssd1 vccd1 vccd1 _17099_/A sky130_fd_sc_hd__a21boi_2
XFILLER_66_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16049_ _15927_/B _15941_/B _15925_/Y vssd1 vssd1 vccd1 vccd1 _16051_/B sky130_fd_sc_hd__a21oi_2
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08940_ _17373_/A _11930_/B _12270_/D _12102_/D vssd1 vssd1 vccd1 vccd1 _08941_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_142_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08871_ _08868_/X _08869_/Y _08844_/X _08908_/A vssd1 vssd1 vccd1 vccd1 _08873_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__xnor2_4
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09354_ _09354_/A _09354_/B _09355_/B vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__or3_4
XFILLER_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_127_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09285_ _12256_/B _12638_/B _12637_/C _12256_/A vssd1 vssd1 vccd1 vccd1 _09285_/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_60_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_109_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10060_ _10086_/A vssd1 vssd1 vccd1 vccd1 _10060_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_102_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13750_ _13749_/A _13749_/B _13751_/A vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__a21o_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10962_ _10962_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__nand2_4
XFILLER_84_992 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12701_ _13628_/B vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13681_ _13681_/A _13681_/B vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10893_ _10893_/A _10893_/B _10893_/C vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__and3_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15420_ _15336_/Y _15346_/B _15335_/Y vssd1 vssd1 vccd1 vccd1 _15422_/B sky130_fd_sc_hd__a21o_2
XFILLER_54_1000 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ _12481_/A _12481_/Y _12630_/X _12631_/Y vssd1 vssd1 vccd1 vccd1 _12676_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_31_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12563_ _12563_/A _12730_/A vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__and2_2
X_15351_ _15352_/A _15352_/B vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__or2_2
XFILLER_157_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_180_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14302_ _14302_/A _14302_/B vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__nor2_2
XFILLER_184_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11514_ _11514_/A _11558_/A _11514_/C vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__or3_4
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12494_ _12494_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__nor2_1
X_15282_ _15283_/A _15283_/B vssd1 vssd1 vccd1 vccd1 _15355_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17021_ _17018_/A _17066_/A _17066_/B vssd1 vssd1 vccd1 vccd1 _17021_/Y sky130_fd_sc_hd__a21oi_1
X_14233_ _14159_/B _14161_/B _14159_/A vssd1 vssd1 vccd1 vccd1 _14235_/B sky130_fd_sc_hd__o21ba_1
X_11445_ _11444_/A _11444_/Y _11396_/X _11421_/Y vssd1 vssd1 vccd1 vccd1 _11453_/B
+ sky130_fd_sc_hd__a211o_4
X_14164_ _14165_/A _14165_/B vssd1 vssd1 vccd1 vccd1 _14164_/X sky130_fd_sc_hd__and2b_1
XFILLER_164_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ _11376_/A _11376_/B _11376_/C vssd1 vssd1 vccd1 vccd1 _11395_/B sky130_fd_sc_hd__nand3_4
XFILLER_180_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10327_ _10559_/A _10360_/D _10326_/C vssd1 vssd1 vccd1 vccd1 _10329_/C sky130_fd_sc_hd__a21o_1
X_13115_ _13248_/B _13115_/B vssd1 vssd1 vccd1 vccd1 _13117_/C sky130_fd_sc_hd__or2_1
X_14095_ _14254_/A _14175_/B _14094_/C vssd1 vssd1 vccd1 vccd1 _14096_/B sky130_fd_sc_hd__a21oi_1
XFILLER_152_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13046_/A _13046_/B _13046_/C vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__nand3_4
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _10372_/A _10257_/B _10257_/A vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__o21ba_2
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10189_ _10207_/A _10161_/X _10188_/A _10188_/Y vssd1 vssd1 vccd1 vccd1 _10192_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16805_ _17063_/A _16787_/Y _16793_/X _16804_/X vssd1 vssd1 vccd1 vccd1 _16805_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14997_ _09712_/B _10791_/C _10036_/D _09892_/D _10542_/A _14982_/A vssd1 vssd1 vccd1
+ vccd1 _14999_/B sky130_fd_sc_hd__mux4_1
XFILLER_93_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16736_ _14925_/Y _15313_/Y _16734_/X _16735_/Y vssd1 vssd1 vccd1 vccd1 _16736_/X
+ sky130_fd_sc_hd__a211o_1
X_13948_ _13948_/A _13948_/B _13948_/C _13948_/D vssd1 vssd1 vccd1 vccd1 _13949_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16667_ _16667_/A _16814_/A _16813_/B _16938_/D vssd1 vssd1 vccd1 vccd1 _16670_/C
+ sky130_fd_sc_hd__or4_2
X_13879_ _14226_/A _14213_/C vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__nand2_4
X_15618_ _15616_/Y _15618_/B vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__nand2b_1
X_16598_ _16507_/A _16507_/B _16505_/X vssd1 vssd1 vccd1 vccd1 _16600_/B sky130_fd_sc_hd__a21boi_2
XFILLER_188_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15549_ _15816_/A _16041_/A vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__nor2_4
XFILLER_187_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09070_ _09051_/A _09051_/B _09051_/C vssd1 vssd1 vccd1 vccd1 _09071_/C sky130_fd_sc_hd__a21oi_4
XFILLER_148_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _17582_/Q _17231_/A2 _17231_/B1 vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__a21o_1
XFILLER_175_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _09960_/A _09960_/C _09960_/B vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_89_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08923_ _08923_/A _08923_/B vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08854_ _08854_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _08856_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08785_ _12088_/B _11870_/B _11867_/C _12088_/A vssd1 vssd1 vccd1 vccd1 _08787_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_168_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_77_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09406_ _09411_/A _09411_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__nor2_2
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09337_ _09334_/A _09335_/Y _09344_/A _09316_/X vssd1 vssd1 vccd1 vccd1 _09344_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09268_ _09268_/A _09411_/A vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__nor2_2
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_154_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _12166_/A _09555_/C _09198_/C vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__a21o_1
XFILLER_101_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11230_ _11229_/Y _16387_/A vssd1 vssd1 vccd1 vccd1 _11717_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_84_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_106_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11161_ _11162_/A _11162_/B _11162_/C vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__a21oi_4
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10112_ _10112_/A _10234_/A vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__nor2_4
XFILLER_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__xnor2_2
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ _14789_/A _10171_/B _10657_/B _10659_/D vssd1 vssd1 vccd1 vccd1 _10162_/A
+ sky130_fd_sc_hd__and4_2
X_14920_ _10560_/D _10321_/C _17302_/A1 _11629_/C _14942_/A _14958_/A vssd1 vssd1
+ vccd1 vccd1 _14920_/X sky130_fd_sc_hd__mux4_1
XFILLER_75_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14851_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15541_/B sky130_fd_sc_hd__and2_1
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_63_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13802_ _14008_/A _13903_/B vssd1 vssd1 vccd1 vccd1 _13803_/B sky130_fd_sc_hd__nand2_1
X_17570_ fanout940/X _17570_/D vssd1 vssd1 vccd1 vccd1 _17570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14782_ _16136_/A _15811_/A vssd1 vssd1 vccd1 vccd1 _15801_/B sky130_fd_sc_hd__or2_1
X_11994_ _12155_/B _11993_/C _11993_/A vssd1 vssd1 vccd1 vccd1 _11994_/X sky130_fd_sc_hd__o21a_2
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16521_ _16522_/A _16522_/B vssd1 vssd1 vccd1 vccd1 _16625_/B sky130_fd_sc_hd__and2_1
X_13733_ _14756_/A1 _13731_/Y _13828_/B _13630_/Y vssd1 vssd1 vccd1 vccd1 _17589_/D
+ sky130_fd_sc_hd__a31o_1
X_10945_ _10953_/A _10945_/B vssd1 vssd1 vccd1 vccd1 _10946_/C sky130_fd_sc_hd__and2_2
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_72_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ _16453_/B _16453_/A vssd1 vssd1 vccd1 vccd1 _16452_/Y sky130_fd_sc_hd__nand2b_1
X_13664_ _14050_/A _14050_/B _13764_/D _13664_/D vssd1 vssd1 vccd1 vccd1 _13778_/A
+ sky130_fd_sc_hd__and4_1
X_10876_ _11122_/B _11391_/B _11480_/C _11266_/A vssd1 vssd1 vccd1 vccd1 _10876_/Y
+ sky130_fd_sc_hd__a22oi_2
X_15403_ _16127_/A _16533_/A _15484_/A vssd1 vssd1 vccd1 vccd1 _15403_/X sky130_fd_sc_hd__and3_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12474_/A _12474_/B _12472_/Y vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__a21bo_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _16292_/B _16562_/B _16562_/C vssd1 vssd1 vccd1 vccd1 _16385_/B sky130_fd_sc_hd__o21a_2
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _13595_/A _13595_/B vssd1 vssd1 vccd1 vccd1 _13597_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15334_ _15334_/A _15334_/B vssd1 vssd1 vccd1 vccd1 _15337_/B sky130_fd_sc_hd__xor2_4
X_12546_ _12845_/S _12546_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12548_/B sky130_fd_sc_hd__and3_2
XFILLER_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15265_ _14899_/X _14968_/X _16446_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _15331_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12477_ _12477_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__nor2_4
X_17004_ _17090_/A _17004_/B vssd1 vssd1 vccd1 vccd1 _17007_/A sky130_fd_sc_hd__nand2_4
XANTENNA_4 _16795_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14216_/A _14216_/B vssd1 vssd1 vccd1 vccd1 _14218_/C sky130_fd_sc_hd__xnor2_2
XFILLER_160_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ _11553_/B _11563_/D vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__nand2_2
XFILLER_172_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15196_ _15175_/B _16008_/C1 _15195_/X vssd1 vssd1 vccd1 vccd1 _17547_/D sky130_fd_sc_hd__a21oi_4
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14147_ _14148_/A _14148_/B vssd1 vssd1 vccd1 vccd1 _14221_/B sky130_fd_sc_hd__and2b_1
X_11359_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11413_/B sky130_fd_sc_hd__and2_2
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_193_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14078_ _14188_/A _14078_/B vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13029_ _13029_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__xnor2_4
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_67_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16719_ _16715_/Y _16717_/Y _16718_/Y vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_23_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_124_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ _09122_/A _09122_/B vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__nor2_4
XFILLER_41_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _09053_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _09055_/C sky130_fd_sc_hd__or2_2
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_171_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ _09956_/A _09956_/B vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__nand2_2
XFILLER_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08906_ _08905_/A _09051_/A _08832_/Y _08875_/X vssd1 vssd1 vccd1 vccd1 _08929_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09914_/B _10029_/A _09914_/A vssd1 vssd1 vccd1 vccd1 _09915_/A sky130_fd_sc_hd__o21a_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08835_/Y _08862_/A _17381_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _08862_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08768_ _08768_/A _08768_/B vssd1 vssd1 vccd1 vccd1 _08780_/A sky130_fd_sc_hd__nor2_2
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10730_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _10730_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_81_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ _10661_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10662_/C sky130_fd_sc_hd__xnor2_4
XFILLER_167_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12400_ _13390_/S _12400_/B vssd1 vssd1 vccd1 vccd1 _12401_/B sky130_fd_sc_hd__or2_2
X_13380_ _13500_/B _13378_/X _13252_/Y _13256_/A vssd1 vssd1 vccd1 vccd1 _13380_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_178_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10592_ _10592_/A vssd1 vssd1 vccd1 vccd1 _10593_/B sky130_fd_sc_hd__inv_2
XFILLER_16_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12333_/A vssd1 vssd1 vccd1 vccd1 _12331_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__nand2b_2
X_15050_ _14796_/A _14796_/B _14796_/C _14796_/D vssd1 vssd1 vccd1 vccd1 _15050_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14001_ _14001_/A _14001_/B vssd1 vssd1 vccd1 vccd1 _14002_/C sky130_fd_sc_hd__xor2_2
X_11213_ _11181_/A _11181_/B _11182_/Y vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__a21o_4
X_12193_ _12360_/A _12193_/B _12193_/C vssd1 vssd1 vccd1 vccd1 _12360_/B sky130_fd_sc_hd__nand3_4
XFILLER_107_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11144_ _11144_/A _11237_/A vssd1 vssd1 vccd1 vccd1 _11145_/C sky130_fd_sc_hd__nand2_2
XFILLER_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_123_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput74 _17467_/Q vssd1 vssd1 vccd1 vccd1 leds[1] sky130_fd_sc_hd__clkbuf_2
Xoutput85 _17444_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[10] sky130_fd_sc_hd__clkbuf_2
Xoutput96 _17454_/Q vssd1 vssd1 vccd1 vccd1 o_wb_data[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_49_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15952_ _15953_/A _15953_/B vssd1 vssd1 vccd1 vccd1 _15954_/A sky130_fd_sc_hd__or2_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ _11075_/A _11075_/B _11075_/C vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__or3_4
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14903_ _14879_/Y _15205_/A _14900_/X _15270_/A _14877_/Y vssd1 vssd1 vccd1 vccd1
+ _14903_/X sky130_fd_sc_hd__a2111o_2
X_10026_ _09865_/B _09975_/X _09991_/Y _10005_/X vssd1 vssd1 vccd1 vccd1 _10027_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_49_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15883_ _15883_/A _15883_/B _15881_/Y vssd1 vssd1 vccd1 vccd1 _15884_/B sky130_fd_sc_hd__or3b_2
X_14834_ _17477_/D _17476_/D vssd1 vssd1 vccd1 vccd1 _14938_/B sky130_fd_sc_hd__nand2b_2
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17553_ fanout935/X _17553_/D vssd1 vssd1 vccd1 vccd1 _17553_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14765_ _14765_/A _17065_/A vssd1 vssd1 vccd1 vccd1 _14765_/X sky130_fd_sc_hd__or2_1
XTAP_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _12174_/A _12174_/B _12174_/D _12129_/B vssd1 vssd1 vccd1 vccd1 _11978_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16504_ _16503_/Y _16504_/B vssd1 vssd1 vccd1 vccd1 _16504_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_186_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13716_ _13818_/A _13714_/Y _13601_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _13717_/B
+ sky130_fd_sc_hd__a211o_1
X_10928_ _11074_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _11057_/C sky130_fd_sc_hd__xnor2_4
X_17484_ fanout927/X _17484_/D vssd1 vssd1 vccd1 vccd1 _17484_/Q sky130_fd_sc_hd__dfxtp_4
X_14696_ _14698_/A _14699_/A vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16435_ _16436_/B _16436_/A vssd1 vssd1 vccd1 vccd1 _16435_/X sky130_fd_sc_hd__and2b_1
XFILLER_60_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13647_ _13529_/B _13535_/B _13527_/X vssd1 vssd1 vccd1 vccd1 _13648_/C sky130_fd_sc_hd__a21o_1
X_10859_ _10859_/A _10859_/B _10859_/C vssd1 vssd1 vccd1 vccd1 _10861_/B sky130_fd_sc_hd__nand3_2
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16367_/A _16367_/B vssd1 vssd1 vccd1 vccd1 _16462_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _14254_/A _16859_/A vssd1 vssd1 vccd1 vccd1 _13579_/B sky130_fd_sc_hd__nand2_2
XFILLER_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15317_ _11100_/A _14931_/X _15316_/X _16977_/A vssd1 vssd1 vccd1 vccd1 _15317_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _12528_/A _12528_/B _12528_/C vssd1 vssd1 vccd1 vccd1 _12530_/B sky130_fd_sc_hd__o21a_1
X_16297_ _14777_/A _16209_/B _16298_/A vssd1 vssd1 vccd1 vccd1 _16394_/A sky130_fd_sc_hd__a21bo_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15248_ _15314_/B _15248_/B _15248_/C vssd1 vssd1 vccd1 vccd1 _15257_/B sky130_fd_sc_hd__and3b_1
XFILLER_172_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_912 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_132_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15179_ _14950_/X _14955_/X _15312_/S vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout308 _08731_/A vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__buf_2
Xfanout319 _14738_/A vssd1 vssd1 vccd1 vccd1 _14290_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09740_/A _09740_/B _09740_/C vssd1 vssd1 vccd1 vccd1 _09832_/A sky130_fd_sc_hd__and3_1
XFILLER_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
.ends

