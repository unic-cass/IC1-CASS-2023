magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< obsli1 >>
rect 0 2272 11146 2338
rect 0 66 28 2244
rect 56 94 84 2272
rect 112 66 140 2244
rect 168 94 196 2272
rect 224 66 252 2244
rect 280 94 308 2272
rect 336 66 364 2244
rect 392 94 420 2272
rect 448 66 476 2244
rect 504 94 532 2272
rect 560 66 588 2244
rect 616 94 644 2272
rect 672 66 700 2244
rect 728 94 756 2272
rect 784 66 812 2244
rect 840 94 868 2272
rect 896 66 924 2244
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 1064 94 1092 2272
rect 1120 66 1148 2244
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1288 94 1316 2272
rect 1344 66 1372 2244
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1512 94 1540 2272
rect 1568 66 1596 2244
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1736 94 1764 2272
rect 1792 66 1820 2244
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1960 94 1988 2272
rect 2016 66 2044 2244
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2184 94 2212 2272
rect 2240 66 2268 2244
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2408 94 2436 2272
rect 2464 66 2492 2244
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2632 94 2660 2272
rect 2688 66 2716 2244
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2856 94 2884 2272
rect 2912 66 2940 2244
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 3080 94 3108 2272
rect 3136 66 3164 2244
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3304 94 3332 2272
rect 3360 66 3388 2244
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3528 94 3556 2272
rect 3584 66 3612 2244
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3752 94 3780 2272
rect 3808 66 3836 2244
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3976 94 4004 2272
rect 4032 66 4060 2244
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4200 94 4228 2272
rect 4256 66 4284 2244
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4424 94 4452 2272
rect 4480 66 4508 2244
rect 4536 94 4564 2272
rect 4592 66 4620 2244
rect 4648 94 4676 2272
rect 4704 66 4732 2244
rect 4760 94 4788 2272
rect 4816 66 4844 2244
rect 4872 94 4900 2272
rect 4928 66 4956 2244
rect 4984 94 5012 2272
rect 5040 66 5068 2244
rect 5096 94 5124 2272
rect 5152 66 5180 2244
rect 5208 94 5236 2272
rect 5264 66 5292 2244
rect 5320 94 5348 2272
rect 5376 66 5404 2244
rect 5432 94 5460 2272
rect 5488 66 5516 2244
rect 5544 94 5572 2272
rect 5600 66 5628 2244
rect 5656 94 5684 2272
rect 5712 66 5740 2244
rect 5768 94 5796 2272
rect 5824 66 5852 2244
rect 5880 94 5908 2272
rect 5936 66 5964 2244
rect 5992 94 6020 2272
rect 6048 66 6076 2244
rect 6104 94 6132 2272
rect 6160 66 6188 2244
rect 6216 94 6244 2272
rect 6272 66 6300 2244
rect 6328 94 6356 2272
rect 6384 66 6412 2244
rect 6440 94 6468 2272
rect 6496 66 6524 2244
rect 6552 94 6580 2272
rect 6608 66 6636 2244
rect 6664 94 6692 2272
rect 6720 66 6748 2244
rect 6776 94 6804 2272
rect 6832 66 6860 2244
rect 6888 94 6916 2272
rect 6944 66 6972 2244
rect 7000 94 7028 2272
rect 7056 66 7084 2244
rect 7112 94 7140 2272
rect 7168 66 7196 2244
rect 7224 94 7252 2272
rect 7280 66 7308 2244
rect 7336 94 7364 2272
rect 7392 66 7420 2244
rect 7448 94 7476 2272
rect 7504 66 7532 2244
rect 7560 94 7588 2272
rect 7616 66 7644 2244
rect 7672 94 7700 2272
rect 7728 66 7756 2244
rect 7784 94 7812 2272
rect 7840 66 7868 2244
rect 7896 94 7924 2272
rect 7952 66 7980 2244
rect 8008 94 8036 2272
rect 8064 66 8092 2244
rect 8120 94 8148 2272
rect 8176 66 8204 2244
rect 8232 94 8260 2272
rect 8288 66 8316 2244
rect 8344 94 8372 2272
rect 8400 66 8428 2244
rect 8456 94 8484 2272
rect 8512 66 8540 2244
rect 8568 94 8596 2272
rect 8624 66 8652 2244
rect 8680 94 8708 2272
rect 8736 66 8764 2244
rect 8792 94 8820 2272
rect 8848 66 8876 2244
rect 8904 94 8932 2272
rect 8960 66 8988 2244
rect 9016 94 9044 2272
rect 9072 66 9100 2244
rect 9128 94 9156 2272
rect 9184 66 9212 2244
rect 9240 94 9268 2272
rect 9296 66 9324 2244
rect 9352 94 9380 2272
rect 9408 66 9436 2244
rect 9464 94 9492 2272
rect 9520 66 9548 2244
rect 9576 94 9604 2272
rect 9632 66 9660 2244
rect 9688 94 9716 2272
rect 9744 66 9772 2244
rect 9800 94 9828 2272
rect 9856 66 9884 2244
rect 9912 94 9940 2272
rect 9968 66 9996 2244
rect 10024 94 10052 2272
rect 10080 66 10108 2244
rect 10136 94 10164 2272
rect 10192 66 10220 2244
rect 10248 94 10276 2272
rect 10304 66 10332 2244
rect 10360 94 10388 2272
rect 10416 66 10444 2244
rect 10472 94 10500 2272
rect 10528 66 10556 2244
rect 10584 94 10612 2272
rect 10640 66 10668 2244
rect 10696 94 10724 2272
rect 10752 66 10780 2244
rect 10808 94 10836 2272
rect 10864 66 10892 2244
rect 10920 94 10948 2272
rect 10976 66 11004 2244
rect 11032 94 11060 2272
rect 11088 66 11146 2244
rect 0 0 11146 66
<< obsm1 >>
rect 0 2272 11146 2338
rect 0 94 28 2272
rect 56 66 84 2244
rect 112 94 140 2272
rect 168 66 196 2244
rect 224 94 252 2272
rect 280 66 308 2244
rect 336 94 364 2272
rect 392 66 420 2244
rect 448 94 476 2272
rect 504 66 532 2244
rect 560 94 588 2272
rect 616 66 644 2244
rect 672 94 700 2272
rect 728 66 756 2244
rect 784 94 812 2272
rect 840 66 868 2244
rect 896 94 924 2272
rect 952 66 980 2244
rect 1008 94 1036 2272
rect 1064 66 1092 2244
rect 1120 94 1148 2272
rect 1176 66 1204 2244
rect 1232 94 1260 2272
rect 1288 66 1316 2244
rect 1344 94 1372 2272
rect 1400 66 1428 2244
rect 1456 94 1484 2272
rect 1512 66 1540 2244
rect 1568 94 1596 2272
rect 1624 66 1652 2244
rect 1680 94 1708 2272
rect 1736 66 1764 2244
rect 1792 94 1820 2272
rect 1848 66 1876 2244
rect 1904 94 1932 2272
rect 1960 66 1988 2244
rect 2016 94 2044 2272
rect 2072 66 2100 2244
rect 2128 94 2156 2272
rect 2184 66 2212 2244
rect 2240 94 2268 2272
rect 2296 66 2324 2244
rect 2352 94 2380 2272
rect 2408 66 2436 2244
rect 2464 94 2492 2272
rect 2520 66 2548 2244
rect 2576 94 2604 2272
rect 2632 66 2660 2244
rect 2688 94 2716 2272
rect 2744 66 2772 2244
rect 2800 94 2828 2272
rect 2856 66 2884 2244
rect 2912 94 2940 2272
rect 2968 66 2996 2244
rect 3024 94 3052 2272
rect 3080 66 3108 2244
rect 3136 94 3164 2272
rect 3192 66 3220 2244
rect 3248 94 3276 2272
rect 3304 66 3332 2244
rect 3360 94 3388 2272
rect 3416 66 3444 2244
rect 3472 94 3500 2272
rect 3528 66 3556 2244
rect 3584 94 3612 2272
rect 3640 66 3668 2244
rect 3696 94 3724 2272
rect 3752 66 3780 2244
rect 3808 94 3836 2272
rect 3864 66 3892 2244
rect 3920 94 3948 2272
rect 3976 66 4004 2244
rect 4032 94 4060 2272
rect 4088 66 4116 2244
rect 4144 94 4172 2272
rect 4200 66 4228 2244
rect 4256 94 4284 2272
rect 4312 66 4340 2244
rect 4368 94 4396 2272
rect 4424 66 4452 2244
rect 4480 94 4508 2272
rect 4536 66 4564 2244
rect 4592 94 4620 2272
rect 4648 66 4676 2244
rect 4704 94 4732 2272
rect 4760 66 4788 2244
rect 4816 94 4844 2272
rect 4872 66 4900 2244
rect 4928 94 4956 2272
rect 4984 66 5012 2244
rect 5040 94 5068 2272
rect 5096 66 5124 2244
rect 5152 94 5180 2272
rect 5208 66 5236 2244
rect 5264 94 5292 2272
rect 5320 66 5348 2244
rect 5376 94 5404 2272
rect 5432 66 5460 2244
rect 5488 94 5516 2272
rect 5544 66 5572 2244
rect 5600 94 5628 2272
rect 5656 66 5684 2244
rect 5712 94 5740 2272
rect 5768 66 5796 2244
rect 5824 94 5852 2272
rect 5880 66 5908 2244
rect 5936 94 5964 2272
rect 5992 66 6020 2244
rect 6048 94 6076 2272
rect 6104 66 6132 2244
rect 6160 94 6188 2272
rect 6216 66 6244 2244
rect 6272 94 6300 2272
rect 6328 66 6356 2244
rect 6384 94 6412 2272
rect 6440 66 6468 2244
rect 6496 94 6524 2272
rect 6552 66 6580 2244
rect 6608 94 6636 2272
rect 6664 66 6692 2244
rect 6720 94 6748 2272
rect 6776 66 6804 2244
rect 6832 94 6860 2272
rect 6888 66 6916 2244
rect 6944 94 6972 2272
rect 7000 66 7028 2244
rect 7056 94 7084 2272
rect 7112 66 7140 2244
rect 7168 94 7196 2272
rect 7224 66 7252 2244
rect 7280 94 7308 2272
rect 7336 66 7364 2244
rect 7392 94 7420 2272
rect 7448 66 7476 2244
rect 7504 94 7532 2272
rect 7560 66 7588 2244
rect 7616 94 7644 2272
rect 7672 66 7700 2244
rect 7728 94 7756 2272
rect 7784 66 7812 2244
rect 7840 94 7868 2272
rect 7896 66 7924 2244
rect 7952 94 7980 2272
rect 8008 66 8036 2244
rect 8064 94 8092 2272
rect 8120 66 8148 2244
rect 8176 94 8204 2272
rect 8232 66 8260 2244
rect 8288 94 8316 2272
rect 8344 66 8372 2244
rect 8400 94 8428 2272
rect 8456 66 8484 2244
rect 8512 94 8540 2272
rect 8568 66 8596 2244
rect 8624 94 8652 2272
rect 8680 66 8708 2244
rect 8736 94 8764 2272
rect 8792 66 8820 2244
rect 8848 94 8876 2272
rect 8904 66 8932 2244
rect 8960 94 8988 2272
rect 9016 66 9044 2244
rect 9072 94 9100 2272
rect 9128 66 9156 2244
rect 9184 94 9212 2272
rect 9240 66 9268 2244
rect 9296 94 9324 2272
rect 9352 66 9380 2244
rect 9408 94 9436 2272
rect 9464 66 9492 2244
rect 9520 94 9548 2272
rect 9576 66 9604 2244
rect 9632 94 9660 2272
rect 9688 66 9716 2244
rect 9744 94 9772 2272
rect 9800 66 9828 2244
rect 9856 94 9884 2272
rect 9912 66 9940 2244
rect 9968 94 9996 2272
rect 10024 66 10052 2244
rect 10080 94 10108 2272
rect 10136 66 10164 2244
rect 10192 94 10220 2272
rect 10248 66 10276 2244
rect 10304 94 10332 2272
rect 10360 66 10388 2244
rect 10416 94 10444 2272
rect 10472 66 10500 2244
rect 10528 94 10556 2272
rect 10584 66 10612 2244
rect 10640 94 10668 2272
rect 10696 66 10724 2244
rect 10752 94 10780 2272
rect 10808 66 10836 2244
rect 10864 94 10892 2272
rect 10920 66 10948 2244
rect 10976 94 11004 2272
rect 11032 66 11060 2244
rect 11088 94 11146 2272
rect 0 0 11146 66
<< obsm2 >>
rect 0 66 28 2338
rect 56 2272 196 2338
rect 56 94 84 2272
rect 112 66 140 2244
rect 0 0 140 66
rect 168 0 196 2272
rect 224 66 252 2338
rect 280 2272 420 2338
rect 280 94 308 2272
rect 336 66 364 2244
rect 224 0 364 66
rect 392 0 420 2272
rect 448 66 476 2338
rect 504 2272 644 2338
rect 504 94 532 2272
rect 560 66 588 2244
rect 448 0 588 66
rect 616 0 644 2272
rect 672 66 700 2338
rect 728 2272 868 2338
rect 728 94 756 2272
rect 784 66 812 2244
rect 672 0 812 66
rect 840 0 868 2272
rect 896 66 924 2338
rect 952 2272 1092 2338
rect 952 94 980 2272
rect 1008 66 1036 2244
rect 896 0 1036 66
rect 1064 0 1092 2272
rect 1120 66 1148 2338
rect 1176 2272 1316 2338
rect 1176 94 1204 2272
rect 1232 66 1260 2244
rect 1120 0 1260 66
rect 1288 0 1316 2272
rect 1344 66 1372 2338
rect 1400 2272 1540 2338
rect 1400 94 1428 2272
rect 1456 66 1484 2244
rect 1344 0 1484 66
rect 1512 0 1540 2272
rect 1568 66 1596 2338
rect 1624 2272 1764 2338
rect 1624 94 1652 2272
rect 1680 66 1708 2244
rect 1568 0 1708 66
rect 1736 0 1764 2272
rect 1792 66 1820 2338
rect 1848 2272 1988 2338
rect 1848 94 1876 2272
rect 1904 66 1932 2244
rect 1792 0 1932 66
rect 1960 0 1988 2272
rect 2016 66 2044 2338
rect 2072 2272 2212 2338
rect 2072 94 2100 2272
rect 2128 66 2156 2244
rect 2016 0 2156 66
rect 2184 0 2212 2272
rect 2240 66 2268 2338
rect 2296 2272 2436 2338
rect 2296 94 2324 2272
rect 2352 66 2380 2244
rect 2240 0 2380 66
rect 2408 0 2436 2272
rect 2464 66 2492 2338
rect 2520 2272 2660 2338
rect 2520 94 2548 2272
rect 2576 66 2604 2244
rect 2464 0 2604 66
rect 2632 0 2660 2272
rect 2688 66 2716 2338
rect 2744 2272 2884 2338
rect 2744 94 2772 2272
rect 2800 66 2828 2244
rect 2688 0 2828 66
rect 2856 0 2884 2272
rect 2912 66 2940 2338
rect 2968 2272 3108 2338
rect 2968 94 2996 2272
rect 3024 66 3052 2244
rect 2912 0 3052 66
rect 3080 0 3108 2272
rect 3136 66 3164 2338
rect 3192 2272 3332 2338
rect 3192 94 3220 2272
rect 3248 66 3276 2244
rect 3136 0 3276 66
rect 3304 0 3332 2272
rect 3360 66 3388 2338
rect 3416 2272 3556 2338
rect 3416 94 3444 2272
rect 3472 66 3500 2244
rect 3360 0 3500 66
rect 3528 0 3556 2272
rect 3584 66 3612 2338
rect 3640 2272 3780 2338
rect 3640 94 3668 2272
rect 3696 66 3724 2244
rect 3584 0 3724 66
rect 3752 0 3780 2272
rect 3808 66 3836 2338
rect 3864 2272 4004 2338
rect 3864 94 3892 2272
rect 3920 66 3948 2244
rect 3808 0 3948 66
rect 3976 0 4004 2272
rect 4032 66 4060 2338
rect 4088 2272 4228 2338
rect 4088 94 4116 2272
rect 4144 66 4172 2244
rect 4032 0 4172 66
rect 4200 0 4228 2272
rect 4256 66 4284 2338
rect 4312 2272 4452 2338
rect 4312 94 4340 2272
rect 4368 66 4396 2244
rect 4256 0 4396 66
rect 4424 0 4452 2272
rect 4480 66 4508 2338
rect 4536 2272 4676 2338
rect 4536 94 4564 2272
rect 4592 66 4620 2244
rect 4480 0 4620 66
rect 4648 0 4676 2272
rect 4704 66 4732 2338
rect 4760 2272 4900 2338
rect 4760 94 4788 2272
rect 4816 66 4844 2244
rect 4704 0 4844 66
rect 4872 0 4900 2272
rect 4928 66 4956 2338
rect 4984 2272 5124 2338
rect 4984 94 5012 2272
rect 5040 66 5068 2244
rect 4928 0 5068 66
rect 5096 0 5124 2272
rect 5152 66 5180 2338
rect 5208 2272 5348 2338
rect 5208 94 5236 2272
rect 5264 66 5292 2244
rect 5152 0 5292 66
rect 5320 0 5348 2272
rect 5376 66 5404 2338
rect 5432 2272 5572 2338
rect 5432 94 5460 2272
rect 5488 66 5516 2244
rect 5376 0 5516 66
rect 5544 0 5572 2272
rect 5600 66 5628 2338
rect 5656 2272 5796 2338
rect 5656 94 5684 2272
rect 5712 66 5740 2244
rect 5600 0 5740 66
rect 5768 0 5796 2272
rect 5824 66 5852 2338
rect 5880 2272 6020 2338
rect 5880 94 5908 2272
rect 5936 66 5964 2244
rect 5824 0 5964 66
rect 5992 0 6020 2272
rect 6048 66 6076 2338
rect 6104 2272 6244 2338
rect 6104 94 6132 2272
rect 6160 66 6188 2244
rect 6048 0 6188 66
rect 6216 0 6244 2272
rect 6272 66 6300 2338
rect 6328 2272 6468 2338
rect 6328 94 6356 2272
rect 6384 66 6412 2244
rect 6272 0 6412 66
rect 6440 0 6468 2272
rect 6496 66 6524 2338
rect 6552 2272 6692 2338
rect 6552 94 6580 2272
rect 6608 66 6636 2244
rect 6496 0 6636 66
rect 6664 0 6692 2272
rect 6720 66 6748 2338
rect 6776 2272 6916 2338
rect 6776 94 6804 2272
rect 6832 66 6860 2244
rect 6720 0 6860 66
rect 6888 0 6916 2272
rect 6944 66 6972 2338
rect 7000 2272 7140 2338
rect 7000 94 7028 2272
rect 7056 66 7084 2244
rect 6944 0 7084 66
rect 7112 0 7140 2272
rect 7168 66 7196 2338
rect 7224 2272 7364 2338
rect 7224 94 7252 2272
rect 7280 66 7308 2244
rect 7168 0 7308 66
rect 7336 0 7364 2272
rect 7392 66 7420 2338
rect 7448 2272 7588 2338
rect 7448 94 7476 2272
rect 7504 66 7532 2244
rect 7392 0 7532 66
rect 7560 0 7588 2272
rect 7616 66 7644 2338
rect 7672 2272 7812 2338
rect 7672 94 7700 2272
rect 7728 66 7756 2244
rect 7616 0 7756 66
rect 7784 0 7812 2272
rect 7840 66 7868 2338
rect 7896 2272 8036 2338
rect 7896 94 7924 2272
rect 7952 66 7980 2244
rect 7840 0 7980 66
rect 8008 0 8036 2272
rect 8064 66 8092 2338
rect 8120 2272 8260 2338
rect 8120 94 8148 2272
rect 8176 66 8204 2244
rect 8064 0 8204 66
rect 8232 0 8260 2272
rect 8288 66 8316 2338
rect 8344 2272 8484 2338
rect 8344 94 8372 2272
rect 8400 66 8428 2244
rect 8288 0 8428 66
rect 8456 0 8484 2272
rect 8512 66 8540 2338
rect 8568 2272 8708 2338
rect 8568 94 8596 2272
rect 8624 66 8652 2244
rect 8512 0 8652 66
rect 8680 0 8708 2272
rect 8736 66 8764 2338
rect 8792 2272 8932 2338
rect 8792 94 8820 2272
rect 8848 66 8876 2244
rect 8736 0 8876 66
rect 8904 0 8932 2272
rect 8960 66 8988 2338
rect 9016 2272 9156 2338
rect 9016 94 9044 2272
rect 9072 66 9100 2244
rect 8960 0 9100 66
rect 9128 0 9156 2272
rect 9184 66 9212 2338
rect 9240 2272 9380 2338
rect 9240 94 9268 2272
rect 9296 66 9324 2244
rect 9184 0 9324 66
rect 9352 0 9380 2272
rect 9408 66 9436 2338
rect 9464 2272 9604 2338
rect 9464 94 9492 2272
rect 9520 66 9548 2244
rect 9408 0 9548 66
rect 9576 0 9604 2272
rect 9632 66 9660 2338
rect 9688 2272 9828 2338
rect 9688 94 9716 2272
rect 9744 66 9772 2244
rect 9632 0 9772 66
rect 9800 0 9828 2272
rect 9856 66 9884 2338
rect 9912 2272 10052 2338
rect 9912 94 9940 2272
rect 9968 66 9996 2244
rect 9856 0 9996 66
rect 10024 0 10052 2272
rect 10080 66 10108 2338
rect 10136 2272 10276 2338
rect 10136 94 10164 2272
rect 10192 66 10220 2244
rect 10080 0 10220 66
rect 10248 0 10276 2272
rect 10304 66 10332 2338
rect 10360 2272 10500 2338
rect 10360 94 10388 2272
rect 10416 66 10444 2244
rect 10304 0 10444 66
rect 10472 0 10500 2272
rect 10528 66 10556 2338
rect 10584 2272 10724 2338
rect 10584 94 10612 2272
rect 10640 66 10668 2244
rect 10528 0 10668 66
rect 10696 0 10724 2272
rect 10752 66 10780 2338
rect 10808 2272 11146 2338
rect 10808 94 10836 2272
rect 10864 66 10892 2244
rect 10752 0 10892 66
rect 10920 0 10948 2272
rect 10976 66 11004 2244
rect 11032 94 11060 2272
rect 11088 66 11146 2244
rect 10976 0 11146 66
<< obsm3 >>
rect 0 2272 11146 2338
rect 0 126 60 2272
rect 120 66 180 2212
rect 240 126 300 2272
rect 360 66 420 2212
rect 480 126 540 2272
rect 600 66 660 2212
rect 720 126 780 2272
rect 840 66 900 2212
rect 960 126 1020 2272
rect 1080 66 1140 2212
rect 1200 126 1260 2272
rect 1320 66 1380 2212
rect 1440 126 1500 2272
rect 1560 66 1620 2212
rect 1680 126 1740 2272
rect 1800 66 1860 2212
rect 1920 126 1980 2272
rect 2040 66 2100 2212
rect 2160 126 2220 2272
rect 2280 66 2340 2212
rect 2400 126 2460 2272
rect 2520 66 2580 2212
rect 2640 126 2700 2272
rect 2760 66 2820 2212
rect 2880 126 2940 2272
rect 3000 66 3060 2212
rect 3120 126 3180 2272
rect 3240 66 3300 2212
rect 3360 126 3420 2272
rect 3480 66 3540 2212
rect 3600 126 3660 2272
rect 3720 66 3780 2212
rect 3840 126 3900 2272
rect 3960 66 4020 2212
rect 4080 126 4140 2272
rect 4200 66 4260 2212
rect 4320 126 4380 2272
rect 4440 66 4500 2212
rect 4560 126 4620 2272
rect 4680 66 4740 2212
rect 4800 126 4860 2272
rect 4920 66 4980 2212
rect 5040 126 5100 2272
rect 5160 66 5220 2212
rect 5280 126 5340 2272
rect 5400 66 5460 2212
rect 5520 126 5580 2272
rect 5640 66 5700 2212
rect 5760 126 5820 2272
rect 5880 66 5940 2212
rect 6000 126 6060 2272
rect 6120 66 6180 2212
rect 6240 126 6300 2272
rect 6360 66 6420 2212
rect 6480 126 6540 2272
rect 6600 66 6660 2212
rect 6720 126 6780 2272
rect 6840 66 6900 2212
rect 6960 126 7020 2272
rect 7080 66 7140 2212
rect 7200 126 7260 2272
rect 7320 66 7380 2212
rect 7440 126 7500 2272
rect 7560 66 7620 2212
rect 7680 126 7740 2272
rect 7800 66 7860 2212
rect 7920 126 7980 2272
rect 8040 66 8100 2212
rect 8160 126 8220 2272
rect 8280 66 8340 2212
rect 8400 126 8460 2272
rect 8520 66 8580 2212
rect 8640 126 8700 2272
rect 8760 66 8820 2212
rect 8880 126 8940 2272
rect 9000 66 9060 2212
rect 9120 126 9180 2272
rect 9240 66 9300 2212
rect 9360 126 9420 2272
rect 9480 66 9540 2212
rect 9600 126 9660 2272
rect 9720 66 9780 2212
rect 9840 126 9900 2272
rect 9960 66 10020 2212
rect 10080 126 10140 2272
rect 10200 66 10260 2212
rect 10320 126 10380 2272
rect 10440 66 10500 2212
rect 10560 126 10620 2272
rect 10680 66 10740 2212
rect 10800 126 10860 2272
rect 10920 66 10980 2212
rect 11040 126 11146 2272
rect 0 0 11146 66
<< obsm4 >>
rect 0 2272 11146 2338
rect 0 66 60 2212
rect 120 2027 420 2272
rect 120 126 180 2027
rect 240 311 300 1967
rect 360 371 420 2027
rect 480 311 540 2212
rect 240 66 540 311
rect 600 126 660 2272
rect 720 66 780 2212
rect 840 126 900 2272
rect 960 66 1020 2212
rect 1080 126 1140 2272
rect 1200 66 1260 2212
rect 1320 126 1380 2272
rect 1440 66 1500 2212
rect 1560 2027 1860 2272
rect 1560 126 1620 2027
rect 1680 311 1740 1967
rect 1800 371 1860 2027
rect 1920 311 1980 2212
rect 1680 66 1980 311
rect 2040 126 2100 2272
rect 2160 66 2220 2212
rect 2280 126 2340 2272
rect 2400 66 2460 2212
rect 2520 126 2580 2272
rect 2640 66 2700 2212
rect 2760 126 2820 2272
rect 2880 66 2940 2212
rect 3000 2027 3300 2272
rect 3000 126 3060 2027
rect 3120 311 3180 1967
rect 3240 371 3300 2027
rect 3360 311 3420 2212
rect 3120 66 3420 311
rect 3480 126 3540 2272
rect 3600 66 3660 2212
rect 3720 126 3780 2272
rect 3840 66 3900 2212
rect 3960 126 4020 2272
rect 4080 66 4140 2212
rect 4200 126 4260 2272
rect 4320 66 4380 2212
rect 4440 2027 4740 2272
rect 4440 126 4500 2027
rect 4560 311 4620 1967
rect 4680 371 4740 2027
rect 4800 311 4860 2212
rect 4560 66 4860 311
rect 4920 126 4980 2272
rect 5040 66 5100 2212
rect 5160 126 5220 2272
rect 5280 66 5340 2212
rect 5400 126 5460 2272
rect 5520 66 5580 2212
rect 5640 126 5700 2272
rect 5760 66 5820 2212
rect 5880 2027 6180 2272
rect 5880 126 5940 2027
rect 6000 311 6060 1967
rect 6120 371 6180 2027
rect 6240 311 6300 2212
rect 6000 66 6300 311
rect 6360 126 6420 2272
rect 6480 66 6540 2212
rect 6600 126 6660 2272
rect 6720 66 6780 2212
rect 6840 126 6900 2272
rect 6960 66 7020 2212
rect 7080 126 7140 2272
rect 7200 66 7260 2212
rect 7320 2027 7620 2272
rect 7320 126 7380 2027
rect 7440 311 7500 1967
rect 7560 371 7620 2027
rect 7680 311 7740 2212
rect 7440 66 7740 311
rect 7800 126 7860 2272
rect 7920 66 7980 2212
rect 8040 126 8100 2272
rect 8160 66 8220 2212
rect 8280 126 8340 2272
rect 8400 66 8460 2212
rect 8520 126 8580 2272
rect 8640 66 8700 2212
rect 8760 2027 9060 2272
rect 8760 126 8820 2027
rect 8880 311 8940 1967
rect 9000 371 9060 2027
rect 9120 311 9180 2212
rect 8880 66 9180 311
rect 9240 126 9300 2272
rect 9360 66 9420 2212
rect 9480 126 9540 2272
rect 9600 66 9660 2212
rect 9720 126 9780 2272
rect 9840 66 9900 2212
rect 9960 126 10020 2272
rect 10080 66 10140 2212
rect 10200 2027 10500 2272
rect 10200 126 10260 2027
rect 10320 311 10380 1967
rect 10440 371 10500 2027
rect 10560 311 10620 2212
rect 10320 66 10620 311
rect 10680 126 10740 2272
rect 10800 66 10860 2212
rect 10920 126 10980 2272
rect 11040 66 11146 2212
rect 0 0 11146 66
<< obsm5 >>
rect 0 2003 11146 2338
rect 0 655 320 2003
rect 640 335 960 1683
rect 1280 655 1600 2003
rect 1920 335 2240 1683
rect 2560 655 2880 2003
rect 3200 335 3520 1683
rect 3840 655 4160 2003
rect 4480 335 4800 1683
rect 5120 655 5440 2003
rect 5760 335 6080 1683
rect 6400 655 6720 2003
rect 7040 335 7360 1683
rect 7680 655 8000 2003
rect 8320 335 8640 1683
rect 8960 655 9280 2003
rect 9600 335 9920 1683
rect 10240 655 11146 2003
rect 0 0 11146 335
<< properties >>
string FIXED_BBOX 0 0 11146 2338
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2113884
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1957848
<< end >>
