magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 1546 850 1570 874 ne
tri 1616 850 1640 874 nw
rect 823 792 899 832
tri 899 792 939 832 sw
rect 823 786 939 792
rect 77 628 287 758
tri 879 726 939 786 ne
tri 939 726 1005 792 sw
tri 939 684 981 726 ne
rect 981 707 1301 726
tri 1301 707 1320 726 sw
tri 1325 707 1412 794 ne
rect 1412 753 1453 794
tri 1453 753 1504 804 sw
rect 1412 707 1592 753
rect 981 684 1320 707
tri 1263 629 1318 684 ne
rect 1318 654 1320 684
tri 1320 654 1373 707 sw
rect 1318 629 1599 654
tri 38 253 77 292 se
rect 77 253 154 628
rect 680 587 684 629
tri 684 587 726 629 sw
rect 680 583 726 587
tri 666 551 698 583 ne
tri 355 488 398 531 se
rect 398 503 652 531
tri 398 488 413 503 nw
tri 351 484 355 488 se
rect 355 484 379 488
tri 340 395 351 406 se
rect 351 395 379 484
tri 379 469 398 488 nw
tri 323 378 340 395 se
rect 340 394 379 395
rect 340 378 346 394
rect 277 361 346 378
tri 346 361 379 394 nw
tri 277 292 346 361 nw
tri 449 339 483 373 sw
tri 604 361 624 381 se
rect 624 343 652 503
rect 698 417 726 583
rect 1200 570 1212 616
tri 1212 570 1258 616 sw
tri 1318 608 1339 629 ne
rect 1339 608 1599 629
tri 1218 530 1258 570 ne
tri 1258 530 1298 570 sw
tri 1258 527 1261 530 ne
tri 726 417 760 451 sw
tri 652 361 686 395 sw
rect 698 389 764 417
tri 746 371 764 389 ne
rect 1261 372 1298 530
tri 1298 372 1332 406 sw
tri 734 343 752 361 sw
tri 1070 343 1088 361 se
rect 443 293 533 339
rect 38 220 154 253
tri 154 220 211 277 sw
tri 449 259 483 293 nw
tri 523 283 533 293 ne
tri 533 287 585 339 sw
rect 624 315 1088 343
rect 1261 326 1572 372
tri 1440 287 1451 298 se
rect 533 283 1451 287
tri 533 259 557 283 ne
rect 557 259 1451 283
tri 1444 252 1451 259 ne
tri 297 220 317 240 se
tri 363 220 383 240 sw
tri 1667 220 1700 253 se
rect 1700 220 1829 253
rect 38 39 1829 220
use sky130_fd_pr__nfet_01v8__example_55959141808496  sky130_fd_pr__nfet_01v8__example_55959141808496_0
timestamp 1676037725
transform -1 0 1744 0 -1 358
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808497  sky130_fd_pr__nfet_01v8__example_55959141808497_0
timestamp 1676037725
transform -1 0 1154 0 1 158
box -1 0 417 1
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_0
timestamp 1676037725
transform -1 0 484 0 1 158
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808498  sky130_fd_pr__nfet_01v8__example_55959141808498_1
timestamp 1676037725
transform -1 0 312 0 1 158
box -1 0 117 1
use sky130_fd_pr__nfet_01v8__example_55959141808582  sky130_fd_pr__nfet_01v8__example_55959141808582_0
timestamp 1676037725
transform -1 0 1186 0 -1 884
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808583  sky130_fd_pr__nfet_01v8__example_55959141808583_0
timestamp 1676037725
transform -1 0 438 0 -1 884
box -1 0 257 1
use sky130_fd_pr__nfet_01v8__example_55959141808583  sky130_fd_pr__nfet_01v8__example_55959141808583_1
timestamp 1676037725
transform -1 0 750 0 -1 884
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808580  sky130_fd_pr__pfet_01v8__example_55959141808580_0
timestamp 1676037725
transform -1 0 1565 0 -1 964
box -1 0 121 1
use sky130_fd_pr__pfet_01v8__example_55959141808580  sky130_fd_pr__pfet_01v8__example_55959141808580_1
timestamp 1676037725
transform 1 0 1621 0 -1 964
box -1 0 121 1
<< properties >>
string GDS_END 43539214
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43520030
<< end >>
