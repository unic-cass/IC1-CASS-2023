magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< metal1 >>
tri 26924 234 27014 324 sw
rect 26924 205 27014 234
tri 26964 155 27014 205 ne
tri 27014 155 27093 234 sw
tri 27014 103 27066 155 ne
rect 27066 103 27849 155
tri 27849 103 27901 155 sw
tri 27827 59 27871 103 ne
rect 27871 81 27901 103
tri 27901 81 27923 103 sw
rect 27871 39 27923 81
rect 27716 -555 28669 -547
tri 28669 -555 28677 -547 sw
rect 27716 -579 28677 -555
tri 28655 -601 28677 -579 ne
tri 28677 -601 28723 -555 sw
tri 28677 -615 28691 -601 ne
tri 27981 -850 27984 -847 se
tri 27981 -899 27984 -896 ne
rect 28691 -1037 28723 -601
tri 28691 -1069 28723 -1037 ne
tri 28723 -1057 28757 -1023 sw
rect 28723 -1069 29018 -1057
tri 28723 -1103 28757 -1069 ne
rect 28757 -1103 29018 -1069
tri 30203 -1921 30266 -1858 ne
tri 30328 -1921 30391 -1858 nw
tri 30173 -2180 30268 -2085 se
tri 36776 -2118 36784 -2110 se
rect 31194 -2137 36784 -2118
rect 31194 -2146 36798 -2137
tri 36768 -2162 36784 -2146 ne
rect 36784 -2162 36798 -2146
tri 30734 -2253 30798 -2189 ne
tri 29988 -2711 30036 -2663 se
rect 29916 -2925 30036 -2711
tri 29966 -2995 30036 -2925 ne
tri 30031 -3184 30105 -3110 se
rect 30105 -3162 30491 -3110
tri 30105 -3184 30127 -3162 nw
tri 29977 -3238 30031 -3184 se
rect 30031 -3238 30051 -3184
tri 30051 -3238 30105 -3184 nw
rect 29689 -3266 30023 -3238
tri 30023 -3266 30051 -3238 nw
tri 27254 -4371 27288 -4337 se
tri 26925 -4410 26964 -4371 se
rect 26964 -4399 27288 -4371
rect 26964 -4410 26977 -4399
tri 26977 -4410 26988 -4399 nw
rect 26702 -4451 26936 -4410
tri 26936 -4451 26977 -4410 nw
tri 26702 -4485 26736 -4451 nw
tri 27162 -5083 27192 -5053 se
tri 27244 -5083 27274 -5053 sw
tri 26788 -5558 26822 -5524 se
tri 26869 -5554 26965 -5458 nw
rect 30798 -5515 30826 -2189
tri 32128 -2255 32146 -2237 se
rect 32146 -2255 32975 -2237
rect 31207 -2256 32975 -2255
tri 32975 -2256 32994 -2237 sw
tri 33972 -2256 33978 -2250 se
rect 31207 -2265 33978 -2256
rect 31207 -2283 32174 -2265
tri 32174 -2283 32192 -2265 nw
tri 32360 -2311 32371 -2300 sw
tri 32541 -2311 32559 -2293 se
rect 32559 -2311 32852 -2293
rect 32360 -2321 32852 -2311
rect 32360 -2339 32587 -2321
tri 32587 -2339 32605 -2321 nw
tri 32360 -2352 32373 -2339 nw
tri 32787 -2358 32824 -2321 ne
rect 32824 -2330 32852 -2321
tri 32852 -2330 32889 -2293 sw
tri 32910 -2302 32947 -2265 ne
rect 32947 -2302 33978 -2265
rect 32824 -2331 35722 -2330
tri 35722 -2331 35723 -2330 sw
rect 32824 -2358 36431 -2331
tri 35693 -2359 35694 -2358 ne
rect 35694 -2359 36431 -2358
tri 36407 -2383 36431 -2359 ne
tri 31207 -2442 31233 -2416 sw
rect 31207 -2470 34575 -2442
rect 31174 -2542 34334 -2498
rect 31174 -2550 31696 -2542
tri 31696 -2550 31704 -2542 nw
tri 34326 -2550 34334 -2542 ne
rect 34334 -2550 34335 -2542
rect 31174 -2574 31226 -2550
tri 31937 -2595 31961 -2571 se
rect 31961 -2595 31976 -2571
rect 31445 -2604 31976 -2595
rect 31445 -2623 31961 -2604
tri 31226 -3212 31260 -3178 sw
tri 31226 -3298 31260 -3264 nw
tri 31226 -3459 31260 -3425 sw
tri 31681 -3459 31715 -3425 se
tri 31767 -3459 31801 -3425 sw
tri 33000 -3459 33016 -3443 se
rect 31226 -3487 33018 -3459
tri 33008 -3495 33016 -3487 ne
tri 31011 -3589 31022 -3578 se
tri 31050 -3589 31061 -3578 sw
tri 31883 -3645 31911 -3617 ne
tri 34353 -3681 34387 -3647 se
tri 34439 -3681 34445 -3675 sw
tri 31011 -3728 31022 -3717 ne
tri 31050 -3728 31061 -3717 nw
tri 35009 -3730 35017 -3722 sw
tri 35009 -3768 35019 -3758 nw
tri 31377 -3812 31411 -3778 sw
rect 31377 -3840 32408 -3812
tri 32382 -3866 32408 -3840 ne
tri 32408 -3865 32461 -3812 sw
tri 34158 -3853 34186 -3825 sw
rect 32408 -3866 32461 -3865
tri 31226 -3912 31260 -3878 sw
tri 31771 -3912 31795 -3888 se
tri 32408 -3919 32461 -3866 ne
tri 32461 -3919 32515 -3865 sw
tri 32743 -3919 32759 -3903 se
rect 34158 -3908 34482 -3853
tri 31226 -3959 31245 -3940 nw
tri 32461 -3947 32489 -3919 ne
rect 32489 -3947 32759 -3919
tri 32751 -3955 32759 -3947 ne
rect 34155 -3910 34482 -3908
rect 34155 -3955 34158 -3910
tri 34158 -3955 34203 -3910 nw
tri 31126 -4112 31160 -4078 sw
rect 31126 -4140 35791 -4112
tri 31126 -4174 31160 -4140 nw
tri 31532 -4418 31566 -4384 sw
rect 32852 -4446 34503 -4418
tri 34503 -4446 34531 -4418 sw
tri 31532 -4477 31539 -4470 nw
tri 33310 -4508 33344 -4474 se
rect 33344 -4502 34042 -4474
rect 33344 -4508 33372 -4502
rect 32626 -4536 33372 -4508
tri 33372 -4536 33406 -4502 nw
rect 34014 -4614 34042 -4502
tri 34457 -4520 34531 -4446 ne
tri 34531 -4467 34552 -4446 sw
rect 34531 -4520 34559 -4467
tri 34531 -4548 34559 -4520 ne
tri 35109 -4662 35147 -4624 nw
tri 32953 -5350 32991 -5312 se
rect 38125 -5336 38157 -5320
tri 38157 -5336 38173 -5320 sw
tri 26162 -5615 26191 -5586 sw
tri 38121 -5896 38125 -5892 se
rect 38125 -5896 38173 -5336
tri 33132 -6006 33157 -5981 se
rect 32949 -6052 33157 -6006
rect 32949 -6093 32995 -6052
tri 33126 -6083 33157 -6052 ne
<< metal2 >>
rect 26270 -790 26444 -715
tri 26444 -790 26519 -715 sw
rect 26270 -845 26884 -790
tri 26390 -920 26465 -845 ne
rect 26465 -920 26884 -845
rect 27871 -913 27923 -89
rect 33875 -130 33916 -78
tri 33717 -232 33819 -130 ne
rect 33819 -208 33916 -130
tri 33916 -208 33990 -134 sw
rect 33819 -232 33967 -208
tri 33967 -232 33990 -208 nw
rect 27984 -702 29111 -632
rect 27984 -847 28112 -702
tri 28112 -784 28194 -702 nw
tri 28270 -756 28324 -702 ne
rect 28324 -707 29111 -702
tri 29111 -707 29186 -632 sw
tri 26632 -1066 26778 -920 ne
tri 27871 -965 27923 -913 ne
tri 27923 -915 27925 -913 sw
rect 27923 -965 27925 -915
tri 27923 -967 27925 -965 ne
tri 27925 -967 27977 -915 sw
tri 27925 -995 27953 -967 ne
rect 27953 -995 28437 -967
tri 28183 -1511 28229 -1465 ne
tri 26343 -2391 26377 -2357 sw
tri 26343 -2477 26377 -2443 nw
tri 26613 -2498 26639 -2472 se
tri 26667 -2498 26701 -2464 sw
tri 26292 -4021 26316 -3997 se
tri 26342 -4015 26344 -4013 sw
rect 26342 -4021 26344 -4015
tri 26087 -4172 26110 -4149 ne
rect 26136 -4151 26137 -4149
tri 26137 -4151 26139 -4149 nw
tri 26771 -4605 26773 -4603 se
tri 27236 -5369 27288 -5317 se
rect 27288 -5339 27340 -4399
tri 28176 -4427 28229 -4374 se
rect 28229 -4422 28257 -1465
tri 28257 -1481 28273 -1465 nw
tri 33590 -2065 33664 -1991 se
rect 33664 -2019 37134 -1991
tri 33664 -2065 33710 -2019 nw
rect 30698 -2146 31155 -2118
tri 33522 -2133 33590 -2065 se
rect 33590 -2133 33596 -2065
tri 33596 -2133 33664 -2065 nw
tri 36574 -2102 36627 -2049 se
rect 36627 -2069 37032 -2049
tri 37032 -2069 37052 -2049 sw
tri 37096 -2057 37134 -2019 ne
tri 37134 -2055 37198 -1991 sw
rect 37134 -2057 37198 -2055
rect 36627 -2077 37052 -2069
tri 37134 -2075 37152 -2057 ne
tri 36627 -2102 36652 -2077 nw
tri 30826 -2189 30869 -2146 nw
tri 31881 -2256 31911 -2226 ne
tri 30707 -2478 30756 -2429 se
rect 30756 -2457 31155 -2429
rect 30756 -2478 30765 -2457
tri 30765 -2478 30786 -2457 nw
rect 29767 -2506 30737 -2478
tri 30737 -2506 30765 -2478 nw
tri 29534 -2554 29582 -2506 sw
tri 29767 -2530 29791 -2506 nw
tri 29530 -2606 29582 -2554 ne
tri 29582 -2587 29615 -2554 sw
rect 29582 -2606 31180 -2587
tri 29582 -2615 29591 -2606 ne
rect 29591 -2615 31180 -2606
rect 30304 -3912 30332 -3458
rect 31911 -3589 31963 -2226
tri 31963 -2272 32009 -2226 nw
rect 33522 -2653 33574 -2133
tri 33574 -2155 33596 -2133 nw
rect 33875 -2166 34143 -2114
tri 34121 -2188 34143 -2166 ne
tri 34143 -2187 34216 -2114 sw
tri 36521 -2155 36574 -2102 se
tri 36574 -2155 36627 -2102 nw
tri 36955 -2122 37000 -2077 ne
rect 34143 -2188 34216 -2187
tri 34143 -2209 34164 -2188 ne
tri 33574 -2653 33596 -2631 sw
tri 33522 -2727 33596 -2653 ne
tri 33596 -2727 33670 -2653 sw
tri 33596 -2749 33618 -2727 ne
rect 33144 -3472 33223 -3443
tri 33223 -3472 33252 -3443 sw
rect 33144 -3495 33252 -3472
tri 33221 -3526 33252 -3495 ne
tri 33252 -3526 33306 -3472 sw
tri 33252 -3554 33280 -3526 ne
rect 33280 -3554 33483 -3526
tri 30332 -3912 30366 -3878 sw
rect 30304 -3940 31174 -3912
tri 31251 -4136 31325 -4062 se
rect 31325 -4084 31377 -3840
tri 31795 -3982 31837 -3940 ne
tri 31325 -4136 31377 -4084 nw
rect 28229 -4427 28252 -4422
tri 28252 -4427 28257 -4422 nw
tri 31243 -4144 31251 -4136 se
rect 31251 -4144 31271 -4136
tri 28153 -4510 28176 -4487 se
rect 28176 -4510 28205 -4427
tri 28205 -4474 28252 -4427 nw
rect 27236 -5821 27288 -5369
tri 27288 -5391 27340 -5339 nw
tri 28296 -5423 28330 -5389 se
rect 31243 -5931 31271 -4144
tri 31271 -4190 31325 -4136 nw
rect 31837 -4942 31889 -3940
tri 31889 -3974 31923 -3940 nw
tri 31889 -4942 31931 -4900 sw
rect 32748 -4909 32800 -4891
tri 31837 -5036 31931 -4942 ne
tri 31931 -5036 32025 -4942 sw
tri 32748 -4961 32800 -4909 ne
tri 32800 -4953 32866 -4887 sw
rect 32800 -4961 32866 -4953
tri 32800 -4975 32814 -4961 ne
tri 31931 -5130 32025 -5036 ne
tri 32025 -5130 32119 -5036 sw
tri 32025 -5224 32119 -5130 ne
tri 32119 -5224 32213 -5130 sw
tri 32792 -5155 32814 -5133 se
rect 32814 -5155 32866 -4961
rect 33455 -5018 33483 -3554
rect 33618 -4628 33670 -2727
rect 33847 -3131 33899 -2844
tri 33899 -2878 33933 -2844 nw
tri 33847 -3138 33854 -3131 ne
tri 33847 -3247 33854 -3240 se
rect 33854 -3247 33899 -3131
rect 33847 -4904 33899 -3247
rect 34055 -4421 34094 -2302
tri 34122 -2411 34164 -2369 se
rect 34164 -2391 34216 -2188
tri 36475 -2201 36521 -2155 se
rect 36521 -2201 36528 -2155
tri 36528 -2201 36574 -2155 nw
rect 36475 -2331 36503 -2201
tri 36503 -2226 36528 -2201 nw
rect 37000 -2367 37052 -2077
rect 34164 -2411 34169 -2391
rect 34122 -4361 34169 -2411
tri 34169 -2438 34216 -2391 nw
rect 37152 -2385 37198 -2057
tri 36660 -2448 36694 -2414 ne
tri 36746 -2436 36768 -2414 nw
rect 37152 -2431 37906 -2385
tri 34501 -3095 34575 -3021 se
rect 34575 -3043 34627 -2494
tri 34627 -2570 34703 -2494 nw
tri 34575 -3095 34627 -3043 nw
tri 34495 -3101 34501 -3095 se
rect 34501 -3101 34547 -3095
rect 34495 -3567 34547 -3101
tri 34547 -3123 34575 -3095 nw
rect 34686 -3108 34738 -3030
tri 34686 -3160 34738 -3108 ne
tri 34738 -3142 34794 -3086 sw
rect 34738 -3160 34794 -3142
tri 34738 -3216 34794 -3160 ne
tri 34794 -3216 34868 -3142 sw
tri 34794 -3261 34839 -3216 ne
rect 34658 -3828 34714 -3614
rect 34839 -3759 34868 -3216
tri 34839 -3788 34868 -3759 ne
tri 34868 -3764 34918 -3714 sw
rect 34868 -3788 35878 -3764
tri 34658 -3884 34714 -3828 ne
tri 34714 -3862 34766 -3810 sw
tri 34868 -3816 34896 -3788 ne
rect 34896 -3816 35878 -3788
rect 34714 -3879 35603 -3862
tri 35603 -3879 35620 -3862 sw
tri 35815 -3879 35878 -3816 ne
rect 34714 -3884 35620 -3879
tri 34351 -3944 34387 -3908 ne
rect 34387 -4090 34439 -3908
tri 34439 -3948 34479 -3908 nw
tri 34714 -3914 34744 -3884 ne
rect 34744 -3914 35620 -3884
tri 35581 -3942 35609 -3914 ne
rect 35609 -3942 35620 -3914
tri 35620 -3942 35683 -3879 sw
tri 35609 -3964 35631 -3942 ne
rect 35631 -4029 35683 -3942
tri 34439 -4090 34457 -4072 sw
tri 35631 -4081 35683 -4029 ne
tri 35683 -4052 35728 -4007 sw
rect 35683 -4081 35728 -4052
rect 34387 -4094 34457 -4090
tri 34387 -4164 34457 -4094 ne
tri 34457 -4164 34531 -4090 sw
tri 35683 -4126 35728 -4081 ne
tri 35728 -4126 35802 -4052 sw
tri 34457 -4216 34509 -4164 ne
rect 34509 -4200 35687 -4164
tri 35687 -4200 35723 -4164 sw
tri 35728 -4200 35802 -4126 ne
tri 35802 -4200 35876 -4126 sw
rect 34509 -4216 35723 -4200
tri 35665 -4252 35701 -4216 ne
rect 35701 -4252 35723 -4216
tri 35723 -4252 35775 -4200 sw
tri 35802 -4252 35854 -4200 ne
rect 35854 -4207 35940 -4200
tri 35940 -4207 35947 -4200 sw
rect 35854 -4252 35947 -4207
tri 35701 -4318 35767 -4252 ne
rect 35767 -4293 35775 -4252
tri 35775 -4293 35816 -4252 sw
tri 35918 -4281 35947 -4252 ne
tri 35947 -4281 36021 -4207 sw
rect 35767 -4318 35816 -4293
tri 34122 -4408 34169 -4361 ne
tri 34169 -4402 34237 -4334 sw
tri 35497 -4336 35515 -4318 se
rect 35515 -4336 35715 -4318
tri 35715 -4336 35733 -4318 sw
tri 35431 -4402 35497 -4336 se
rect 35497 -4345 35733 -4336
tri 35733 -4345 35742 -4336 sw
rect 35497 -4364 35742 -4345
tri 35497 -4402 35535 -4364 nw
tri 35695 -4402 35733 -4364 ne
rect 35733 -4367 35742 -4364
tri 35742 -4367 35764 -4345 sw
tri 35767 -4367 35816 -4318 ne
tri 35816 -4367 35890 -4293 sw
tri 35947 -4355 36021 -4281 ne
tri 36021 -4355 36095 -4281 sw
rect 35733 -4402 35764 -4367
tri 35764 -4402 35799 -4367 sw
rect 34169 -4408 34237 -4402
tri 34094 -4421 34100 -4415 sw
rect 34055 -4450 34100 -4421
tri 34055 -4495 34100 -4450 ne
tri 34100 -4465 34144 -4421 sw
tri 34169 -4465 34226 -4408 ne
rect 34226 -4465 34237 -4408
tri 34237 -4465 34300 -4402 sw
tri 35425 -4408 35431 -4402 se
rect 35431 -4408 35471 -4402
rect 34100 -4495 34144 -4465
tri 34144 -4495 34174 -4465 sw
tri 34100 -4569 34174 -4495 ne
tri 34174 -4517 34196 -4495 sw
tri 34226 -4517 34278 -4465 ne
rect 34278 -4517 34828 -4465
rect 34174 -4569 34196 -4517
tri 34196 -4569 34248 -4517 sw
tri 34174 -4621 34226 -4569 ne
rect 34226 -4621 34311 -4569
rect 34776 -4840 34828 -4517
tri 33847 -4956 33899 -4904 ne
tri 33899 -4908 33925 -4882 sw
tri 35054 -4908 35106 -4856 se
rect 35106 -4908 35246 -4856
rect 33899 -4956 35076 -4908
tri 33899 -4960 33903 -4956 ne
rect 33903 -4960 35076 -4956
tri 35076 -4960 35128 -4908 nw
tri 33483 -5018 33494 -5007 sw
rect 33455 -5053 33494 -5018
tri 33455 -5092 33494 -5053 ne
tri 33494 -5092 33568 -5018 sw
tri 35373 -5092 35425 -5040 se
rect 35425 -5060 35471 -4408
tri 35471 -4428 35497 -4402 nw
tri 35733 -4468 35799 -4402 ne
tri 35799 -4419 35816 -4402 sw
tri 35816 -4419 35868 -4367 ne
rect 35868 -4419 35890 -4367
rect 35799 -4468 35816 -4419
tri 35816 -4468 35865 -4419 sw
tri 35868 -4441 35890 -4419 ne
tri 35890 -4441 35964 -4367 sw
tri 36021 -4429 36095 -4355 ne
tri 36095 -4429 36169 -4355 sw
tri 35799 -4534 35865 -4468 ne
tri 35865 -4493 35890 -4468 sw
tri 35890 -4493 35942 -4441 ne
rect 35942 -4493 35964 -4441
rect 35865 -4534 35890 -4493
tri 35890 -4534 35931 -4493 sw
tri 35942 -4515 35964 -4493 ne
tri 35964 -4515 36038 -4441 sw
tri 36095 -4503 36169 -4429 ne
tri 36169 -4503 36243 -4429 sw
tri 35865 -4600 35931 -4534 ne
tri 35931 -4567 35964 -4534 sw
tri 35964 -4567 36016 -4515 ne
rect 36016 -4567 36038 -4515
rect 35931 -4600 35964 -4567
tri 35964 -4600 35997 -4567 sw
tri 36016 -4589 36038 -4567 ne
tri 36038 -4589 36112 -4515 sw
tri 36169 -4577 36243 -4503 ne
tri 36243 -4577 36317 -4503 sw
tri 35931 -4666 35997 -4600 ne
tri 35997 -4641 36038 -4600 sw
tri 36038 -4641 36090 -4589 ne
rect 36090 -4641 36112 -4589
rect 35997 -4666 36038 -4641
tri 36038 -4666 36063 -4641 sw
tri 36090 -4663 36112 -4641 ne
tri 36112 -4663 36186 -4589 sw
tri 36243 -4651 36317 -4577 ne
tri 36317 -4651 36391 -4577 sw
rect 39702 -4619 39812 -4573
tri 35997 -4686 36017 -4666 ne
tri 35983 -4872 36017 -4838 se
rect 36017 -4872 36063 -4666
tri 36112 -4737 36186 -4663 ne
tri 36186 -4737 36260 -4663 sw
tri 36317 -4725 36391 -4651 ne
tri 36391 -4725 36465 -4651 sw
tri 36186 -4811 36260 -4737 ne
tri 36260 -4811 36334 -4737 sw
tri 36391 -4777 36443 -4725 ne
rect 36443 -4777 36515 -4725
tri 36063 -4872 36092 -4843 sw
tri 36260 -4885 36334 -4811 ne
tri 36334 -4885 36408 -4811 sw
tri 36334 -4937 36386 -4885 ne
rect 36386 -4937 36526 -4885
rect 35425 -5092 35439 -5060
tri 35439 -5092 35471 -5060 nw
tri 33494 -5138 33540 -5092 ne
rect 33540 -5138 35393 -5092
tri 35393 -5138 35439 -5092 nw
tri 32777 -5170 32792 -5155 se
rect 32792 -5170 32799 -5155
tri 32524 -5222 32576 -5170 se
rect 32576 -5222 32799 -5170
tri 32799 -5222 32866 -5155 nw
tri 32119 -5252 32147 -5224 ne
rect 32147 -6295 32213 -5224
tri 32504 -5242 32524 -5222 se
rect 32524 -5242 32556 -5222
tri 32265 -5436 32299 -5402 ne
tri 32351 -5423 32372 -5402 nw
rect 32504 -5695 32556 -5242
tri 32556 -5264 32598 -5222 nw
tri 33263 -5262 33264 -5261 se
rect 33263 -5264 33264 -5262
tri 33316 -5264 33350 -5230 sw
rect 39766 -5259 39812 -4619
tri 33111 -5346 33165 -5292 se
tri 33215 -5346 33239 -5322 sw
tri 33570 -5325 33636 -5259 se
rect 33636 -5305 39812 -5259
tri 33636 -5325 33656 -5305 nw
tri 33504 -5391 33570 -5325 se
tri 33570 -5391 33636 -5325 nw
rect 32991 -5434 33043 -5402
tri 33043 -5434 33077 -5400 sw
tri 33461 -5434 33504 -5391 se
rect 33504 -5434 33527 -5391
tri 33527 -5434 33570 -5391 nw
rect 32991 -5460 33492 -5434
tri 32991 -5469 33000 -5460 ne
rect 33000 -5469 33492 -5460
tri 33492 -5469 33527 -5434 nw
tri 32956 -5507 32990 -5473 sw
tri 32504 -5747 32556 -5695 ne
tri 32556 -5738 32621 -5673 sw
rect 32556 -5747 32621 -5738
tri 32556 -5812 32621 -5747 ne
tri 32621 -5812 32695 -5738 sw
tri 32621 -5834 32643 -5812 ne
rect 32643 -6188 32695 -5812
tri 34800 -5876 34824 -5852 sw
rect 33209 -6073 33236 -5981
tri 33236 -6073 33328 -5981 sw
tri 33589 -6018 33619 -5988 se
tri 33671 -6018 33705 -5984 sw
tri 37354 -6053 37358 -6049 ne
rect 33209 -6109 33328 -6073
tri 33290 -6147 33328 -6109 ne
tri 33328 -6147 33402 -6073 sw
tri 38173 -6089 38207 -6055 se
tri 33328 -6221 33402 -6147 ne
tri 33402 -6221 33476 -6147 sw
tri 33402 -6264 33445 -6221 ne
rect 33445 -6264 35057 -6221
tri 32147 -6361 32213 -6295 ne
tri 32213 -6298 32244 -6267 sw
tri 32697 -6298 32727 -6268 se
tri 35023 -6298 35057 -6264 ne
rect 32213 -6361 32727 -6298
tri 32213 -6364 32216 -6361 ne
rect 32216 -6364 32727 -6361
tri 32697 -6394 32727 -6364 ne
tri 26259 -6801 26293 -6767 se
tri 26321 -6801 26355 -6767 sw
tri 41412 -8324 41444 -8292 se
tri 41195 -8404 41229 -8370 nw
tri 41410 -8404 41444 -8370 ne
<< metal3 >>
tri 34559 -3787 34653 -3693 se
tri 34653 -3787 34718 -3722 nw
tri 34467 -3879 34559 -3787 se
rect 34559 -3879 34561 -3787
tri 34561 -3879 34653 -3787 nw
rect 26319 -4665 26385 -4334
tri 26319 -4725 26379 -4665 ne
rect 26379 -4697 26385 -4665
tri 26385 -4697 26445 -4637 sw
rect 26379 -6055 26445 -4697
rect 32722 -8329 32788 -6270
tri 34373 -7363 34467 -7269 se
rect 34467 -7297 34533 -3879
tri 34533 -3907 34561 -3879 nw
tri 34467 -7363 34533 -7297 nw
tri 34279 -7457 34373 -7363 se
tri 34373 -7457 34467 -7363 nw
tri 34185 -7551 34279 -7457 se
tri 34279 -7551 34373 -7457 nw
tri 34091 -7645 34185 -7551 se
tri 34185 -7645 34279 -7551 nw
tri 33997 -7739 34091 -7645 se
tri 34091 -7739 34185 -7645 nw
tri 33903 -7833 33997 -7739 se
tri 33997 -7833 34091 -7739 nw
tri 33809 -7927 33903 -7833 se
tri 33903 -7927 33997 -7833 nw
tri 33715 -8021 33809 -7927 se
tri 33809 -8021 33903 -7927 nw
tri 33621 -8115 33715 -8021 se
tri 33715 -8115 33809 -8021 nw
tri 33527 -8209 33621 -8115 se
tri 33621 -8209 33715 -8115 nw
tri 32722 -8395 32788 -8329 ne
tri 32788 -8382 32869 -8301 sw
tri 33433 -8303 33527 -8209 se
tri 33527 -8303 33621 -8209 nw
tri 33354 -8382 33433 -8303 se
rect 33433 -8382 33435 -8303
rect 32788 -8395 33435 -8382
tri 33435 -8395 33527 -8303 nw
tri 32788 -8448 32841 -8395 ne
rect 32841 -8448 33382 -8395
tri 33382 -8448 33435 -8395 nw
use sky130_fd_io__gpiov2_amux_decoder  sky130_fd_io__gpiov2_amux_decoder_0
timestamp 1676037725
transform 1 0 31774 0 1 -5388
box -341 -792 8677 3339
use sky130_fd_io__gpiov2_amux_drvr  sky130_fd_io__gpiov2_amux_drvr_0
timestamp 1676037725
transform 1 0 9862 0 1 6253
box 16159 -15244 28245 -4293
use sky130_fd_io__gpiov2_amux_ls  sky130_fd_io__gpiov2_amux_ls_0
timestamp 1676037725
transform 1 0 25054 0 1 -16031
box 1038 -423 16864 16947
<< properties >>
string GDS_END 44030200
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43961016
<< end >>
