magic
tech sky130A
magscale 1 2
timestamp 1676037725
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 361 163 642 203
rect 1 27 642 163
rect 29 -17 63 27
rect 361 21 642 27
<< locali >>
rect 108 417 346 483
rect 480 299 526 493
rect 17 215 85 265
rect 492 152 526 299
rect 480 83 526 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 299 69 527
rect 119 265 153 377
rect 197 333 281 383
rect 382 367 438 527
rect 197 299 446 333
rect 412 265 446 299
rect 119 199 266 265
rect 412 199 458 265
rect 119 181 168 199
rect 21 147 168 181
rect 412 165 446 199
rect 21 53 84 147
rect 298 131 446 165
rect 560 292 611 527
rect 118 17 264 113
rect 298 61 332 131
rect 366 17 442 97
rect 560 17 611 185
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 108 417 346 483 6 A
port 1 nsew signal input
rlabel locali s 17 215 85 265 6 B_N
port 2 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 361 21 642 27 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 29 -17 63 27 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 27 642 163 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 361 163 642 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 480 83 526 152 6 X
port 7 nsew signal output
rlabel locali s 492 152 526 299 6 X
port 7 nsew signal output
rlabel locali s 480 299 526 493 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1004888
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 999424
<< end >>
