magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< pdiff >>
rect 22593 771 22806 1297
<< locali >>
rect 18667 697 18705 731
<< viali >>
rect 18633 697 18667 731
rect 18705 697 18739 731
<< metal1 >>
tri 22870 3602 22922 3654 se
rect 22922 3602 23394 3654
rect 23446 3602 23458 3654
rect 23510 3602 23516 3654
rect 8579 3548 16095 3576
tri 22836 3568 22870 3602 se
rect 22870 3568 22888 3602
tri 22888 3568 22922 3602 nw
rect 8579 3424 8607 3548
rect 8579 3372 8585 3424
rect 8637 3372 8649 3424
rect 8701 3372 8707 3424
rect 8750 3372 8756 3424
rect 8808 3372 8820 3424
rect 8872 3372 8878 3424
rect 1961 3188 2003 3242
rect 1878 2542 1916 2592
rect 8583 2577 8619 3372
tri 8726 3348 8750 3372 se
rect 8750 3348 8793 3372
tri 8651 3273 8726 3348 se
rect 8726 3339 8793 3348
tri 8793 3339 8826 3372 nw
rect 11364 3339 11370 3391
rect 11422 3339 11434 3391
rect 11486 3358 15853 3391
rect 11486 3339 11492 3358
rect 8726 3273 8727 3339
tri 8727 3273 8793 3339 nw
tri 14707 3279 14721 3293 se
rect 14721 3279 15717 3293
rect 14707 3277 15717 3279
rect 8651 2867 8703 3273
tri 8703 3249 8727 3273 nw
rect 14707 3255 15595 3277
rect 14707 2951 14759 3255
tri 14759 3225 14789 3255 nw
tri 15575 3241 15589 3255 ne
rect 15589 3225 15595 3255
rect 15647 3225 15659 3277
rect 15711 3225 15717 3277
rect 15351 3212 15403 3218
tri 15403 3192 15422 3211 sw
rect 15403 3160 15595 3192
rect 15351 3148 15595 3160
rect 15403 3140 15595 3148
rect 15647 3140 15659 3192
rect 15711 3140 15717 3192
tri 15403 3119 15424 3140 nw
rect 15772 3128 15853 3358
rect 15351 3090 15403 3096
rect 15772 3076 15778 3128
rect 15830 3076 15842 3128
rect 15894 3076 15900 3128
rect 15772 2843 15778 2895
rect 15830 2843 15842 2895
rect 15894 2843 15900 2895
rect 8651 2803 8703 2815
rect 9220 2765 9239 2785
rect 12737 2780 12755 2800
rect 8651 2660 8703 2751
rect 8651 2608 8758 2660
rect 6259 2534 6292 2567
rect 8583 2541 8677 2577
rect 1812 2105 1851 2137
rect 5073 1350 5127 1393
rect 8641 1228 8677 2541
rect 5637 1176 5689 1223
rect 8616 1192 8677 1228
rect 8706 1219 8758 2608
rect 16067 2585 16095 3548
tri 22784 3516 22836 3568 se
tri 22836 3516 22888 3568 nw
tri 22732 3464 22784 3516 se
tri 22784 3464 22836 3516 nw
tri 22712 3444 22732 3464 se
rect 22268 3412 22732 3444
tri 22732 3412 22784 3464 nw
rect 18170 3363 18222 3369
rect 18170 3299 18222 3311
rect 18170 3241 18222 3247
rect 23347 2699 23388 2748
rect 20492 2228 20529 2255
rect 22879 1981 22916 2029
rect 23229 1983 23269 2035
rect 10372 1944 10390 1957
rect 10401 1922 10407 1974
rect 10459 1922 10473 1974
rect 10525 1922 10531 1974
rect 12382 1915 12414 1942
rect 11941 1260 11976 1292
rect 7820 1037 7860 1069
rect 8616 1062 8652 1192
rect 8706 1155 8758 1167
rect 8706 1097 8758 1103
rect 9373 1219 9425 1225
rect 9373 1155 9425 1167
rect 9425 1103 10075 1128
rect 9373 1097 10075 1103
rect 9425 1096 10075 1097
rect 8608 1056 8660 1062
rect 8608 992 8660 1004
rect 8608 934 8660 940
rect 10043 965 10075 1096
rect 10326 1019 10690 1051
rect 10326 965 10358 1019
rect 10043 933 10358 965
rect 10658 889 10690 1019
rect 17242 1004 17284 1058
rect 17596 924 17635 966
rect 10658 857 11037 889
rect 18024 864 18076 870
rect 18024 803 18076 812
tri 18076 803 18106 833 sw
rect 18024 800 18691 803
rect 18076 770 18691 800
rect 18076 751 18081 770
tri 18081 751 18100 770 nw
rect 18024 742 18076 748
tri 18595 744 18621 770 ne
rect 18621 737 18691 770
rect 18621 731 18751 737
rect 18621 697 18633 731
rect 18667 697 18705 731
rect 18739 697 18751 731
rect 18621 691 18751 697
rect 12171 335 12212 369
rect -288 -4434 -248 -4402
rect 563 -5404 595 -5362
rect -800 -5553 -782 -5528
rect -1082 -6366 -1043 -6334
rect 709 -6389 742 -6356
rect -296 -6437 -275 -6412
<< via1 >>
rect 23394 3602 23446 3654
rect 23458 3602 23510 3654
rect 8585 3372 8637 3424
rect 8649 3372 8701 3424
rect 8756 3372 8808 3424
rect 8820 3372 8872 3424
rect 11370 3339 11422 3391
rect 11434 3339 11486 3391
rect 15595 3225 15647 3277
rect 15659 3225 15711 3277
rect 15351 3160 15403 3212
rect 15351 3096 15403 3148
rect 15595 3140 15647 3192
rect 15659 3140 15711 3192
rect 15778 3076 15830 3128
rect 15842 3076 15894 3128
rect 8651 2815 8703 2867
rect 15778 2843 15830 2895
rect 15842 2843 15894 2895
rect 8651 2751 8703 2803
rect 18170 3311 18222 3363
rect 18170 3247 18222 3299
rect 10407 1922 10459 1974
rect 10473 1922 10525 1974
rect 8706 1167 8758 1219
rect 8706 1103 8758 1155
rect 9373 1167 9425 1219
rect 9373 1103 9425 1155
rect 8608 1004 8660 1056
rect 8608 940 8660 992
rect 18024 812 18076 864
rect 18024 748 18076 800
<< metal2 >>
rect 23388 3602 23394 3654
rect 23446 3602 23458 3654
rect 23510 3602 23516 3654
rect 8579 3372 8585 3424
rect 8637 3372 8649 3424
rect 8701 3372 8707 3424
rect 8750 3372 8756 3424
rect 8808 3372 8820 3424
rect 8872 3394 11310 3424
rect 8872 3372 8878 3394
tri 11248 3339 11303 3394 ne
rect 11303 3391 11310 3394
tri 11310 3391 11343 3424 sw
rect 11303 3339 11370 3391
rect 11422 3339 11434 3391
rect 11486 3339 11492 3391
rect 11532 3388 15341 3424
rect 8651 2867 8703 2873
rect 8651 2803 8703 2815
rect 8651 2745 8703 2751
rect 11532 2766 11568 3388
rect 15305 3218 15341 3388
rect 18170 3363 18222 3369
rect 18170 3299 18222 3311
rect 15589 3225 15595 3277
rect 15647 3225 15659 3277
rect 15711 3247 18170 3277
rect 15711 3241 18222 3247
rect 15711 3225 15717 3241
rect 15305 3212 15403 3218
rect 15305 3182 15351 3212
rect 15351 3148 15403 3160
rect 15589 3140 15595 3192
rect 15647 3140 15659 3192
rect 15711 3156 18310 3192
rect 15711 3140 15717 3156
rect 15351 3090 15403 3096
rect 15772 3076 15778 3128
rect 15830 3076 15842 3128
rect 15894 3076 15900 3128
rect 15772 2895 15853 3076
rect 15772 2843 15778 2895
rect 15830 2843 15842 2895
rect 15894 2843 15951 2895
tri 15907 2799 15951 2843 ne
tri 15951 2840 16006 2895 sw
rect 15951 2799 17964 2840
tri 15951 2788 15962 2799 ne
rect 15962 2788 17964 2799
rect 11532 2730 11668 2766
rect 11632 2301 11668 2730
rect 11632 2265 11732 2301
rect 10401 1922 10407 1974
rect 10459 1922 10473 1974
rect 10525 1958 10531 1974
rect 10525 1922 10746 1958
rect 10710 1661 10746 1922
rect 11696 1661 11732 2265
rect 18274 1869 18310 3156
rect 23388 2977 23516 3602
rect 10710 1625 11732 1661
rect 18032 1833 18310 1869
rect 5644 1266 5693 1311
rect 8706 1219 8758 1225
rect 8706 1155 8758 1167
rect 9373 1219 9425 1225
rect 9373 1155 9425 1167
rect 8758 1103 9373 1148
rect 8706 1097 9425 1103
rect 8608 1056 9204 1062
rect 8660 1006 9204 1056
rect 8608 992 8660 1004
rect 8608 934 8660 940
rect 18032 870 18068 1833
rect 21015 1377 21043 1404
rect 5631 828 5679 869
rect 18024 864 18076 870
rect 18024 800 18076 812
rect 18024 742 18076 748
rect 5630 656 5678 697
rect -435 -7766 -426 -7710
rect -370 -7766 -271 -7710
rect -215 -7766 -206 -7710
rect -435 -7850 -206 -7766
rect -435 -7906 -426 -7850
rect -370 -7906 -271 -7850
rect -215 -7906 -206 -7850
<< via2 >>
rect -426 -7766 -370 -7710
rect -271 -7766 -215 -7710
rect -426 -7906 -370 -7850
rect -271 -7906 -215 -7850
<< metal3 >>
rect -437 -7710 -204 -126
rect -437 -7766 -426 -7710
rect -370 -7766 -271 -7710
rect -215 -7766 -204 -7710
rect -437 -7850 -204 -7766
rect -437 -7906 -426 -7850
rect -370 -7906 -271 -7850
rect -215 -7906 -204 -7850
rect -437 -7908 -204 -7906
rect -431 -7911 -210 -7908
use sky130_fd_io__gpio_ovtv2_amux_decoder_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_decoder_i2c_fix_0
timestamp 1676037725
transform 1 0 11738 0 1 2297
box -2660 -4046 6639 1104
use sky130_fd_io__gpio_ovtv2_amux_drvr_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_drvr_i2c_fix_0
timestamp 1676037725
transform 1 0 981 0 1 558
box -262 -463 24132 3162
use sky130_fd_io__gpio_ovtv2_amux_ls_i2c_fix  sky130_fd_io__gpio_ovtv2_amux_ls_i2c_fix_0
timestamp 1676037725
transform 1 0 1902 0 1 606
box -3270 -8769 21967 3114
<< labels >>
flabel metal2 s 5630 656 5678 697 3 FreeSans 400 0 0 0 PD_CSD_VSWITCH_H
port 2 nsew
flabel metal2 s 5644 1266 5693 1311 3 FreeSans 400 0 0 0 NGA_PAD_VSWITCH_H
port 3 nsew
flabel metal2 s 5631 828 5679 869 3 FreeSans 400 0 0 0 NGA_AMX_VSWITCH_H
port 4 nsew
flabel metal2 s 21015 1377 21043 1404 3 FreeSans 400 0 0 0 HLD_I_H_N
port 5 nsew
flabel metal1 s -288 -4434 -248 -4402 3 FreeSans 400 0 0 0 VSWITCH
port 7 nsew
flabel metal1 s 1812 2105 1851 2137 3 FreeSans 400 0 0 0 VSSA
port 8 nsew
flabel metal1 s 6259 2534 6292 2567 3 FreeSans 400 90 0 0 VDDA
port 9 nsew
flabel metal1 s 23347 2699 23388 2748 3 FreeSans 400 90 0 0 PU_CSD_VDDIOQ_H_N
port 10 nsew
flabel metal1 s 22879 1981 22916 2029 3 FreeSans 400 90 0 0 PGB_PAD_VDDIOQ_H_N
port 11 nsew
flabel metal1 s 1878 2542 1916 2592 3 FreeSans 400 90 0 0 PGB_AMX_VDDA_H_N
port 12 nsew
flabel metal1 s 23229 1983 23269 2035 3 FreeSans 400 90 0 0 PGA_PAD_VDDIOQ_H_N
port 13 nsew
flabel metal1 s 1961 3188 2003 3242 3 FreeSans 400 90 0 0 PGA_AMX_VDDA_H_N
port 14 nsew
flabel metal1 s 17596 924 17635 966 3 FreeSans 400 90 0 0 D_B
port 15 nsew
flabel metal1 s 17242 1004 17284 1058 3 FreeSans 400 90 0 0 NMIDA_VCCD
port 16 nsew
flabel metal1 s 5073 1350 5127 1393 3 FreeSans 400 0 0 0 NGB_PAD_VSWITCH_H
port 17 nsew
flabel metal1 s 5637 1176 5689 1223 3 FreeSans 400 0 0 0 NGB_AMX_VSWITCH_H
port 18 nsew
flabel metal1 s 563 -5404 595 -5362 3 FreeSans 400 90 0 0 AMUX_EN_VDDA_H_N
port 19 nsew
flabel metal1 s 7820 1037 7860 1069 3 FreeSans 400 0 0 0 VSWITCH
port 7 nsew
flabel metal1 s 12171 335 12212 369 3 FreeSans 520 0 0 0 VSSD
port 20 nsew
flabel metal1 s -1082 -6366 -1043 -6334 3 FreeSans 400 0 0 0 VSSA
port 8 nsew
flabel metal1 s 20492 2228 20529 2255 3 FreeSans 400 0 0 0 VDDIO_Q
port 21 nsew
flabel metal1 s 709 -6389 742 -6356 3 FreeSans 400 0 0 0 VDDA
port 9 nsew
flabel metal1 s 11941 1260 11976 1292 3 FreeSans 400 0 0 0 VCCD
port 22 nsew
flabel metal1 s 12382 1915 12414 1942 3 FreeSans 520 0 0 0 OUT
port 23 nsew
flabel metal1 s -800 -5553 -782 -5528 3 FreeSans 400 90 0 0 ENABLE_VSWITCH_H
port 24 nsew
flabel metal1 s -296 -6437 -275 -6412 3 FreeSans 520 90 0 0 ENABLE_VDDA_H
port 25 nsew
flabel metal1 s 9220 2765 9239 2785 3 FreeSans 520 90 0 0 ANALOG_SEL
port 26 nsew
flabel metal1 s 12737 2780 12755 2800 3 FreeSans 400 90 0 0 ANALOG_POL
port 27 nsew
flabel metal1 s 10372 1944 10390 1957 3 FreeSans 400 0 0 0 ANALOG_EN
port 28 nsew
flabel comment s 16902 1461 16902 1461 0 FreeSans 1600 0 0 0 VDDA
flabel comment s 7294 1461 7294 1461 0 FreeSans 1600 0 0 0 VDDA
<< properties >>
string GDS_END 30224952
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30213802
<< end >>
