magic
tech sky130A
magscale 1 2
timestamp 1676037725
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_0
timestamp 1676037725
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_1
timestamp 1676037725
transform 1 0 1600 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_2
timestamp 1676037725
transform 1 0 3256 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 33932816
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 33931374
<< end >>
