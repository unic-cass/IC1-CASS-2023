* NGSPICE file created from wb_buttons_leds.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt wb_buttons_leds buttons clk i_wb_addr[0] i_wb_addr[10] i_wb_addr[11] i_wb_addr[12]
+ i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16] i_wb_addr[17] i_wb_addr[18]
+ i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21] i_wb_addr[22] i_wb_addr[23]
+ i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27] i_wb_addr[28] i_wb_addr[29]
+ i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3] i_wb_addr[4] i_wb_addr[5]
+ i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc i_wb_data[0] i_wb_data[10]
+ i_wb_data[11] i_wb_data[12] i_wb_data[13] i_wb_data[14] i_wb_data[15] i_wb_data[16]
+ i_wb_data[17] i_wb_data[18] i_wb_data[19] i_wb_data[1] i_wb_data[20] i_wb_data[21]
+ i_wb_data[22] i_wb_data[23] i_wb_data[24] i_wb_data[25] i_wb_data[26] i_wb_data[27]
+ i_wb_data[28] i_wb_data[29] i_wb_data[2] i_wb_data[30] i_wb_data[31] i_wb_data[3]
+ i_wb_data[4] i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8] i_wb_data[9] i_wb_stb
+ i_wb_we led_enb[0] led_enb[1] led_enb[2] led_enb[3] led_enb[4] led_enb[5] led_enb[6]
+ led_enb[7] led_enb[8] led_enb[9] leds[0] leds[10] leds[11] leds[1] leds[2] leds[3]
+ leds[4] leds[5] leds[6] leds[7] leds[8] leds[9] o_wb_ack o_wb_data[0] o_wb_data[10]
+ o_wb_data[11] o_wb_data[12] o_wb_data[13] o_wb_data[14] o_wb_data[15] o_wb_data[16]
+ o_wb_data[17] o_wb_data[18] o_wb_data[19] o_wb_data[1] o_wb_data[20] o_wb_data[21]
+ o_wb_data[22] o_wb_data[23] o_wb_data[24] o_wb_data[25] o_wb_data[26] o_wb_data[27]
+ o_wb_data[28] o_wb_data[29] o_wb_data[2] o_wb_data[30] o_wb_data[31] o_wb_data[3]
+ o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7] o_wb_data[8] o_wb_data[9] o_wb_stall
+ reset vccd1 vssd1 led_enb[11] led_enb[10]
XFILLER_0_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09671_ _05834_ _05888_ _05899_ _05910_ _05921_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a32o_1
X_18869_ clknet_4_7_0_clk _00035_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09938_ _05573_ _05649_ _06722_ _05693_ vssd1 vssd1 vccd1 vccd1 _08832_ sky130_fd_sc_hd__and4_1
X_09869_ _08060_ _08071_ _05682_ _06062_ vssd1 vssd1 vccd1 vccd1 _08082_ sky130_fd_sc_hd__and4b_1
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11900_ _01902_ _01901_ vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__nand2_1
X_12880_ _02972_ vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__clkbuf_4
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _05399_ _05355_ _00217_ _00909_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__nand4_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _04773_ _04774_ vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__xor2_2
XFILLER_0_67_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _01853_ _01854_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__xnor2_2
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13501_ _06711_ _00509_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10713_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00806_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _04608_ _04609_ _04625_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__nand3_1
XFILLER_0_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _01781_ _01782_ _01741_ _01756_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__o211ai_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16220_ _03239_ _06418_ vssd1 vssd1 vccd1 vccd1 _06589_ sky130_fd_sc_hd__or2_1
X_13432_ _03043_ _03113_ _01677_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__mux2_1
X_10644_ _00719_ _00720_ _00735_ _00736_ vssd1 vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16151_ _03126_ _06512_ _06513_ vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10575_ _07080_ cla_inst.in1\[30\] _07755_ _07047_ vssd1 vssd1 vccd1 vccd1 _00668_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _03475_ _03477_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer7 net169 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15102_ _05375_ _05376_ vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _02357_ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__inv_2
X_16082_ _03311_ _06368_ _06438_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__and3_1
X_13294_ _03396_ _03400_ _03401_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15033_ _05198_ _05202_ _05196_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__o21a_1
X_12245_ _05747_ _00878_ _02337_ _02245_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__a22oi_1
X_12176_ _02265_ _02267_ vssd1 vssd1 vccd1 vccd1 _02269_ sky130_fd_sc_hd__nand2_1
X_11127_ _00514_ _00813_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__nor2_2
X_16984_ _06874_ _06957_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__or2_1
X_11058_ ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel vssd1 vssd1 vccd1 vccd1
+ _01151_ sky130_fd_sc_hd__clkbuf_4
X_18723_ _00516_ _09183_ net69 vssd1 vssd1 vccd1 vccd1 _09249_ sky130_fd_sc_hd__a21oi_1
X_15935_ _06272_ _06280_ vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10009_ cla_inst.in2\[25\] vssd1 vssd1 vccd1 vccd1 _09352_ sky130_fd_sc_hd__buf_2
X_18654_ net62 _03086_ _09193_ vssd1 vssd1 vccd1 vccd1 _09199_ sky130_fd_sc_hd__mux2_1
X_15866_ _06157_ _06205_ _06206_ vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__or3_1
X_17605_ _08086_ _08096_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14817_ _04965_ _04966_ _05065_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__o211ai_4
X_18585_ salida\[12\] _09141_ _09142_ salida\[44\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09148_ sky130_fd_sc_hd__a221o_1
X_15797_ _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17536_ _02846_ _02847_ _08021_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__o21a_2
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14748_ _04854_ _04859_ _04852_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17467_ _06969_ net145 vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__nand2_1
X_14679_ _04750_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16418_ sel_op\[2\] sel_op\[3\] sel_op\[1\] vssd1 vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__nor3_1
X_17398_ _07869_ _07870_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16349_ _03049_ _06612_ _06728_ _06626_ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_898 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18019_ _08464_ _08545_ _08532_ vssd1 vssd1 vccd1 vccd1 _08547_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09723_ _06460_ _06482_ _05083_ _05072_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__a31oi_4
X_09654_ _05736_ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__buf_4
X_09585_ _04984_ _03750_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__and2_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10360_ _05017_ _06062_ _00451_ _00452_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__nand4_2
XFILLER_0_143_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10291_ _09240_ _09326_ _09287_ vssd1 vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__o21a_1
X_12030_ _02108_ _02121_ vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13981_ _09172_ _04154_ _00563_ _00358_ vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a22o_1
X_15720_ _05890_ _05983_ vssd1 vssd1 vccd1 vccd1 _06049_ sky130_fd_sc_hd__and2b_1
X_12932_ _01113_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__buf_2
X_15651_ _09351_ _09311_ _07744_ _02991_ vssd1 vssd1 vccd1 vccd1 _05974_ sky130_fd_sc_hd__a22o_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _02954_ _02955_ vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__and2_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _00592_ _01112_ _04773_ _04771_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__a31oi_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _08835_ _08837_ _08833_ vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__a21bo_1
X_11814_ _01906_ _01822_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15582_ _05897_ _05898_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__nor2_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _02884_ _02886_ vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17321_ _07654_ _07658_ _07785_ vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__or3b_1
X_14533_ _04756_ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__inv_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _01660_ _01662_ vssd1 vssd1 vccd1 vccd1 _01838_ sky130_fd_sc_hd__xor2_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17252_ _07113_ _06655_ _07489_ _07595_ vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__and4_1
XFILLER_0_153_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14464_ _04678_ _04680_ _04533_ _04535_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _01760_ _01761_ _01768_ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _06567_ _06570_ _00357_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13415_ _07047_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__inv_2
X_10627_ _00553_ _00542_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__and2b_1
X_17183_ _07634_ _07636_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__nand2_1
X_14395_ _04598_ _04599_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16134_ _01672_ _03188_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__or2_1
X_13346_ _03453_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__xnor2_1
X_10558_ _00646_ _00472_ _00649_ _00650_ vssd1 vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_59_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16065_ _06420_ vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ _03379_ _03380_ _03381_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10489_ _00535_ _00536_ net186 _00375_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15016_ _05262_ _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or2_1
X_12228_ _02320_ _02312_ vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _02247_ _02250_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16967_ _07399_ _07400_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__and2_1
X_18706_ _09235_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__buf_1
X_15918_ _06260_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__xor2_1
X_16898_ _07212_ _07214_ _07325_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ _06183_ _06187_ _06188_ vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__a21oi_1
X_18637_ _09176_ _09184_ vssd1 vssd1 vccd1 vccd1 _09185_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18568_ salida\[6\] _09114_ _09118_ salida\[38\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17519_ _08001_ _08002_ vssd1 vssd1 vccd1 vccd1 _08003_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18499_ _03197_ _06317_ vssd1 vssd1 vccd1 vccd1 _09067_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09706_ _06288_ _06298_ vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__nor2_1
X_09637_ ApproximateM_inst.lob_16.lob2.genblk1\[7\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05562_ sky130_fd_sc_hd__buf_2
X_09568_ _04777_ _04788_ _04799_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09499_ _03399_ vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__buf_4
X_11530_ _01185_ _01184_ _01183_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11461_ _03892_ _00180_ _00130_ _03881_ vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__a22o_1
X_13200_ _01504_ _00557_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__nand2_1
X_10412_ _00497_ _00504_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__xor2_2
X_14180_ _04369_ _04370_ vssd1 vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__and2_1
X_11392_ _01483_ _01484_ vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _04984_ _05845_ _00613_ _00612_ _00443_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a32o_1
X_10343_ _00432_ _00434_ _00433_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10274_ _00365_ _00366_ vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__nor2_2
X_13062_ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__clkbuf_4
X_12013_ _02047_ _02048_ _02049_ net328 vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__o31ai_2
X_17870_ _08383_ _08384_ vssd1 vssd1 vccd1 vccd1 _08385_ sky130_fd_sc_hd__xnor2_1
X_16821_ _07103_ _07138_ vssd1 vssd1 vccd1 vccd1 _07242_ sky130_fd_sc_hd__and2_1
X_16752_ _07165_ _07166_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__and2_1
X_13964_ _05834_ _03455_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nand2_1
X_15703_ _06028_ _06030_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__nor2_1
Xmax_cap5 _02383_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__clkbuf_1
X_12915_ _09166_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__buf_2
X_16683_ _02975_ _07089_ _07092_ _06645_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__a211o_1
X_13895_ _04058_ _04059_ vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__xor2_1
X_15634_ _05934_ _05936_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__or2_1
X_18422_ _01502_ _02891_ _02894_ vssd1 vssd1 vccd1 vccd1 _08985_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12846_ _02920_ _02938_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__or2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _03108_ _07390_ _08845_ _04668_ _07592_ vssd1 vssd1 vccd1 vccd1 _08910_ sky130_fd_sc_hd__a32o_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ _04076_ _04084_ _03536_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__mux2_1
X_12777_ _02866_ _02868_ vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__nand2_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _07767_ _07768_ vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__nor2_1
X_14516_ _04735_ _04736_ _04584_ _04704_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__a211oi_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18284_ _08833_ _08834_ vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__and2_1
X_11728_ _04416_ _00179_ _00129_ _04340_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15496_ _03537_ _03913_ _05082_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17235_ _06368_ _06438_ _06425_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__a21oi_1
X_14447_ _04480_ _04662_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11659_ _01702_ _01704_ _01750_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__nor3_1
XFILLER_0_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17166_ _07494_ _07588_ _07616_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__nor3_1
X_14378_ _02059_ _08224_ _04439_ _04437_ vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16117_ _03028_ vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__buf_4
X_13329_ _09166_ _09172_ _00218_ _00178_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__and4_1
X_17097_ _07541_ _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _06400_ _06401_ _05557_ vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17999_ _03198_ _05807_ vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09422_ op_code\[1\] vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ _05399_ _05355_ _03804_ _03914_ vssd1 vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__nand4_4
X_12700_ _02764_ _02765_ vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__xnor2_1
X_13680_ _03820_ _03822_ _03817_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__o21ai_1
X_10892_ _00981_ _00984_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _02686_ _02721_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15350_ _05452_ _05566_ vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ _02611_ _02654_ vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14301_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__nand2_2
XFILLER_0_81_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11513_ _01550_ _01561_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__or2_1
X_15281_ _05554_ _05555_ _05570_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12493_ _02585_ _02527_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__xnor2_1
Xwire133 _04284_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_1
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17020_ _00593_ _07355_ vssd1 vssd1 vccd1 vccd1 _07459_ sky130_fd_sc_hd__nor2_1
X_14232_ _04299_ _04300_ _04312_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nor3_1
XFILLER_0_135_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11444_ _04635_ _04362_ _00176_ vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14163_ _04350_ _04352_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__and2_2
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11375_ _01394_ _01413_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ _03465_ _00439_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__and2_1
X_10326_ _00417_ _00416_ _09342_ _00379_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__o211ai_2
X_14094_ _04099_ _04132_ _07962_ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__and3_1
X_18971_ clknet_4_5_0_clk _09402_ vssd1 vssd1 vccd1 vccd1 salida\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _06680_ _08441_ vssd1 vssd1 vccd1 vccd1 _08443_ sky130_fd_sc_hd__nor2_1
X_13045_ _01220_ _03136_ _03040_ vssd1 vssd1 vccd1 vccd1 _03137_ sky130_fd_sc_hd__o21a_1
X_10257_ _00348_ _00337_ _00338_ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__nand3_1
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10188_ _00278_ _00279_ _00280_ vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__nand3_1
X_17853_ _08283_ _08284_ _08282_ vssd1 vssd1 vccd1 vccd1 _08367_ sky130_fd_sc_hd__o21ai_1
X_16804_ _07215_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__xor2_1
X_17784_ _08257_ _08258_ _08291_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__a21oi_1
X_14996_ _05260_ _05261_ vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__and2_1
X_13947_ _04109_ _04115_ vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__xnor2_1
X_16735_ _07139_ _07148_ vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16666_ _02800_ _07073_ _04238_ vssd1 vssd1 vccd1 vccd1 _07074_ sky130_fd_sc_hd__a21oi_1
X_13878_ _04025_ _04026_ _04040_ vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15617_ _05861_ net118 _05937_ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__o21bai_1
X_18405_ _08912_ _08915_ vssd1 vssd1 vccd1 vccd1 _08966_ sky130_fd_sc_hd__nand2_1
X_12829_ _02903_ _02904_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__and2_2
X_16597_ _00494_ _02983_ _06487_ _06485_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__or4_2
XFILLER_0_146_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15548_ _05757_ _05861_ _05862_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__nor3_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18336_ _03206_ _08873_ _08874_ _08891_ vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__o31ai_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18267_ _08815_ _08816_ _06508_ vssd1 vssd1 vccd1 vccd1 _08817_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15479_ _05700_ _05702_ _05787_ vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17218_ _07673_ _07674_ _06649_ vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__and3b_2
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18198_ _08586_ _08668_ vssd1 vssd1 vccd1 vccd1 _08742_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17149_ _06657_ net145 vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09971_ cla_inst.in2\[30\] vssd1 vssd1 vccd1 vccd1 _09166_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ _00203_ _00134_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10111_ _00203_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__clkbuf_4
X_11091_ _05464_ _03837_ _04056_ _05508_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ _00126_ vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__inv_2
X_14850_ _03651_ _03662_ _07755_ _08169_ vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__nand4_2
Xhold85 op_code\[0\] vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__buf_1
X_13801_ _04548_ _08169_ _03953_ _03954_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__o2bb2a_1
Xhold96 net108 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _05025_ _05026_ vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__nor2_1
X_11993_ _04351_ _04373_ _07548_ _07581_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16520_ _06913_ _06914_ _04247_ vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__mux2_2
X_13732_ _03836_ _03715_ _03879_ _03880_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10944_ _01029_ _01030_ _01035_ vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16451_ _06781_ _06782_ _06780_ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__a21bo_1
X_13663_ _03802_ _03803_ _03789_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__a21o_1
X_10875_ _04001_ _00165_ _00921_ _00920_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15402_ _05575_ _05576_ _05587_ vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__and3_1
X_12614_ _02701_ _02704_ _02705_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__a211oi_1
X_16382_ _06764_ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__clkbuf_4
X_13594_ _03518_ _03521_ _03730_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18121_ _08654_ _08657_ vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__xnor2_1
X_15333_ _05574_ _05592_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__or2_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ _07036_ _07973_ _00871_ _09179_ vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__nand4_2
XFILLER_0_108_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052_ _08497_ _08530_ _08581_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__and3_1
X_15264_ _05339_ _05472_ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__and2b_1
X_12476_ _02510_ _02512_ vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__xnor2_1
X_17003_ _07438_ _07440_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__nand2_1
X_14215_ _02963_ _04404_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11427_ _03509_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__buf_4
XANTENNA_5 _00206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _05461_ _05462_ _05477_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__or3_1
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _04332_ _04333_ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _01337_ _01377_ _01440_ _01441_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _00204_ _00166_ _00260_ vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__and3_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18954_ clknet_4_1_0_clk _09415_ vssd1 vssd1 vccd1 vccd1 salida\[7\] sky130_fd_sc_hd__dfxtp_1
X_14077_ _03576_ _03579_ _03060_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__mux2_1
X_11289_ _01279_ net140 _00794_ _01381_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__o211ai_4
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _03120_ vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__buf_4
X_17905_ _02173_ _08423_ vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__nor2_1
X_18885_ clknet_4_13_0_clk _00039_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17836_ _08294_ _08312_ vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer17 _01858_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer28 net337 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17767_ _08271_ _08272_ vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__nand2_1
Xrebuffer39 _04882_ vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_1
X_14979_ _05240_ _05242_ vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xor2_2
X_16718_ _07035_ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__clkbuf_4
X_17698_ _08074_ _08076_ _08197_ vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__o21a_1
XFILLER_0_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16649_ _07053_ _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18319_ _08840_ _08841_ _08872_ vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09954_ _08681_ _08973_ _08984_ _08995_ vssd1 vssd1 vccd1 vccd1 _09005_ sky130_fd_sc_hd__nand4_4
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _08148_ _08246_ vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__xor2_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _00750_ _00751_ _00585_ _00599_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10591_ _00682_ _00683_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _00992_ _05638_ _00196_ _00871_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__and4_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12261_ _07973_ _04220_ _00774_ _07984_ vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _04014_ _04013_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__or2b_1
X_11212_ _01293_ _01294_ _01303_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__nand3_1
X_12192_ _02195_ _02198_ _02284_ vssd1 vssd1 vccd1 vccd1 _02285_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _01204_ _01233_ _01234_ _01235_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__or4_4
Xoutput75 net75 vssd1 vssd1 vccd1 vccd1 leds[3] sky130_fd_sc_hd__buf_2
Xoutput86 net86 vssd1 vssd1 vccd1 vccd1 o_wb_data[12] sky130_fd_sc_hd__clkbuf_4
Xoutput97 net97 vssd1 vssd1 vccd1 vccd1 o_wb_data[22] sky130_fd_sc_hd__clkbuf_4
X_11074_ _03728_ _00218_ _01153_ _01152_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__a31o_1
X_15951_ _06287_ vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__inv_2
X_14902_ _05141_ _05142_ _05157_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__nor3_1
X_10025_ _00105_ _00117_ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__and2_1
X_18670_ _09209_ _09210_ vssd1 vssd1 vccd1 vccd1 _09211_ sky130_fd_sc_hd__and2_1
X_15882_ _06221_ _06223_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__xnor2_1
X_17621_ _08001_ _08002_ _08004_ vssd1 vssd1 vccd1 vccd1 _08114_ sky130_fd_sc_hd__a21o_1
X_14833_ _05082_ _05084_ _03081_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__mux2_1
X_14764_ _05001_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__or2_1
X_17552_ _06421_ _08030_ _08031_ _08033_ _08038_ vssd1 vssd1 vccd1 vccd1 _08040_ sky130_fd_sc_hd__a311o_1
X_11976_ _02056_ _02066_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__xor2_1
X_13715_ _09353_ _00398_ _03705_ _03704_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__a31o_1
X_16503_ _06888_ _06896_ vssd1 vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__xor2_2
X_10927_ _00980_ _01018_ _01019_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__nor3_2
X_17483_ _07955_ _07963_ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__xnor2_1
X_14695_ _04932_ _04933_ vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nor2_2
X_13646_ _03784_ _03785_ _03606_ net324 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__a211oi_4
X_16434_ _06769_ _06821_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__or2_1
X_10858_ _04493_ _04416_ _03388_ _00949_ vssd1 vssd1 vccd1 vccd1 _00951_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _04241_ _06739_ _06746_ _03117_ vssd1 vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__a211o_1
X_13577_ _03700_ _03711_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10789_ _00877_ _00881_ vssd1 vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__nand2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _05607_ _05610_ vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18104_ _07604_ _07623_ _08638_ vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12528_ _02540_ _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__and2_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16296_ _00494_ _06509_ _06427_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15247_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ _08563_ _08564_ vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12459_ _07243_ _00145_ _00129_ _07221_ vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__a22o_1
X_15178_ _05364_ vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14129_ _04123_ _04145_ _04313_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__o211a_2
X_18937_ clknet_4_3_0_clk _00091_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[23\] sky130_fd_sc_hd__dfxtp_1
X_09670_ _04591_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__buf_6
X_18868_ clknet_4_5_0_clk _00034_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__dfxtp_1
X_17819_ _03041_ _06511_ _02985_ vssd1 vssd1 vccd1 vccd1 _08330_ sky130_fd_sc_hd__and3b_1
X_18799_ _09308_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09937_ _08800_ _08811_ vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__xor2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _08039_ _06613_ _08049_ _06019_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09799_ _07210_ _07297_ _07308_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__nand3_4
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11830_ _06591_ _00774_ _00909_ _00806_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__a22o_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11761_ _01657_ _01656_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__and2b_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _03625_ _03626_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _00803_ _00804_ vssd1 vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__xor2_2
XFILLER_0_49_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _04628_ _04629_ _04674_ _04675_ vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__and4bb_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11692_ _01742_ _01753_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__and2_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13431_ _03105_ _03110_ _03048_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__mux2_1
X_10643_ _00733_ _00734_ _00721_ _00722_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_153_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ _01113_ _06509_ _09354_ vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13362_ _01504_ _00716_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10574_ _06711_ _07384_ _00478_ _00319_ _08158_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__a32o_1
Xrebuffer8 _03781_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_1
X_15101_ _01745_ _03067_ vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12313_ _02402_ _02404_ vssd1 vssd1 vccd1 vccd1 _02406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16081_ _00558_ _06437_ vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__and2_1
X_13293_ _04558_ _07962_ _03397_ _03398_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__a22o_1
X_15032_ _05299_ _05300_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__or2_1
X_12244_ _02244_ vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ _02265_ _02267_ vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__or2_4
X_11126_ _01132_ _01205_ _01216_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__a21oi_2
X_16983_ _07416_ _07418_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__nand2_1
X_18722_ _09247_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__clkbuf_1
X_11057_ _01037_ _01036_ _01028_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__a21o_1
X_15934_ _06278_ _06279_ vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__nand2_1
X_10008_ _09350_ vssd1 vssd1 vccd1 vccd1 _09351_ sky130_fd_sc_hd__clkbuf_4
X_18653_ _09198_ vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__buf_1
X_15865_ _06037_ _06163_ _02992_ _05652_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__o211a_1
X_17604_ _08087_ _08095_ vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14816_ _05063_ _05064_ _04967_ _04928_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a211o_1
X_18584_ net293 _09140_ _09147_ _09144_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__o211a_1
X_15796_ _06086_ _06130_ vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17535_ _02846_ _02847_ _04238_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__a21oi_1
X_14747_ _04845_ _04988_ _04986_ _04987_ vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__o211ai_4
X_11959_ _02042_ _02050_ _02027_ _02051_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_129_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14678_ _04906_ _04914_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17466_ _07943_ _07944_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13629_ _03761_ _03762_ _03767_ vssd1 vssd1 vccd1 vccd1 _03768_ sky130_fd_sc_hd__nand3_1
X_16417_ _04340_ _04362_ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17397_ _06875_ _07314_ vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16348_ _02982_ _06619_ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16279_ _06652_ vssd1 vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18018_ _08464_ _08532_ _08545_ vssd1 vssd1 vccd1 vccd1 _08546_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09722_ _06471_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09653_ _05682_ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09584_ _03717_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__buf_6
XFILLER_0_89_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10290_ _07624_ _00240_ _00382_ vssd1 vssd1 vccd1 vccd1 _00383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_131_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13980_ _09166_ _09172_ _04154_ _00563_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__and4_1
X_12931_ _03023_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__buf_2
X_15650_ _03015_ _03142_ _05884_ _05883_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__a31o_1
X_12862_ _00904_ _02953_ _02952_ _02945_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__o211ai_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _04822_ _04824_ _04830_ vssd1 vssd1 vccd1 vccd1 _09356_ sky130_fd_sc_hd__a21bo_1
X_11813_ _01823_ _01821_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__or2_1
X_15581_ _09351_ _07744_ _05896_ vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__and3_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _02873_ _02877_ _02885_ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__a21oi_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _04741_ _04742_ _04753_ vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__nand3_2
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _07654_ _07658_ _07785_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__o21ba_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _01835_ _01832_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _04533_ _04535_ _04678_ _04680_ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a211oi_2
X_17251_ _07707_ _07709_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__nand2_1
X_11675_ _01766_ _01767_ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__xnor2_1
X_16202_ _06532_ _06568_ vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__nor2_2
X_13414_ _02977_ _00494_ _03533_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__or3_2
XFILLER_0_153_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10626_ _00543_ _00552_ vssd1 vssd1 vccd1 vccd1 _00719_ sky130_fd_sc_hd__and2_1
X_17182_ _07630_ _07332_ _07632_ _07633_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__o22ai_1
X_14394_ _04603_ _04604_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16133_ _01863_ _03186_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13345_ _02972_ _03456_ _03457_ vssd1 vssd1 vccd1 vccd1 _03458_ sky130_fd_sc_hd__and3_1
X_10557_ _05834_ _07123_ _00647_ _00648_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _02965_ _06418_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13276_ _03379_ _03380_ _03381_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__nand3_1
XFILLER_0_110_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10488_ _00578_ _00579_ _00396_ _00538_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__o211a_1
X_15015_ _05262_ _05282_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12227_ _02313_ _02319_ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__xnor2_1
X_12158_ _02247_ _02250_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__xor2_1
X_11109_ _01051_ _01052_ _01039_ _01050_ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a211oi_1
X_12089_ _02178_ _02181_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__or2_1
X_16966_ _06766_ _07106_ _07398_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__o21ai_1
X_18705_ _09209_ _09234_ vssd1 vssd1 vccd1 vccd1 _09235_ sky130_fd_sc_hd__and2_1
X_15917_ _06219_ _06261_ vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__nand2_1
X_16897_ _07215_ _07223_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__or2_1
X_18636_ net35 _03029_ _09183_ vssd1 vssd1 vccd1 vccd1 _09184_ sky130_fd_sc_hd__mux2_1
X_15848_ _06183_ _06187_ _03202_ vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18567_ net252 _09098_ _09134_ _09126_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15779_ _06111_ _06112_ vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _07860_ _07865_ _07862_ vssd1 vssd1 vccd1 vccd1 _08002_ sky130_fd_sc_hd__a21bo_1
X_18498_ _06413_ _07274_ _09065_ _06720_ vssd1 vssd1 vccd1 vccd1 _09066_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17449_ _06426_ _06441_ _07916_ _07924_ _07926_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__o311a_1
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09705_ _04088_ _03892_ _04395_ _04886_ vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09636_ _05442_ _05540_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__xnor2_2
X_09567_ _03509_ _03914_ _03476_ _03531_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09498_ _03837_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _04088_ _04121_ _00180_ _00130_ vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _00501_ _00503_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__xnor2_2
X_11391_ _01473_ _01482_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13130_ _00625_ _00626_ vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__nand2_1
X_10342_ _00432_ _00433_ _00434_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__nand3_1
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13061_ _00665_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__clkbuf_4
X_10273_ _00355_ _00356_ _00364_ vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12012_ _02103_ _02104_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__and2b_1
X_16820_ _07103_ _07138_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__or2_1
X_16751_ _00214_ _06673_ _02533_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__or3b_1
X_13963_ _04131_ _04133_ vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__nor2_1
X_15702_ _06024_ _06027_ vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__nor2_1
Xmax_cap6 _03753_ vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__buf_1
X_12914_ _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__buf_2
X_13894_ net119 _03893_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__nor2_2
X_16682_ _03921_ _07090_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18421_ _08981_ _08982_ vssd1 vssd1 vccd1 vccd1 _08983_ sky130_fd_sc_hd__xnor2_1
X_15633_ _05924_ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__inv_2
X_12845_ _02936_ _02937_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__or2b_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _08906_ _08907_ vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _02866_ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__or2_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ _05804_ _05623_ _05807_ _03125_ _05880_ vssd1 vssd1 vccd1 vccd1 _09367_ sky130_fd_sc_hd__a221o_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _07735_ _07765_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__and2_1
X_14515_ _04584_ _04704_ _04735_ _04736_ vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__o211a_4
X_11727_ _01816_ _01819_ vssd1 vssd1 vccd1 vccd1 _01820_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18283_ _03143_ _08428_ _01417_ vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__or3b_1
X_15495_ _05084_ _05088_ _03081_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17234_ _06484_ _07688_ _07689_ _07692_ _06462_ vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__a311o_1
XFILLER_0_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14446_ _04653_ _04661_ vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__xnor2_1
X_11658_ _01702_ _01704_ _01750_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ _00183_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14377_ _04451_ _04452_ vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17165_ _07494_ _07588_ _07616_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11589_ _05682_ _08409_ _01578_ _01577_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13328_ _03005_ _01264_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16116_ _03050_ _02607_ _03170_ _06470_ _06475_ vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__o311a_1
X_17096_ _07539_ _07426_ _07540_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ _03202_ _03362_ _03363_ vssd1 vssd1 vccd1 vccd1 _03364_ sky130_fd_sc_hd__and3_1
X_16047_ _01359_ _03056_ vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17998_ _06915_ _08141_ _08524_ _06721_ vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__o211a_1
X_16949_ _07333_ _07334_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__or2b_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _03195_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18619_ net269 _09157_ _09170_ _09162_ vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960_ _01039_ _01050_ _01051_ _01052_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09619_ _05355_ vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__buf_6
X_10891_ _00982_ _00983_ vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12630_ _07711_ _00193_ _02685_ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _02643_ _02652_ _02613_ _02653_ vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_109_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14300_ _04500_ _04499_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__or2b_1
X_11512_ _01551_ _01560_ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15280_ _05554_ _05555_ _05570_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12492_ _02460_ _02472_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ _04332_ _04333_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__or2b_1
X_11443_ _04362_ _00176_ _00145_ _04635_ vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire145 _07389_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
XFILLER_0_22_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14162_ _04338_ _04183_ _04349_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__nand3_1
X_11374_ _01465_ _01464_ _01462_ vssd1 vssd1 vccd1 vccd1 _01467_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ _03629_ _03596_ _05039_ _04460_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__nand4_2
X_10325_ _00379_ _09342_ _00416_ _00417_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a211o_2
XFILLER_0_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14093_ _04273_ _04275_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__or2b_1
X_18970_ clknet_4_4_0_clk _09401_ vssd1 vssd1 vccd1 vccd1 salida\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _06390_ _06790_ _08440_ _04336_ vssd1 vssd1 vccd1 vccd1 _08441_ sky130_fd_sc_hd__a22o_1
X_13044_ _03028_ _01136_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__nor2_1
X_10256_ _00337_ _00338_ _00348_ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__a21o_2
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ _08363_ _08364_ vssd1 vssd1 vccd1 vccd1 _08366_ sky130_fd_sc_hd__nand2_1
X_10187_ _08344_ _08354_ _08333_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__a21bo_1
X_16803_ _07220_ _07222_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__xnor2_1
X_17783_ _08277_ _08290_ vssd1 vssd1 vccd1 vccd1 _08291_ sky130_fd_sc_hd__xnor2_1
X_14995_ _05244_ _05245_ _05259_ vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16734_ _07146_ _07147_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__and2_1
X_13946_ _04113_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16665_ _02798_ _02830_ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__or2b_1
X_13877_ _04028_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18404_ _08964_ vssd1 vssd1 vccd1 vccd1 _08965_ sky130_fd_sc_hd__buf_1
X_15616_ _05934_ _05936_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12828_ _00592_ _00214_ _00886_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__and3_1
X_16596_ _06703_ _06707_ _06709_ _06715_ _03062_ _03081_ vssd1 vssd1 vccd1 vccd1 _06998_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18335_ _08880_ _08886_ _08890_ vssd1 vssd1 vccd1 vccd1 _08891_ sky130_fd_sc_hd__and3b_1
X_15547_ _05859_ _05860_ _05771_ _05808_ vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__o211a_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _01239_ _01246_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18266_ _08752_ _08754_ _08751_ vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__a21o_1
X_15478_ _05703_ _05706_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17217_ _07669_ _07670_ _07672_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__or3_1
XFILLER_0_142_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14429_ _04641_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__or2_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18197_ _08739_ _08740_ vssd1 vssd1 vccd1 vccd1 _08741_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17148_ _07594_ _07597_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09970_ _09145_ _09037_ _09048_ vssd1 vssd1 vccd1 vccd1 _09158_ sky130_fd_sc_hd__and3_1
X_17079_ _07521_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10110_ cla_inst.in2\[21\] vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__clkbuf_4
X_11090_ _05213_ _04864_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__and2_1
X_10041_ _00132_ vssd1 vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__buf_4
Xsplit9 _03366_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_8
X_13800_ _03953_ _03954_ _04548_ _07374_ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__and4bb_1
Xhold86 salida\[0\] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold97 _00007_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _05023_ _05024_ _05019_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__a21oi_1
X_11992_ _04690_ _00127_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__nand2_1
X_13731_ _03877_ _03878_ _03667_ _03838_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10943_ _01029_ _01030_ _01035_ vssd1 vssd1 vccd1 vccd1 _01036_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16450_ _02972_ _06837_ _06838_ vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13662_ _03789_ _03802_ _03803_ vssd1 vssd1 vccd1 vccd1 _03805_ sky130_fd_sc_hd__nand3_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10874_ _00918_ net190 _00966_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15401_ _05700_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_ sky130_fd_sc_hd__xnor2_1
X_12613_ _02664_ _02663_ _02658_ vssd1 vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__a21oi_1
X_13593_ _03727_ _03729_ vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__nand2_1
X_16381_ _06758_ _06761_ _00132_ vssd1 vssd1 vccd1 vccd1 _06764_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_94_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18120_ _08655_ _08656_ vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__or2_1
X_15332_ _05604_ _05605_ _05610_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__or3b_1
X_12544_ _07243_ _01031_ _09179_ _07221_ vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18051_ _08497_ _08530_ _08581_ vssd1 vssd1 vccd1 vccd1 _08582_ sky130_fd_sc_hd__a21oi_2
X_15263_ _05480_ _05496_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__or2_1
X_12475_ _02482_ _02532_ _02567_ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17002_ _06749_ _07216_ _07437_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__a21o_1
X_11426_ _03574_ _03662_ _09188_ _07591_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__and4_1
X_14214_ _04068_ _04070_ _04236_ _04405_ _04408_ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__o311a_1
X_15194_ _05461_ _05462_ _05477_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__o21ai_2
XANTENNA_6 _00309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14145_ _04146_ _04167_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__or2b_1
X_11357_ _01448_ _01446_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__or3_4
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10308_ _00258_ _00259_ vssd1 vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__and2_1
X_18953_ clknet_4_1_0_clk _09414_ vssd1 vssd1 vccd1 vccd1 salida\[6\] sky130_fd_sc_hd__dfxtp_1
X_14076_ _03537_ _04256_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__and2_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _00779_ _00793_ _00792_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__a21o_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__buf_2
X_17904_ _02846_ _02850_ _02469_ vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__a21oi_2
X_10239_ _00303_ _00304_ _08529_ _08659_ vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__a211o_1
X_18884_ clknet_4_8_0_clk _00038_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_17835_ _08316_ _08317_ vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__nand2_1
Xrebuffer18 net332 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17766_ _08266_ _08270_ vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__nand2_1
X_14978_ _05121_ _05122_ _05241_ vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__o21ai_2
Xrebuffer29 net216 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_1
X_16717_ _07127_ _07128_ vssd1 vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__and2b_1
X_13929_ _03574_ _08757_ _04093_ _04094_ vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__o2bb2a_1
X_17697_ _08188_ _08196_ vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ _07050_ _07052_ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ _06976_ _06978_ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18318_ _08870_ _08871_ vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__xor2_1
XFILLER_0_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18249_ _08716_ _08722_ _08720_ vssd1 vssd1 vccd1 vccd1 _08797_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09953_ _08659_ _08670_ _06373_ _08322_ vssd1 vssd1 vccd1 vccd1 _08995_ sky130_fd_sc_hd__o211ai_4
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _08202_ _08213_ _08235_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__or3_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10590_ _00362_ _00223_ _00680_ _00681_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12260_ _02243_ _02251_ vssd1 vssd1 vccd1 vccd1 _02353_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11211_ _01293_ _01294_ _01303_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__a21o_1
X_12191_ _02132_ _02283_ vssd1 vssd1 vccd1 vccd1 _02284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ _01077_ _01203_ _01181_ _01201_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput76 net76 vssd1 vssd1 vccd1 vccd1 leds[4] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 vssd1 vssd1 vccd1 vccd1 o_wb_data[13] sky130_fd_sc_hd__clkbuf_4
X_11073_ _01149_ _01150_ _01165_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__and3_2
X_15950_ _04823_ _06289_ _06290_ _06291_ _06296_ vssd1 vssd1 vccd1 vccd1 _09375_ sky130_fd_sc_hd__a32o_1
Xoutput98 net98 vssd1 vssd1 vccd1 vccd1 o_wb_data[23] sky130_fd_sc_hd__clkbuf_4
X_14901_ _05141_ _05142_ _05157_ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__o21a_1
X_10024_ _00114_ _00116_ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__nor2_1
X_15881_ _06178_ _06222_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__or2_1
X_17620_ _08111_ _08112_ vssd1 vssd1 vccd1 vccd1 _08113_ sky130_fd_sc_hd__xor2_1
X_14832_ _03097_ _03106_ _03062_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17551_ _06462_ _08035_ _08037_ vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__or3b_1
X_14763_ _05004_ _05007_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__or2_1
X_11975_ _02027_ _02051_ _02042_ _02050_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16502_ _06893_ _06894_ vssd1 vssd1 vccd1 vccd1 _06896_ sky130_fd_sc_hd__xnor2_2
X_13714_ _03653_ _03659_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__or2_1
X_10926_ _00978_ _00979_ net195 _00955_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__a211oi_2
X_17482_ _07956_ _07961_ vssd1 vssd1 vccd1 vccd1 _07963_ sky130_fd_sc_hd__xnor2_1
X_14694_ _04758_ _04803_ _04931_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__and3_1
X_16433_ _06800_ _06820_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__xor2_1
X_13645_ _03606_ _03753_ _03784_ _03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__o211a_2
XFILLER_0_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10857_ _04416_ _03399_ _00949_ _04493_ vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _03916_ _06745_ vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__nor2_1
X_13576_ _03447_ _03710_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__xor2_1
X_10788_ _00207_ vssd1 vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__buf_4
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _07604_ _07623_ _08638_ vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__and3_1
X_15315_ _05608_ _05609_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__nand2_1
X_12527_ _02538_ _02539_ vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16295_ _06649_ _06669_ _06670_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18034_ _08469_ _08480_ _08468_ vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15246_ _05532_ _05533_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__nor2_1
X_12458_ _07984_ _07973_ _00145_ _00196_ vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__nand4_2
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11409_ _01501_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15177_ _05457_ _05458_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__nor2_1
X_12389_ _02479_ _02481_ vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__and2_1
X_14128_ _04299_ _04300_ _04312_ vssd1 vssd1 vccd1 vccd1 _04314_ sky130_fd_sc_hd__o21ai_2
X_18936_ clknet_4_2_0_clk _00090_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[22\] sky130_fd_sc_hd__dfxtp_1
X_14059_ _04065_ _04072_ _04236_ _04238_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__a31o_1
X_18867_ clknet_4_7_0_clk net304 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__dfxtp_1
X_17818_ _02985_ _06511_ _01695_ vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18798_ _09298_ _09307_ vssd1 vssd1 vccd1 vccd1 _09308_ sky130_fd_sc_hd__and2_1
XFILLER_0_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17749_ _08212_ _08211_ vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09936_ _05834_ _06094_ _06624_ _06602_ vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _06019_ _08039_ _06613_ _08049_ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__and4_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _07178_ _07199_ _07189_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__a21o_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _06971_ _04460_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__nand2_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _08452_ _05910_ _05899_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a21bo_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__inv_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10642_ _00721_ _00722_ _00733_ _00734_ vssd1 vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__a211o_2
X_13430_ _03549_ _03550_ _02489_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13361_ _03473_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10573_ _06993_ _00665_ _00501_ _00500_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15100_ _05373_ _05374_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__xor2_1
Xrebuffer9 _03810_ vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlymetal6s2s_1
X_12312_ _02402_ _02404_ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__nand2_1
X_13292_ _04558_ _06732_ _03397_ _03398_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__nand4_1
X_16080_ _00593_ _00248_ _06436_ vssd1 vssd1 vccd1 vccd1 _06437_ sky130_fd_sc_hd__and3_1
X_15031_ _05188_ _05206_ _05298_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__a21oi_1
X_12243_ _02208_ _02331_ _02335_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12174_ _02234_ _02239_ _02266_ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__a21oi_2
X_11125_ _01217_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__inv_2
X_16982_ _06968_ _06946_ _07026_ _06890_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__a22o_1
X_18721_ _09245_ _09246_ vssd1 vssd1 vccd1 vccd1 _09247_ sky130_fd_sc_hd__and2_1
X_11056_ _01037_ _01028_ _01036_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__nand3_1
X_15933_ _06273_ _06276_ vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__nand2_1
X_10007_ _09349_ vssd1 vssd1 vccd1 vccd1 _09350_ sky130_fd_sc_hd__clkbuf_4
X_18652_ _09176_ _09196_ vssd1 vssd1 vccd1 vccd1 _09198_ sky130_fd_sc_hd__and2_1
X_15864_ _06155_ _06204_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__xnor2_1
X_17603_ _08092_ _08094_ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__xnor2_1
X_14815_ _04967_ _04928_ _05063_ _05064_ vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_59_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18583_ salida\[11\] _09141_ _09142_ salida\[43\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09147_ sky130_fd_sc_hd__a221o_1
X_15795_ _06086_ _06130_ vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17534_ _08016_ _08018_ _08019_ vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__a21oi_1
X_14746_ _04986_ _04987_ _04845_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__a211o_1
X_11958_ _02009_ _02024_ _02026_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _05355_ _04384_ _04471_ _05399_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__a22o_1
X_17465_ _02347_ _06891_ vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__nand2_1
X_14677_ _04907_ _04913_ vssd1 vssd1 vccd1 vccd1 _04914_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11889_ _01868_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__xor2_1
X_16416_ _05213_ _03003_ _03004_ _06523_ vssd1 vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13628_ _03765_ _03766_ vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__xor2_2
XFILLER_0_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17396_ _07867_ _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16347_ _06724_ _06726_ _03061_ vssd1 vssd1 vccd1 vccd1 _06727_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13559_ _03689_ _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16278_ _06427_ _06651_ vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18017_ _08537_ _08544_ vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__xor2_1
X_15229_ _05426_ _05427_ _05515_ vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__o21a_1
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09721_ _05497_ vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__buf_6
X_18919_ clknet_4_8_0_clk _00073_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09652_ _05627_ _05660_ _05682_ _05715_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__and4b_1
XFILLER_0_78_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _04941_ _04952_ _04962_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__nand3_2
XFILLER_0_145_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold150 salida\[3\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_1
XFILLER_0_130_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09919_ _08615_ _05888_ _06417_ _06406_ vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__a31o_1
X_12930_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _02945_ _02952_ _02953_ _00904_ vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__a211o_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _02976_ _03038_ _04826_ _04829_ _03121_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__o32a_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _04132_ _04984_ _07559_ _07602_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__nand4_4
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _09351_ _07744_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__a21oi_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _02876_ _02875_ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__and2b_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14531_ _04741_ _04742_ _04753_ vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__a21oi_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _01832_ _01835_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__and2b_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17250_ _06756_ _07410_ _07708_ _06542_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14462_ _04676_ _04677_ _04566_ _04538_ vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ _01722_ _01723_ _01724_ _01732_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__a31o_1
X_16201_ _00210_ _06528_ _06530_ _06533_ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__or4_4
X_13413_ _03032_ _03085_ _03089_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10625_ _00714_ _00717_ vssd1 vssd1 vccd1 vccd1 _00718_ sky130_fd_sc_hd__xor2_2
X_17181_ _07630_ _07126_ _07632_ _07633_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__or4_1
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14393_ _04304_ _04600_ _04601_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16132_ _06488_ _06492_ _03061_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__mux2_1
X_10556_ _05834_ _08876_ _00647_ _00648_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__nand4_2
X_13344_ _07091_ _00513_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _03292_ _03217_ vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10487_ _00396_ _00538_ _00578_ _00579_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a211oi_2
X_13275_ _03207_ _03209_ _03208_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _05281_ vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__inv_2
X_12226_ _02317_ _02318_ vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__nor2_1
X_12157_ _02248_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__xnor2_2
X_11108_ _01181_ _01198_ _01199_ _01200_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__nand4_2
X_12088_ _08713_ _00147_ _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and4_1
X_16965_ _06766_ _07106_ _07398_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__or3_1
X_11039_ _01126_ _01130_ _01131_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__nand3_1
X_18704_ net52 _03056_ _09182_ vssd1 vssd1 vccd1 vccd1 _09234_ sky130_fd_sc_hd__mux2_1
X_15916_ _06178_ _06221_ vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nand2_1
X_16896_ _07322_ _07323_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__nand2_1
X_18635_ _09182_ vssd1 vssd1 vccd1 vccd1 _09183_ sky130_fd_sc_hd__buf_2
X_15847_ _06184_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and2_1
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ salida\[5\] _09114_ _09118_ salida\[37\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09134_ sky130_fd_sc_hd__a221o_1
X_15778_ _06032_ _06110_ vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17517_ _07855_ _07876_ _08000_ vssd1 vssd1 vccd1 vccd1 _08001_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14729_ _01520_ _07722_ _07406_ _03651_ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18497_ _03155_ _09064_ vssd1 vssd1 vccd1 vccd1 _09065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17448_ _06376_ _06372_ _06375_ _06598_ _07925_ vssd1 vssd1 vccd1 vccd1 _07926_ sky130_fd_sc_hd__a311o_1
X_17379_ _07840_ _07849_ vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09704_ _04121_ _04395_ _04657_ _04088_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__a22oi_2
X_09635_ _05475_ _05529_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09566_ _03465_ _03410_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09497_ _03793_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__buf_8
XFILLER_0_93_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _07363_ _00502_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ _01473_ _01482_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10341_ _03377_ _04384_ _04886_ _03356_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__a22o_1
X_13060_ _01677_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__clkbuf_4
X_10272_ _00355_ _00356_ _00364_ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12011_ _02088_ _02089_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__xor2_1
X_16750_ _02533_ _06510_ _00214_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a21bo_1
X_13962_ _05453_ _00645_ _00502_ _09248_ vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15701_ _06024_ _06027_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__and2_1
X_12913_ _03005_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__clkbuf_4
Xmax_cap7 _01329_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_1
X_16681_ _06741_ _06736_ _06738_ _06731_ _03912_ _03077_ vssd1 vssd1 vccd1 vccd1 _07090_
+ sky130_fd_sc_hd__mux4_2
X_13893_ _04055_ _04057_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__nand2_2
X_18420_ _08926_ _08928_ _08925_ vssd1 vssd1 vccd1 vccd1 _08982_ sky130_fd_sc_hd__a21o_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15632_ _04080_ _05623_ _05881_ _03125_ _05953_ vssd1 vssd1 vccd1 vccd1 _09368_ sky130_fd_sc_hd__a221o_1
X_12844_ _02913_ _02935_ _02934_ _02933_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _08903_ _08905_ vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__nand2_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15563_ _05875_ _05877_ _05879_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__a21oi_2
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _02867_ _01808_ vssd1 vssd1 vccd1 vccd1 _02868_ sky130_fd_sc_hd__nor2_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17302_ _07735_ _07765_ vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__nor2_1
X_14514_ _04723_ _04724_ _04734_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__or3_4
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18282_ _01417_ _06512_ _03143_ vssd1 vssd1 vccd1 vccd1 _08833_ sky130_fd_sc_hd__a21bo_1
X_11726_ _01817_ _01818_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__xor2_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15494_ _05803_ _03918_ _03547_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17233_ _06369_ _06790_ _07691_ _06368_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__a22o_1
X_14445_ _04654_ _04660_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11657_ _01748_ _01749_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _00562_ _00570_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__or2b_1
X_17164_ _07603_ net238 vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__xor2_1
X_14376_ _04581_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__a21oi_1
X_11588_ _01670_ _01676_ _01679_ _01680_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16115_ _03027_ _03166_ _02685_ _02983_ vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__a211o_1
X_13327_ _03258_ _03261_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10539_ _00620_ _00621_ _00631_ vssd1 vssd1 vccd1 vccd1 _00632_ sky130_fd_sc_hd__o21ai_2
X_17095_ _07539_ _07426_ _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16046_ _06398_ _06399_ _05368_ vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__a21o_1
X_13258_ _03358_ _03361_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12209_ _02290_ net322 _02151_ _02301_ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__o211a_4
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13189_ _03278_ _03288_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17997_ _06392_ _06546_ _08523_ _00813_ vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__o2bb2a_1
X_16948_ _07342_ _07343_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__or2b_1
X_16879_ _07301_ _07304_ vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__nor2_1
X_09420_ op_code\[2\] op_code\[3\] vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nand2_4
X_18618_ salida\[26\] _09159_ _09160_ salida\[58\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09170_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18549_ _09115_ net27 net1 vssd1 vssd1 vccd1 vccd1 _09120_ sky130_fd_sc_hd__or3b_1
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _05290_ vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__buf_8
XFILLER_0_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10890_ _05290_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel _03739_
+ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _00983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ _04558_ _04591_ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12560_ _02605_ _02606_ _02612_ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11511_ _01564_ _01601_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__nand4_2
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12491_ _02531_ _02583_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__nor2_1
X_14230_ _04161_ _04335_ _04378_ _04379_ vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__a211o_1
XFILLER_0_151_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11442_ _01533_ _01534_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__or2_1
Xwire146 _07216_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XFILLER_0_123_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11373_ _01462_ _01464_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__nand3b_4
X_14161_ _04338_ _04183_ _04349_ vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13112_ _03377_ _05039_ _04384_ _03356_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__a22o_1
X_10324_ _00396_ _00397_ _00415_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__and3_1
X_14092_ _04271_ _04272_ net174 _04095_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__a211o_1
X_10255_ _00340_ _00347_ vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _03368_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__a21o_1
X_13043_ _01672_ _03134_ _03040_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o21a_1
X_17851_ _08349_ _08350_ _08362_ vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__nand3_1
X_10186_ _00275_ _00277_ _00276_ vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__a21o_1
X_16802_ _06579_ _07126_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__or2_1
X_17782_ _08287_ _08288_ vssd1 vssd1 vccd1 vccd1 _08290_ sky130_fd_sc_hd__nor2_1
X_14994_ _05244_ _05245_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__o21ai_1
X_16733_ _07142_ _07144_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__nand2_1
X_13945_ _04690_ _07722_ _04111_ _04112_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__o2bb2a_1
X_16664_ _03206_ _07071_ vssd1 vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__nor2_1
X_13876_ _03823_ _04038_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__xor2_1
X_15615_ _05935_ _05860_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__nor2_1
X_18403_ _08961_ _08963_ vssd1 vssd1 vccd1 vccd1 _08964_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12827_ _02918_ _02919_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__nand2_1
X_16595_ _06343_ _06345_ _06995_ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__nand3_1
X_18334_ _08888_ _06402_ _06403_ _07084_ _08889_ vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__a311o_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15546_ _05771_ _05808_ _05859_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__a211oi_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _02176_ _02846_ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__and3_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18265_ _08813_ _08814_ vssd1 vssd1 vccd1 vccd1 _08815_ sky130_fd_sc_hd__nor2_1
X_11709_ _01771_ _01781_ _01800_ _01801_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15477_ _05784_ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ _02713_ _02781_ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__nor2_1
X_17216_ _07669_ _07670_ _07672_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__o21a_1
X_14428_ _04630_ _04640_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__and2_1
X_18196_ _08696_ _08738_ vssd1 vssd1 vccd1 vccd1 _08740_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17147_ _06542_ _07113_ _07489_ _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__and4_1
XFILLER_0_142_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14359_ _04315_ _04331_ _04487_ _04488_ vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17078_ _06875_ _07035_ vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16029_ _02988_ _03111_ vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _00126_ _00128_ _00106_ _00132_ vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__and4b_1
Xhold87 net109 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _04438_ _09188_ _07591_ _04646_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold98 net111 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _03667_ _03838_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__o211a_1
X_10942_ _01032_ _01033_ _01034_ vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13661_ _03800_ _03801_ _03794_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10873_ _00961_ _00965_ vssd1 vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15400_ _05600_ _05601_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12612_ _02664_ _02658_ _02663_ vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__and3_1
X_16380_ net237 _06579_ _06657_ _06762_ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__and4bb_1
X_13592_ _03724_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _05503_ _05506_ _05603_ vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12543_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _00196_ vssd1
+ vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__and2_1
X_18050_ _08578_ _08580_ vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15262_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ _02542_ _02566_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17001_ _06665_ _07318_ _07437_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__or3b_1
X_14213_ _04233_ _04235_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a21boi_1
X_11425_ _01516_ _01517_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15193_ _05473_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__xnor2_1
XANTENNA_7 _00443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ _04330_ _04331_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ _01444_ _01445_ _01370_ _01374_ vssd1 vssd1 vccd1 vccd1 _01449_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _00164_ _00399_ vssd1 vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18952_ clknet_4_1_0_clk _09413_ vssd1 vssd1 vccd1 vccd1 salida\[5\] sky130_fd_sc_hd__dfxtp_1
X_14075_ _03912_ _04254_ _04255_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__o21ai_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _01279_ _01286_ _01287_ vssd1 vssd1 vccd1 vccd1 _01380_ sky130_fd_sc_hd__nor3_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17903_ _08413_ _08418_ _08421_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__a21oi_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _06765_ _03037_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__nand2_2
X_10238_ _00326_ _00327_ _00329_ vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__nand3_4
X_18883_ clknet_4_9_0_clk _00037_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_10169_ _00250_ _00251_ _00261_ vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__o21ai_1
X_17834_ _03041_ _06464_ net116 _08346_ vssd1 vssd1 vccd1 vccd1 _09396_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ _05123_ _05134_ vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__or2b_1
X_17765_ _08266_ _08270_ vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__or2_1
Xrebuffer19 _01849_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_1
X_13928_ _04093_ _04094_ _03574_ _08757_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16716_ _06560_ _06951_ _06816_ _07125_ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__or4_4
X_17696_ _08194_ _08195_ vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16647_ _07050_ _07052_ vssd1 vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__and2_1
X_13859_ _04019_ _03847_ vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16578_ _06888_ _06896_ _06977_ vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15529_ _05831_ _05749_ _05840_ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18317_ _08802_ _08807_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _08794_ _08795_ vssd1 vssd1 vccd1 vccd1 _08796_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ _08620_ _08622_ _08719_ vssd1 vssd1 vccd1 vccd1 _08721_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09952_ _08951_ _08962_ _08930_ _08941_ vssd1 vssd1 vccd1 vccd1 _08984_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _07853_ _08224_ _07810_ vssd1 vssd1 vccd1 vccd1 _08235_ sky130_fd_sc_hd__a21oi_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11210_ _01299_ _01302_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__xnor2_1
X_12190_ _02129_ _02130_ _02131_ _02123_ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_102_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11141_ _01231_ _01232_ _01218_ _01228_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11072_ _01156_ _01163_ _01164_ vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a21bo_1
Xoutput77 net77 vssd1 vssd1 vccd1 vccd1 leds[5] sky130_fd_sc_hd__buf_2
XFILLER_0_37_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput88 net88 vssd1 vssd1 vccd1 vccd1 o_wb_data[14] sky130_fd_sc_hd__clkbuf_4
Xoutput99 net99 vssd1 vssd1 vccd1 vccd1 o_wb_data[24] sky130_fd_sc_hd__clkbuf_4
X_14900_ _05155_ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__xnor2_1
X_10023_ _00115_ _00108_ _00111_ _00113_ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__a22oi_1
X_15880_ _06128_ _06180_ vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__nor2_1
X_14831_ _03033_ _03091_ _03062_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__mux2_1
X_17550_ _03119_ _05423_ _06505_ _08036_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__o22a_1
X_14762_ _07635_ _01866_ _05005_ _05002_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11974_ _02056_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__or2b_1
X_16501_ _06749_ _06762_ vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__nand2_1
X_13713_ _03701_ _03709_ _03860_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__a21bo_1
X_10925_ _01016_ _01017_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__nand2_1
X_17481_ _07959_ _07960_ vssd1 vssd1 vccd1 vccd1 _07961_ sky130_fd_sc_hd__xnor2_1
X_14693_ _04758_ _04803_ _04931_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16432_ _06801_ _06818_ vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__xnor2_1
X_13644_ _03772_ _03773_ _03783_ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__or3_4
X_10856_ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00949_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _03077_ _06741_ _06744_ _06487_ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__o2bb2a_1
X_13575_ _03701_ _03709_ vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__xnor2_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _00877_ _00878_ _00879_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _07195_ _07741_ vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__nor2_1
X_15314_ _03368_ _03072_ _05494_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__nand3_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12526_ net137 _02614_ _02604_ _02613_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_124_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16294_ _06659_ _06668_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18033_ _08548_ _08562_ vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__xor2_1
X_15245_ _05324_ _05439_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__nand2_1
X_12457_ _02545_ _02548_ _02549_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__nand3_1
XFILLER_0_112_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11408_ _01447_ _01450_ _01499_ _01500_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__a211o_1
X_15176_ _05430_ _05342_ _05456_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__and3_1
X_12388_ _02409_ _02480_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14127_ _04299_ _04300_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__or3_4
XFILLER_0_50_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11339_ _01430_ _01431_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18935_ clknet_4_2_0_clk _00089_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[21\] sky130_fd_sc_hd__dfxtp_2
X_14058_ _02968_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__clkbuf_8
X_13009_ _00593_ _03101_ _02505_ vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__mux2_1
X_18866_ clknet_4_5_0_clk net309 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__dfxtp_1
X_17817_ _08252_ _08223_ _08326_ vssd1 vssd1 vccd1 vccd1 _08328_ sky130_fd_sc_hd__nand3_1
X_18797_ _02998_ net49 _09301_ vssd1 vssd1 vccd1 vccd1 _09307_ sky130_fd_sc_hd__mux2_1
X_17748_ _08216_ _08217_ vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17679_ _07109_ _07665_ vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_876 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09935_ _08735_ _08789_ vssd1 vssd1 vccd1 vccd1 _08800_ sky130_fd_sc_hd__xnor2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ cla_inst.in1\[19\] vssd1 vssd1 vccd1 vccd1 _08049_ sky130_fd_sc_hd__clkbuf_4
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09797_ _07265_ _07286_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__nand2_2
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _05235_ _05878_ vssd1 vssd1 vccd1 vccd1 _00803_ sky130_fd_sc_hd__nand2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11690_ _01741_ _01756_ _01781_ _01782_ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__a211o_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _00723_ _00524_ _00732_ vssd1 vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ _00184_ _00174_ _03815_ _03914_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10572_ _00513_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__buf_4
XFILLER_0_8_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12311_ _02334_ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13291_ _04515_ _04438_ _00308_ _06689_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__nand4_2
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15030_ _05188_ _05206_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ _07613_ _02205_ _02334_ vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12173_ _02235_ _02238_ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11124_ _01132_ _01205_ _01216_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__and3_1
X_16981_ _06816_ _06880_ _06944_ _07115_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__or4_1
X_18720_ net58 _03155_ _09182_ vssd1 vssd1 vccd1 vccd1 _09246_ sky130_fd_sc_hd__mux2_1
X_11055_ _01079_ _01146_ _01145_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__a21o_1
X_15932_ _06273_ _06276_ vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__or2_1
X_10006_ cla_inst.in2\[26\] vssd1 vssd1 vccd1 vccd1 _09349_ sky130_fd_sc_hd__buf_2
X_15863_ _06153_ _06157_ _06158_ vssd1 vssd1 vccd1 vccd1 _06204_ sky130_fd_sc_hd__or3_1
X_18651_ net61 _03166_ _09193_ vssd1 vssd1 vccd1 vccd1 _09196_ sky130_fd_sc_hd__mux2_1
X_14814_ _05014_ _05015_ _05062_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__a21o_1
X_17602_ _07630_ _07516_ _07982_ _07980_ vssd1 vssd1 vccd1 vccd1 _08094_ sky130_fd_sc_hd__o31a_1
X_15794_ _06128_ _06129_ vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__nand2_1
X_18582_ _09127_ vssd1 vssd1 vccd1 vccd1 _09146_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14745_ _02200_ _03153_ _04846_ vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17533_ _08016_ _08018_ _06649_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__o21ai_1
X_11957_ _02043_ _02047_ _02048_ _02049_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__or4_4
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ _05399_ _05355_ _04449_ _04471_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__and4_1
X_17464_ _06764_ _07593_ vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__nor2_1
X_14676_ _04911_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11888_ _01971_ _01973_ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16415_ _06578_ _06764_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__or2_1
X_13627_ _03990_ _00308_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__nand2_1
X_10839_ _00916_ _00914_ _00915_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__nand3_1
X_17395_ _07207_ _07751_ net146 _06947_ vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16346_ _03049_ _06609_ _06725_ _06467_ vssd1 vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13558_ _03690_ _03482_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ _02553_ _02600_ _02599_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__nand3_1
X_16277_ _00218_ _06568_ _06650_ _03313_ vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__o22a_4
XFILLER_0_113_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13489_ _03610_ _03613_ _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15228_ _05512_ _05514_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__xnor2_1
X_18016_ _08541_ _08542_ _08543_ vssd1 vssd1 vccd1 vccd1 _08544_ sky130_fd_sc_hd__or3_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15159_ _05437_ _05438_ vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09720_ _05017_ vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__buf_6
X_18918_ clknet_4_11_0_clk _00072_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_09651_ _05704_ vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__clkbuf_8
X_18849_ clknet_4_6_0_clk net294 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__dfxtp_1
X_09582_ _03946_ _03957_ _03706_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold140 net104 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 net106 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09918_ _06460_ vssd1 vssd1 vccd1 vccd1 _08615_ sky130_fd_sc_hd__buf_6
X_09849_ _07853_ _07744_ _07766_ vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__a21o_1
X_12860_ _00900_ _00903_ _00902_ vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__o21a_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _01897_ _01898_ _01876_ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__a21oi_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _01450_ _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__nand2_2
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _04603_ _04752_ vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__xnor2_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _01833_ _01834_ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__xnor2_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14461_ _04566_ _04538_ _04676_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__o211a_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11673_ _01764_ _01765_ vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__or2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _06564_ _06566_ _03313_ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ _03355_ _03362_ _03529_ _03530_ _02969_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__a311o_1
X_10624_ _00163_ _00716_ vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__nand2_1
X_17180_ _07042_ _07303_ _07130_ _07302_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__o22a_1
X_14392_ _04600_ _04601_ _04304_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16131_ _06467_ _06491_ vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__nand2_1
X_13343_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__buf_4
X_10555_ _05453_ _00645_ _06732_ _05715_ vssd1 vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__nand4_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16062_ op_code\[3\] op_code\[2\] vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__nand2b_2
X_13274_ _01521_ _05050_ net240 _03378_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__nand4_1
X_10486_ _00577_ _00576_ _00373_ _00370_ vssd1 vssd1 vccd1 vccd1 _00579_ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15013_ _05278_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__xor2_2
X_12225_ _02315_ _02316_ _02302_ _02314_ vssd1 vssd1 vccd1 vccd1 _02318_ sky130_fd_sc_hd__a211oi_2
X_12156_ _02233_ _02232_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__and2b_1
X_11107_ _01179_ _01180_ _01166_ _01178_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__a211o_1
X_12087_ _05301_ _00130_ _09212_ _05279_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a22o_1
X_16964_ _07393_ _07397_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__nand2_1
X_18703_ net51 _09190_ _09233_ vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__o21a_1
X_11038_ _01096_ _01125_ _01124_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__a21o_1
X_15915_ _06258_ _06259_ vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__nand2_1
X_16895_ _07310_ _07321_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__nand2_1
X_18634_ _09181_ vssd1 vssd1 vccd1 vccd1 _09182_ sky130_fd_sc_hd__clkbuf_4
X_15846_ _06076_ _06079_ _06185_ vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__a21o_1
X_18565_ net250 _09098_ _09133_ _09126_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__o211a_1
X_15777_ _06032_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and2_1
X_12989_ _03063_ _03078_ _03081_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__mux2_2
XFILLER_0_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17516_ _07856_ _07857_ _07874_ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14728_ _04730_ _04833_ _04862_ _04863_ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__a211oi_4
X_18496_ _03011_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _09064_ sky130_fd_sc_hd__a21o_1
X_14659_ _00877_ _01112_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__nand2_1
X_17447_ _06376_ _06375_ _06372_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17378_ _07841_ _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16329_ _01677_ _02370_ _03175_ vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09703_ _04984_ _04700_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__nand2_4
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09634_ _05235_ _05486_ _05475_ _05519_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nand4_2
X_09565_ _03356_ _03377_ _03914_ _03476_ vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nand4_1
XFILLER_0_78_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09496_ _04001_ _04012_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__nand2_8
XFILLER_0_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10340_ _03465_ _04395_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _00361_ _00363_ vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12010_ _02098_ _02101_ _02102_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__a21boi_1
X_13961_ _05453_ _09248_ _04130_ vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__a21boi_1
X_12912_ cla_inst.in2\[31\] vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__clkbuf_4
X_15700_ _06025_ _06026_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nor2_1
X_16680_ _07086_ _07088_ _04247_ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__mux2_2
X_13892_ _04052_ _04053_ _04054_ vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__o21ai_1
X_12843_ _02933_ _02934_ _02935_ _02913_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o211a_1
X_15631_ _05947_ _05951_ _05952_ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__a21oi_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15562_ _05875_ _05877_ _03202_ vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__o21ai_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _08903_ _08905_ vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__or2_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _01806_ vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__inv_2
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14513_ _04723_ _04724_ _04734_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _07738_ _07764_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__xnor2_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _00146_ _01537_ _01536_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18281_ _03056_ _06463_ _08831_ vssd1 vssd1 vccd1 vccd1 _09403_ sky130_fd_sc_hd__a21oi_2
X_15493_ _05087_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14444_ _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17232_ _04725_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11656_ _01744_ _01747_ _01698_ vssd1 vssd1 vccd1 vccd1 _01749_ sky130_fd_sc_hd__o21ai_1
X_10607_ _00568_ _00569_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__nand2_1
X_17163_ _07606_ _07614_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _04581_ _04582_ _04583_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__and3_4
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _01673_ _01675_ vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__and2_1
X_16114_ _06469_ _06473_ _03099_ vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__mux2_1
X_13326_ _03286_ _03287_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10538_ _00622_ _00630_ vssd1 vssd1 vccd1 vccd1 _00631_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17094_ _07411_ _07414_ _07412_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__o21a_1
X_16045_ _02994_ _04900_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__or2_1
X_13257_ _03358_ _03361_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__nand2_1
X_10469_ _00203_ _00399_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12208_ _02134_ _02149_ _02150_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _03286_ _03287_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__xor2_2
XFILLER_0_19_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12139_ _07243_ _00949_ _03421_ _07221_ vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a22o_1
X_17996_ _03000_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__a21oi_1
X_16947_ _07339_ _07340_ vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16878_ _06816_ _07302_ _07303_ _06764_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__o22a_1
X_18617_ net263 _09157_ _09169_ _09162_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__o211a_1
X_15829_ _06104_ _06108_ _06166_ vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__a21o_1
X_18548_ net28 _09109_ vssd1 vssd1 vccd1 vccd1 _09119_ sky130_fd_sc_hd__or2_1
X_18479_ _09036_ _09008_ _09043_ vssd1 vssd1 vccd1 vccd1 _09045_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09617_ _05279_ _05301_ _05322_ _05333_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09548_ _04580_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09479_ _03826_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11510_ _01562_ _01563_ _01525_ _01540_ vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ _02580_ _02582_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__nor2_1
X_11441_ _01529_ _01532_ _01530_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire136 _03205_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__buf_1
XFILLER_0_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _04347_ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__nand2_1
X_11372_ _01382_ _01392_ _00821_ _01463_ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a211o_2
XFILLER_0_150_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _00620_ _00621_ _00631_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__nor3_1
X_10323_ _00396_ _00397_ _00415_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a21oi_1
X_14091_ net173 _04095_ _04271_ _04272_ vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13042_ _03028_ _01692_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nor2_1
X_10254_ _00341_ _00346_ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17850_ _08349_ _08350_ _08362_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__a21o_1
X_10185_ _00275_ _00276_ _00277_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__nand3_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16801_ _07217_ _07219_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__nand2_1
X_17781_ _08279_ _08286_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__nor2_1
X_14993_ _05256_ _05258_ vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__xnor2_1
X_16732_ _07142_ _07144_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__or2_1
X_13944_ _04111_ _04112_ _04548_ _07722_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_89_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13875_ _04029_ _04037_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__xnor2_2
X_16663_ _07068_ _07070_ vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__xor2_1
X_18402_ _08907_ _08946_ _08960_ vssd1 vssd1 vccd1 vccd1 _08963_ sky130_fd_sc_hd__and3_1
X_15614_ _05846_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__inv_2
X_12826_ _02916_ _02917_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__nand2_1
X_16594_ _06343_ _06345_ _06995_ vssd1 vssd1 vccd1 vccd1 _06996_ sky130_fd_sc_hd__a21o_1
X_18333_ _08888_ _06403_ _06402_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__a21oi_1
X_15545_ _05858_ _05846_ _05847_ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__and3_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _02330_ _02849_ vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__nor2_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11708_ _01790_ _01799_ _01798_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15476_ _05665_ _05668_ _05783_ vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__or3_1
X_18264_ _03055_ _06511_ _01359_ vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__and3b_1
X_12688_ _06993_ _07646_ _02779_ _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_154_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14427_ _04630_ _04640_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__nor2_1
X_17215_ _07671_ _07558_ vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _01730_ _01726_ _01725_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__and3b_1
XFILLER_0_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18195_ _08696_ _08738_ vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14358_ _04425_ _04382_ _04540_ _04541_ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17146_ _07595_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13309_ _05410_ _05301_ _07004_ _07102_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__nand4_2
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17077_ _07519_ _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__nand2_1
X_14289_ _04487_ _04488_ _04315_ _04331_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16028_ _06377_ _06378_ _06379_ vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17979_ _08502_ _08503_ vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold88 _00008_ vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _02003_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__xor2_1
Xhold99 _00010_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _03531_ _03509_ _00130_ _07548_ vssd1 vssd1 vccd1 vccd1 _01034_ sky130_fd_sc_hd__nand4_2
X_13660_ _03794_ _03800_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ _00963_ _00964_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12611_ _02701_ _02702_ _02703_ vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__nand3_1
XFILLER_0_38_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13591_ _03724_ _03725_ _03726_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15330_ _05624_ vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__inv_2
X_12542_ _02602_ _02598_ _02601_ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__nand3_1
XFILLER_0_94_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15261_ _05526_ _05527_ _05548_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__or3_1
X_12473_ _02544_ _02557_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_136_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14212_ _04233_ _04235_ _04065_ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__o21bai_1
X_17000_ _07435_ _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__xnor2_1
X_11424_ _04984_ _00181_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15192_ _05350_ _05358_ _05474_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_8 _00461_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14143_ _04315_ _04316_ _04328_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__nor3_2
X_11355_ _01352_ _01354_ _01351_ vssd1 vssd1 vccd1 vccd1 _01448_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_104_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _00398_ vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__clkbuf_8
X_18951_ clknet_4_1_0_clk _09412_ vssd1 vssd1 vccd1 vccd1 salida\[4\] sky130_fd_sc_hd__dfxtp_1
X_14074_ _03080_ _02981_ _03560_ vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__or3_1
X_11286_ _01290_ _01308_ _01309_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__nor3_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17902_ _06559_ _08419_ vssd1 vssd1 vccd1 vccd1 _08421_ sky130_fd_sc_hd__or2_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _03082_ _03116_ _03117_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__mux2_1
X_10237_ _00326_ _00327_ _00329_ vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__a21o_1
X_18882_ clknet_4_9_0_clk _00036_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17833_ _06649_ _08327_ _08328_ _08345_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__a31o_1
X_10168_ _00252_ _00260_ vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__xnor2_1
X_17764_ _08268_ _08269_ vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__nand2_1
X_14976_ _05228_ _05239_ vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__xnor2_2
X_10099_ _00191_ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16715_ _07124_ _06816_ _07126_ net237 vssd1 vssd1 vccd1 vccd1 _07127_ sky130_fd_sc_hd__o22a_1
X_13927_ _03345_ net172 cla_inst.in1\[22\] cla_inst.in1\[20\] vssd1 vssd1 vccd1 vccd1
+ _04094_ sky130_fd_sc_hd__and4_1
X_17695_ _08090_ _08091_ _08088_ vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16646_ _06952_ _06958_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__o21ai_1
X_13858_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12809_ _01458_ _01460_ _02900_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__nor3_1
X_16577_ _06867_ _06887_ vssd1 vssd1 vccd1 vccd1 _06977_ sky130_fd_sc_hd__or2b_1
X_13789_ _03728_ _07962_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18316_ _08868_ _08869_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15528_ _05831_ _05749_ _05840_ vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18247_ _08712_ _08726_ _08793_ vssd1 vssd1 vccd1 vccd1 _08795_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15459_ _05763_ _05765_ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ _08620_ _08622_ _08719_ vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17129_ _07577_ _06845_ _02979_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09951_ _08930_ _08941_ _08951_ _08962_ vssd1 vssd1 vccd1 vccd1 _08973_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _08169_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__buf_6
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ _01218_ _01228_ _01231_ _01232_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11071_ _01157_ _01158_ _01162_ vssd1 vssd1 vccd1 vccd1 _01164_ sky130_fd_sc_hd__nand3_1
XFILLER_0_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput78 net78 vssd1 vssd1 vccd1 vccd1 leds[6] sky130_fd_sc_hd__buf_2
Xoutput89 net89 vssd1 vssd1 vccd1 vccd1 o_wb_data[15] sky130_fd_sc_hd__clkbuf_4
X_10022_ _00107_ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__buf_4
X_14830_ _05077_ _05079_ _03202_ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14761_ _05003_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__inv_2
X_11973_ _02061_ _02062_ _02065_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a21bo_1
X_16500_ _06527_ _06809_ _06891_ _06892_ vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__a31o_1
X_13712_ _03702_ _03708_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nand2_1
X_10924_ _01014_ _01015_ _00989_ _00997_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__a211o_1
X_14692_ _04928_ _04929_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__or2_1
X_17480_ _07106_ _07332_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16431_ _06809_ _06817_ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13643_ net329 _03773_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__o21ai_2
X_10855_ _00942_ _00947_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ _03702_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__xor2_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _03164_ _06742_ vssd1 vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__nand2_1
X_10786_ _00870_ _00875_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__xnor2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _07390_ _07650_ _08535_ _08534_ vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__a31o_1
X_15313_ _05491_ _05493_ vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__or2b_1
X_12525_ _02616_ _02617_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _06659_ _06668_ vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18032_ _08559_ _08560_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__and2_1
X_15244_ _05528_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__xnor2_1
X_12456_ _00832_ _00171_ _02494_ _02493_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11407_ _01430_ _01498_ _01496_ _01497_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__a211oi_2
X_15175_ _05430_ _05342_ _05456_ vssd1 vssd1 vccd1 vccd1 _05457_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12387_ _02360_ _02408_ _02406_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14126_ _04301_ _04311_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__xnor2_1
X_11338_ _01429_ _01347_ _01423_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__or3_1
X_18934_ clknet_4_8_0_clk _00088_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[20\] sky130_fd_sc_hd__dfxtp_2
X_14057_ _04065_ _04072_ _04236_ vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__a21oi_1
X_11269_ _01355_ _01361_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__nor2_1
X_13008_ _00248_ vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__clkbuf_4
X_18865_ clknet_4_4_0_clk net268 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__dfxtp_1
X_17816_ _08252_ _08223_ _08326_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__a21o_1
X_18796_ _09306_ vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__clkbuf_1
X_17747_ _08249_ _02329_ _08227_ _08250_ _02969_ vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__a311oi_2
X_14959_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17678_ _08174_ _08175_ vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__nand2_1
X_16629_ _00398_ _07032_ vssd1 vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09934_ _08768_ _08778_ vssd1 vssd1 vccd1 vccd1 _08789_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09865_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _08039_ sky130_fd_sc_hd__clkbuf_4
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _06982_ _07156_ _07265_ _07276_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__nand4_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ _00723_ _00524_ _00732_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _00496_ _00505_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12310_ _05235_ _09219_ _02332_ _02333_ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13290_ _04438_ _05704_ _06689_ _04646_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ _08713_ _00127_ _02332_ _02333_ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ _02111_ _02119_ vssd1 vssd1 vccd1 vccd1 _02265_ sky130_fd_sc_hd__xnor2_1
X_11123_ _01209_ _01214_ _01215_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16980_ _07413_ _07414_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__xnor2_1
X_11054_ _01079_ _01145_ _01146_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__nand3_2
X_15931_ _06274_ _06250_ _06275_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or3b_1
X_10005_ _06938_ _08311_ _09344_ _09347_ vssd1 vssd1 vccd1 vccd1 _09348_ sky130_fd_sc_hd__a211o_4
X_18650_ _09195_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15862_ _06199_ _06201_ vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nor2_1
X_17601_ _08090_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__xor2_1
X_14813_ _05014_ _05015_ _05062_ vssd1 vssd1 vccd1 vccd1 _05063_ sky130_fd_sc_hd__nand3_2
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18581_ net306 _09140_ _09143_ _09144_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__o211a_1
X_15793_ _06058_ _06087_ _06126_ vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nand3_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17532_ _07900_ _07903_ _07901_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__o21ai_4
X_14744_ _04982_ _04983_ _04985_ vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11956_ _01964_ _02046_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907_ _08713_ _04580_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__nand2_1
X_17463_ _07938_ _07941_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__xnor2_1
X_14675_ _00106_ _05486_ _04909_ _04910_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__o2bb2a_1
X_11887_ _01979_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16414_ _06572_ _06756_ vssd1 vssd1 vccd1 vccd1 _06800_ sky130_fd_sc_hd__nor2_1
X_13626_ _06689_ _03763_ _03764_ vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__a21bo_1
X_10838_ _00929_ _00930_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17394_ _07302_ _07303_ _07126_ _07318_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__or4_1
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16345_ _02982_ _06614_ vssd1 vssd1 vccd1 vccd1 _06725_ sky130_fd_sc_hd__or2_1
X_10769_ _07853_ _00318_ _00861_ vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__and3_2
X_13557_ _03478_ _03479_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12508_ _02553_ _02599_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__a21o_1
X_13488_ _04690_ _07112_ _03611_ _03612_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__a22o_1
X_16276_ _03410_ _06528_ _06565_ _06539_ _06520_ vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__o32a_1
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18015_ _08459_ _08460_ _08540_ vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__and3_1
X_15227_ _05513_ _05381_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__nand2_1
X_12439_ _02479_ _02481_ vssd1 vssd1 vccd1 vccd1 _02532_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15158_ _05316_ _05433_ _05436_ vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__o21ai_2
X_14109_ _04291_ _04292_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__nand2_1
X_15089_ _05360_ _05362_ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18917_ clknet_4_13_0_clk _00071_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09650_ _05693_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__buf_6
X_18848_ clknet_4_6_0_clk net307 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__dfxtp_1
X_09581_ _04842_ _04930_ _04919_ vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__a21o_1
X_18779_ _09292_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold130 net85 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _00033_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 salida\[2\] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_1
XFILLER_0_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09917_ _08539_ _08594_ vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__xnor2_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _07788_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__clkbuf_8
X_09779_ cla_inst.in1\[25\] vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__buf_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _01747_ _01901_ _01902_ vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__a21bo_2
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _01446_ _01449_ _01448_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__o21ai_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11741_ _01591_ _01590_ vssd1 vssd1 vccd1 vccd1 _01834_ sky130_fd_sc_hd__and2b_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _04628_ _04629_ _04674_ _04675_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a2bb2o_1
X_11672_ _01763_ _01762_ _01716_ _01713_ vssd1 vssd1 vccd1 vccd1 _01765_ sky130_fd_sc_hd__o211a_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13411_ _03355_ _03362_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__a21oi_1
X_10623_ _00715_ vssd1 vssd1 vccd1 vccd1 _00716_ sky130_fd_sc_hd__buf_6
XFILLER_0_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14391_ _04447_ _04455_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13342_ _00509_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16130_ _06489_ _06490_ _01677_ vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ _05464_ _07962_ _05715_ _05453_ vssd1 vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _03574_ _05050_ net241 _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__a22o_1
X_16061_ _06200_ _06246_ vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__or2_1
X_10485_ _00370_ _00373_ _00576_ _00577_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15012_ _01873_ _03067_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__nand2_1
X_12224_ _02302_ _02314_ _02315_ _02316_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _07352_ _04056_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__nand2_1
X_11106_ _01196_ _01197_ _01187_ _01192_ vssd1 vssd1 vccd1 vccd1 _01199_ sky130_fd_sc_hd__o211ai_2
X_12086_ _02178_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__inv_2
X_16963_ _06655_ _07394_ _07396_ _07113_ vssd1 vssd1 vccd1 vccd1 _07397_ sky130_fd_sc_hd__a22o_1
X_18702_ _06776_ _09183_ net69 vssd1 vssd1 vccd1 vccd1 _09233_ sky130_fd_sc_hd__a21oi_1
X_11037_ _01127_ _01129_ vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__nand2_1
X_15914_ _06257_ _06236_ vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__or2b_1
X_16894_ _07310_ _07321_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__or2_1
X_18633_ _09119_ _09180_ vssd1 vssd1 vccd1 vccd1 _09181_ sky130_fd_sc_hd__or2_1
X_15845_ _06074_ _06137_ vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18564_ salida\[4\] _09114_ _09118_ salida\[36\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09133_ sky130_fd_sc_hd__a221o_1
X_15776_ _06108_ _06109_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__nand2_1
X_12988_ _03080_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__buf_4
X_17515_ _07997_ _07998_ vssd1 vssd1 vccd1 vccd1 _07999_ sky130_fd_sc_hd__nor2_1
X_14727_ _04867_ _04868_ _04879_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11939_ _06008_ _05584_ _03421_ _04220_ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and4_1
X_18495_ _03155_ _06451_ vssd1 vssd1 vccd1 vccd1 _09063_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ _02974_ _03119_ _05306_ _07923_ vssd1 vssd1 vccd1 vccd1 _07924_ sky130_fd_sc_hd__o31a_1
X_14658_ _04891_ _04892_ vssd1 vssd1 vccd1 vccd1 _04893_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _03741_ _03746_ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or2_1
X_17377_ _07843_ _07847_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14589_ _04816_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16328_ _03089_ _06495_ _06706_ _06626_ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_858 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16259_ _06470_ _06631_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09702_ _06234_ _06245_ _06256_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__nand3_1
X_09633_ _05464_ _05388_ _05497_ _05508_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _04318_ _04744_ _04755_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__nand3_2
XFILLER_0_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09495_ _03815_ vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__buf_8
XFILLER_0_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10270_ _00362_ _00134_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13960_ _00645_ _09256_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__nand2_1
X_12911_ _04493_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__or3_4
X_13891_ _04052_ _04053_ _04054_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15630_ _05947_ _05951_ _03202_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__o21ai_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _02895_ _02915_ vssd1 vssd1 vccd1 vccd1 _02935_ sky130_fd_sc_hd__nand2_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _05789_ _05796_ _05876_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__a21oi_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _02853_ _02865_ vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__xnor2_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _07762_ _07763_ vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__nor2_1
X_14512_ _04726_ _04732_ vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__xnor2_2
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _04690_ _00218_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__nand2_1
X_18280_ _03206_ _08812_ _08818_ _08830_ vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__o211a_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _04823_ _05797_ _05798_ _05801_ vssd1 vssd1 vccd1 vccd1 _09365_ sky130_fd_sc_hd__a31o_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17231_ _03913_ _06913_ _03920_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14443_ _00107_ _06482_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nand2_1
X_11655_ _01698_ _01744_ _01747_ vssd1 vssd1 vccd1 vccd1 _01748_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10606_ _00349_ _00531_ _00529_ _00530_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__a211oi_2
X_17162_ _07488_ _07612_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__xnor2_1
X_14374_ _04435_ _04441_ _04434_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__a21bo_1
X_11586_ _01677_ _01678_ _01672_ vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16113_ _02983_ _02563_ _03173_ _06470_ _06472_ vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__o311a_1
X_13325_ _03278_ _03288_ vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__nand2_1
X_10537_ _00628_ _00629_ vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__and2b_1
X_17093_ _07409_ _07424_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16044_ _06396_ _06397_ _05162_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__a21o_1
X_10468_ _00204_ _00248_ _00410_ vssd1 vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__and3_1
X_13256_ _02963_ _03359_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _02148_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__inv_2
X_13187_ _00666_ _00674_ _00672_ vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__a21oi_2
X_10399_ _00341_ _00346_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _02203_ _02228_ _02229_ vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__nor3_1
X_17995_ _06426_ _06445_ _08521_ vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__or3_1
X_12069_ _02079_ _02078_ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__nor2_1
X_16946_ _03101_ _06464_ _07351_ _07378_ vssd1 vssd1 vccd1 vccd1 _09387_ sky130_fd_sc_hd__o2bb2a_1
X_16877_ _07115_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__clkbuf_4
X_18616_ salida\[25\] _09159_ _09160_ salida\[57\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09169_ sky130_fd_sc_hd__a221o_1
X_15828_ _06095_ _06165_ vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__xnor2_1
X_18547_ _09117_ vssd1 vssd1 vccd1 vccd1 _09118_ sky130_fd_sc_hd__buf_2
X_15759_ _06089_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18478_ _09036_ _09008_ _09043_ vssd1 vssd1 vccd1 vccd1 _09044_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ _07902_ _07903_ _07904_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09616_ net234 vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__buf_6
XFILLER_0_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09547_ _04569_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__buf_6
X_09478_ ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03826_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11440_ _01529_ _01530_ _01532_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_135_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire148 net149 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ _00821_ _01463_ _01382_ _01392_ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13110_ _00696_ _00697_ _00743_ _00744_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__nor4_2
X_10322_ _00400_ _00414_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ _01521_ _05964_ _04269_ _04270_ vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _02976_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__nor2_1
X_10253_ _00342_ _00345_ vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10184_ _03377_ _04471_ _03903_ _03356_ vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16800_ net334 _06951_ _06961_ _07218_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__or4_4
X_17780_ _08279_ _08286_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__and2_1
X_14992_ _05143_ _05153_ _05151_ vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16731_ _06665_ _07143_ vssd1 vssd1 vccd1 vccd1 _07144_ sky130_fd_sc_hd__or2_1
X_13943_ _04635_ _04427_ cla_inst.in1\[27\] _07004_ vssd1 vssd1 vccd1 vccd1 _04112_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16662_ _06983_ _06985_ _06981_ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__a21o_1
X_13874_ _04030_ _04036_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__xnor2_2
X_18401_ _08907_ _08946_ _08960_ vssd1 vssd1 vccd1 vccd1 _08961_ sky130_fd_sc_hd__a21oi_1
X_15613_ _05931_ _05933_ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__or2_1
X_12825_ _02916_ _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__or2_1
X_16593_ _06346_ _06926_ _02358_ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a21o_1
X_18332_ _01417_ _03143_ vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15544_ _05846_ _05847_ _05858_ vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__a21oi_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12756_ _02847_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _01790_ _01798_ _01799_ vssd1 vssd1 vccd1 vccd1 _01800_ sky130_fd_sc_hd__or3_4
X_18263_ _01359_ _06512_ _03056_ vssd1 vssd1 vccd1 vccd1 _08813_ sky130_fd_sc_hd__a21boi_1
X_15475_ _05665_ _05668_ _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__o21ai_1
X_12687_ _07091_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_127_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17214_ _07554_ _07555_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__and2b_1
X_14426_ _04638_ _04639_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__or2_1
X_11638_ _01725_ _01726_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__a21boi_1
X_18194_ _08736_ _08737_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17145_ _04725_ _06889_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__and2_1
X_14357_ _04540_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11569_ _03399_ _01659_ _01661_ vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ _05301_ _07004_ _07102_ _05279_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17076_ _06944_ _06957_ _07207_ _06969_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__a2bb2o_1
X_14288_ _04315_ _04331_ _04487_ _04488_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16027_ _02989_ _03693_ vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__nand2_1
X_13239_ _03295_ _03296_ _03339_ _03340_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a22o_2
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17978_ _08403_ _08448_ _08501_ vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__or3_1
XFILLER_0_34_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16929_ _07168_ _07170_ _07259_ _07359_ vssd1 vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold89 net110 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ net242 _00196_ _09179_ _03345_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10871_ _00910_ _00912_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _02662_ _02695_ _02700_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__o21bai_1
X_13590_ _03512_ _03514_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12541_ _02616_ _02629_ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15260_ _05526_ _05527_ _05548_ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__o21ai_1
X_12472_ _02558_ _02560_ _02562_ _02564_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__nor4_1
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14211_ _03745_ _04402_ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__nand2_1
X_11423_ _00197_ _01509_ _01515_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__a21bo_1
X_15191_ _05351_ _05357_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_9 _00516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14142_ _04315_ _04316_ _04328_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__o21a_1
X_11354_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10305_ _04143_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__buf_4
X_11285_ _01312_ _01332_ _01333_ _01334_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__nand4_2
X_14073_ _03561_ _03575_ _03060_ vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__mux2_1
X_18950_ clknet_4_5_0_clk _09411_ vssd1 vssd1 vccd1 vccd1 salida\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17901_ _08413_ _08418_ vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__nor2_1
X_10236_ _08800_ _08811_ _00328_ vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__a21o_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13024_ _02975_ vssd1 vssd1 vccd1 vccd1 _03117_ sky130_fd_sc_hd__buf_4
X_18881_ clknet_4_15_0_clk net318 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dfxtp_1
X_17832_ _06508_ _08332_ _08334_ _08343_ vssd1 vssd1 vccd1 vccd1 _08345_ sky130_fd_sc_hd__a31o_1
X_10167_ _00258_ _00259_ vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17763_ _06957_ _07035_ _07487_ _07593_ vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__or4_2
X_14975_ _05237_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__and2_1
X_10098_ _00175_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16714_ _07125_ vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__buf_2
X_13926_ _03509_ _05606_ _05246_ _03531_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__a22oi_2
X_17694_ _08192_ _08193_ vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16645_ _06959_ _06962_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__nand2_1
X_13857_ _04016_ _04017_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12808_ _01458_ _01460_ _02900_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__o21a_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16576_ _06967_ _06975_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__xor2_1
X_13788_ _00308_ _03940_ _03941_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_146_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18315_ _08795_ _08842_ _08867_ vssd1 vssd1 vccd1 vccd1 _08869_ sky130_fd_sc_hd__and3_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15527_ _05838_ _05839_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ _02776_ _02778_ _02798_ _02800_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18246_ _08712_ _08726_ _08793_ vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__or3_1
X_15458_ _05449_ _01317_ _05764_ _05761_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_127_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14409_ _04619_ _04620_ vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__and2_1
X_18177_ _08717_ _08718_ vssd1 vssd1 vccd1 vccd1 _08719_ sky130_fd_sc_hd__nor2_1
X_15389_ _05688_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17128_ _06469_ _06498_ _02980_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09950_ _06667_ _06798_ vssd1 vssd1 vccd1 vccd1 _08962_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17059_ _07499_ _07500_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _08191_ _07820_ vssd1 vssd1 vccd1 vccd1 _08213_ sky130_fd_sc_hd__and2b_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11070_ _01157_ _01158_ _01162_ vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput79 net79 vssd1 vssd1 vccd1 vccd1 leds[7] sky130_fd_sc_hd__buf_2
X_10021_ _00107_ _00108_ _00111_ _00113_ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__and4_1
X_14760_ _05002_ _06482_ _07635_ _05003_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__and4b_1
XFILLER_0_98_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11972_ _02023_ _02063_ _02064_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__or3_1
XFILLER_0_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13711_ _03700_ _03711_ vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__nand2_1
X_10923_ _00989_ _00997_ _01014_ _01015_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__o211ai_4
X_14691_ net202 _04883_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16430_ _06522_ _06525_ _06816_ _01113_ vssd1 vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__a211o_1
X_13642_ _03774_ _03781_ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__xnor2_2
X_10854_ _00943_ _00946_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__xnor2_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _03083_ _03166_ _03086_ _03169_ _06477_ _03161_ vssd1 vssd1 vccd1 vccd1 _06742_
+ sky130_fd_sc_hd__mux4_1
X_13573_ _03705_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10785_ _00172_ vssd1 vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__clkbuf_8
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _08553_ _08554_ _08552_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__o21ai_2
X_15312_ _05604_ _05605_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__or2_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _02561_ _02615_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _06665_ _06666_ _06582_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18031_ _08473_ _08475_ _08558_ vssd1 vssd1 vccd1 vccd1 _08560_ sky130_fd_sc_hd__or3_1
X_15243_ _05434_ _05438_ _05530_ vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ _05671_ _09212_ _02546_ _02547_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__a31o_1
X_11406_ _01496_ _01497_ _01430_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__o211a_1
X_15174_ _05443_ _05455_ vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__xnor2_1
X_12386_ _02475_ _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ _04309_ _04310_ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11337_ _01347_ _01423_ _01429_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_132_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18933_ clknet_4_12_0_clk _00087_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[19\] sky130_fd_sc_hd__dfxtp_2
X_14056_ _04233_ _04235_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__xnor2_2
X_11268_ _01358_ _01360_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ _03091_ _03097_ _03099_ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__mux2_1
X_10219_ _05464_ _06689_ _08757_ _05508_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__a22o_1
X_11199_ _01007_ _01012_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__and2_1
X_18864_ clknet_4_4_0_clk net270 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__dfxtp_1
X_17815_ _08324_ _08325_ vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18795_ _09298_ _09305_ vssd1 vssd1 vccd1 vccd1 _09306_ sky130_fd_sc_hd__and2_1
X_17746_ _08249_ _08227_ _02329_ vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__a21oi_1
X_14958_ _05109_ _05110_ _05111_ _05108_ _05106_ vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _03130_ _03172_ _03060_ vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__mux2_1
X_17677_ _07126_ _07195_ _07318_ _07608_ vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__or4_1
X_14889_ _00125_ _00459_ _05322_ _00151_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16628_ _04864_ _06812_ _06529_ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__or3_4
XFILLER_0_58_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16559_ _06954_ _06956_ _00172_ vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a21bo_4
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18229_ _00789_ _07743_ _07390_ _03311_ vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09933_ _05366_ _08757_ _05246_ _05508_ vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _07352_ _07112_ _07265_ _07276_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__a22o_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _07254_ cla_inst.in1\[24\] _05693_ _07232_ vssd1 vssd1 vccd1 vccd1 _07276_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10570_ _00497_ _00504_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12240_ _05301_ _07548_ _07591_ _05279_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12171_ _02256_ _02261_ _02262_ _02263_ vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__or4_4
X_11122_ _01129_ _01213_ _01210_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__nand3_2
XFILLER_0_102_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11053_ _01020_ _01021_ _01078_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__o21ai_1
X_15930_ _06200_ _03072_ _06249_ vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__a21o_1
X_10004_ _09341_ _09345_ _09343_ _09346_ vssd1 vssd1 vccd1 vccd1 _09347_ sky130_fd_sc_hd__a2bb2oi_2
X_15861_ _06200_ _03149_ _06198_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__a21oi_1
X_17600_ _07630_ _07511_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__or2_1
X_14812_ _05059_ _05060_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__nor2_1
X_18580_ _09125_ vssd1 vssd1 vccd1 vccd1 _09144_ sky130_fd_sc_hd__buf_2
X_15792_ _06058_ _06087_ _06126_ vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17531_ _08014_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_87_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14743_ _04982_ _04983_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nand3_4
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_160 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_160/HI led_enb[9] sky130_fd_sc_hd__conb_1
XFILLER_0_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11955_ _00845_ _01962_ _01963_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10906_ _00948_ _00952_ vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__nand2_1
X_17462_ _07829_ _07830_ _07939_ vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__a21boi_2
X_14674_ _04909_ _04910_ cla_inst.in2\[25\] _05486_ vssd1 vssd1 vccd1 vccd1 _04911_
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_86_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11886_ _01945_ _01976_ _01978_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16413_ _03083_ _06464_ _06748_ _06799_ vssd1 vssd1 vccd1 vccd1 _09411_ sky130_fd_sc_hd__o2bb2a_1
X_13625_ _03782_ cla_inst.in1\[22\] _08746_ _03848_ vssd1 vssd1 vccd1 vccd1 _03764_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10837_ _03717_ _03432_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__nand2_1
X_17393_ _07863_ _07865_ vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16344_ _03049_ _03064_ _06626_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__and3_1
X_13556_ _03687_ _03688_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__nand2_1
X_10768_ _00120_ _07123_ vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__and2_4
X_12507_ _05595_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel _07548_
+ _07581_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16275_ _06516_ vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__buf_4
X_13487_ _05017_ _07156_ _03611_ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__nand4_2
X_10699_ _00785_ _00791_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18014_ _07039_ _08150_ _08538_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15226_ _05378_ _05379_ vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__or2b_1
X_12438_ _02526_ _02530_ vssd1 vssd1 vccd1 vccd1 _02531_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15157_ _05316_ _05433_ _05436_ vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12369_ _02400_ _02461_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__nor2_1
X_14108_ _06460_ _09311_ _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__a22o_1
X_15088_ _05247_ _05254_ _05361_ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14039_ _04214_ _04215_ _04171_ _04172_ vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__o211a_1
X_18916_ clknet_4_9_0_clk _00070_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_129_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ clknet_4_1_0_clk net278 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__dfxtp_1
X_09580_ _04842_ _04919_ _04930_ vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__nand3_1
X_18778_ _09273_ _09291_ vssd1 vssd1 vccd1 vccd1 _09292_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17729_ _08023_ _08129_ _08130_ vssd1 vssd1 vccd1 vccd1 _08232_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold120 net97 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 _00015_ vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 net305 sky130_fd_sc_hd__buf_1
Xhold153 salida\[1\] vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_1
XFILLER_0_0_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09916_ _08550_ _08583_ vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _07777_ _07820_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__or2_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _07080_ vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _05224_ _03673_ vssd1 vssd1 vccd1 vccd1 _01833_ sky130_fd_sc_hd__nand2_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _01713_ _01716_ _01762_ _01763_ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a211oi_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13410_ _03527_ _03528_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__nand2_1
X_10622_ _03750_ vssd1 vssd1 vccd1 vccd1 _00715_ sky130_fd_sc_hd__buf_12
X_14390_ _04454_ _04448_ vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13341_ _05736_ _09248_ _03244_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__a31o_1
X_10553_ _00644_ _00645_ _05758_ _05975_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16060_ _06200_ _06246_ _06248_ _06414_ vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__a211o_1
X_13272_ _03531_ _03366_ net224 _04569_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__nand4_2
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10484_ _00555_ _00556_ _00575_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15011_ _05276_ _05277_ vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nor2_1
X_12223_ _02154_ _02157_ _02156_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12154_ _02244_ _02246_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__or2_1
X_11105_ _01187_ _01192_ _01196_ _01197_ vssd1 vssd1 vccd1 vccd1 _01198_ sky130_fd_sc_hd__a211o_1
X_12085_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ _00129_
+ _01031_ vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__and4_1
X_16962_ _03324_ _03003_ _06814_ _07289_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__a211oi_4
X_18701_ _09231_ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__buf_1
X_11036_ _06982_ _05845_ _01127_ _01128_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__nand4_2
X_15913_ _06236_ _06257_ vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__or2b_1
X_16893_ _07317_ _07320_ vssd1 vssd1 vccd1 vccd1 _07321_ sky130_fd_sc_hd__xnor2_1
X_15844_ _06071_ _06134_ _06136_ vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__a21o_1
X_18632_ net24 net27 _09111_ _09178_ vssd1 vssd1 vccd1 vccd1 _09180_ sky130_fd_sc_hd__or4_1
X_15775_ _06100_ _06107_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__or2_1
X_18563_ net259 _09098_ _09132_ _09126_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__o211a_1
X_12987_ _03079_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__buf_4
X_17514_ _07851_ _07878_ _07996_ vssd1 vssd1 vccd1 vccd1 _07998_ sky130_fd_sc_hd__nor3_1
X_14726_ _04882_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11938_ _06982_ _04012_ _02029_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__a31o_1
X_18494_ _02951_ _09060_ _09061_ _02968_ vssd1 vssd1 vccd1 vccd1 _09062_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17445_ _06680_ _07918_ _07922_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__nor3_1
XFILLER_0_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14657_ _04760_ _04763_ _04761_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11869_ _04700_ vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__buf_6
XFILLER_0_67_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ _02963_ _03742_ _03745_ vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ _07845_ _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14588_ net243 _04686_ _04815_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16327_ _01677_ _02125_ _03179_ vssd1 vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__or3_1
X_13539_ _03652_ _03669_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__xor2_2
XFILLER_0_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16258_ _03086_ _03169_ _00881_ _03094_ _06477_ _02983_ vssd1 vssd1 vccd1 vccd1 _06631_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15209_ _05491_ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16189_ _06508_ _06514_ _06555_ _06462_ vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09701_ _04788_ _04799_ _04777_ vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__a21bo_1
X_09632_ _05399_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09563_ _03968_ _03979_ _04307_ vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09494_ _03990_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12910_ _03771_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel vssd1
+ vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__or2_4
X_13890_ _03879_ _03882_ vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__nor2_1
X_12841_ _00884_ _02921_ _02932_ vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _05786_ _05788_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ _02863_ _02864_ vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__and2_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _04730_ _04731_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__and2_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _01813_ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _03573_ _05307_ _05800_ _03124_ vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _03081_ _07686_ _07687_ _02973_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__a211o_1
X_14442_ _04655_ _04656_ vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__nor2_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11654_ _01745_ cla_inst.in2\[20\] _01746_ _01357_ vssd1 vssd1 vccd1 vccd1 _01747_
+ sky130_fd_sc_hd__and4_4
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10605_ _00555_ _00556_ _00575_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17161_ _07607_ _07611_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14373_ _04573_ _04574_ _04579_ vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__a21o_1
X_11585_ _05888_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ _03049_ _02370_ _03175_ vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__or3_1
X_13324_ _03431_ _03433_ _03374_ _03264_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__a211oi_4
X_10536_ _00626_ _00627_ _00623_ vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__a21o_1
X_17092_ _07483_ _07430_ _07535_ vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16043_ _02997_ _01112_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13255_ _00757_ _00906_ _00758_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__o21ba_1
X_10467_ _00408_ _00409_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__and2_1
X_12206_ _02295_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__nor3_1
X_13186_ _03279_ _03285_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__xnor2_2
X_10398_ net184 net340 _00489_ _00490_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_102_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12137_ _02203_ _02228_ _02229_ vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__or3_1
X_17994_ _03044_ _06444_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__nor2_1
X_12068_ _02135_ _02159_ _02160_ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__o21ba_1
X_16945_ _07353_ _03202_ _07354_ _07377_ vssd1 vssd1 vccd1 vccd1 _07378_ sky130_fd_sc_hd__a31o_1
X_11019_ _05758_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__buf_4
X_16876_ _06944_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18615_ net287 _09157_ _09168_ _09162_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__o211a_1
X_15827_ _06163_ _06164_ vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15758_ _03010_ _03012_ _03149_ _03067_ vssd1 vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__and4_1
X_18546_ net27 _09115_ _09116_ vssd1 vssd1 vccd1 vccd1 _09117_ sky130_fd_sc_hd__nor3_2
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14709_ _04819_ _04816_ vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__nand2_1
X_15689_ _05947_ _05951_ _05945_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__o21a_1
X_18477_ _09041_ _09042_ vssd1 vssd1 vccd1 vccd1 _09043_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17428_ _07902_ _07903_ _06516_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17359_ _02977_ _07657_ net168 _06753_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__nand4_1
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09615_ _05311_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09546_ cla_inst.in1\[16\] vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09477_ _03804_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__buf_6
XFILLER_0_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire116 _08251_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire149 _09108_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11370_ _00797_ _00820_ _00819_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10321_ _00412_ _00413_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13040_ _02977_ _03131_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__or2_1
X_10252_ _00343_ _00344_ vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__and2b_1
X_10183_ _03465_ _04886_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__and2_1
X_14991_ _05132_ _05255_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__xnor2_1
X_13942_ _00294_ cla_inst.in1\[27\] _07004_ _04351_ vssd1 vssd1 vccd1 vccd1 _04111_
+ sky130_fd_sc_hd__a22oi_1
X_16730_ _07042_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__clkbuf_4
X_16661_ _07066_ _07067_ vssd1 vssd1 vccd1 vccd1 _07068_ sky130_fd_sc_hd__or2b_1
X_13873_ _04033_ _04035_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__xnor2_2
X_15612_ _05929_ _05930_ _05892_ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__a21oi_1
X_18400_ _08958_ _08959_ vssd1 vssd1 vccd1 vccd1 _08960_ sky130_fd_sc_hd__nand2_1
X_12824_ _01496_ _01500_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__nor2_2
XFILLER_0_97_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16592_ _06990_ _06991_ _06836_ vssd1 vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15543_ _05855_ _05857_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__and2_1
X_18331_ _06426_ _06448_ _08881_ _08882_ _08885_ vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__o311a_1
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _02466_ _02398_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__xnor2_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _01236_ _01789_ _01760_ _01769_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a211oi_2
X_18262_ _08773_ _08810_ vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__xnor2_2
X_15474_ _05781_ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__xor2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _07613_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14425_ _04496_ _04631_ _04637_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__o21a_1
X_17213_ _07586_ _07587_ _07667_ vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__o21a_1
X_11637_ _01727_ _01728_ _01729_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or3_1
X_18193_ _08660_ _08697_ _08734_ vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17144_ _06572_ _07487_ _07593_ _06563_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__o22a_1
X_14356_ _04560_ _04562_ _03539_ vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__mux2_1
X_11568_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel _03826_ _03388_
+ _06008_ vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13307_ _03414_ _03415_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__xor2_2
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10519_ _03881_ _03892_ _05028_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__and3_1
X_17075_ _06880_ _06944_ _06957_ _07115_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__or4_1
X_14287_ _04470_ _04472_ _04486_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11499_ _08713_ _00165_ _01590_ _01591_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16026_ _02989_ _03693_ vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__or2_1
X_13238_ _03295_ _03296_ _03339_ _03340_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__nand4_4
XFILLER_0_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13169_ _00655_ _00657_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__nand2_2
X_17977_ _08403_ _08448_ _08501_ vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__o21ai_2
X_16928_ _07165_ _07358_ _07258_ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__a21oi_1
X_16859_ _07240_ _07244_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18529_ _09097_ vssd1 vssd1 vccd1 vccd1 _09098_ sky130_fd_sc_hd__buf_2
XFILLER_0_153_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10870_ _00775_ _00962_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel vssd1 vssd1 vccd1 vccd1
+ _04384_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _02590_ _02632_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12471_ _00846_ _00214_ _02563_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_124_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14210_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__inv_2
X_11422_ _01151_ _00196_ _00871_ _03848_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15190_ _05339_ _05472_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14141_ _04317_ _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11353_ _01370_ _01374_ _01444_ _01445_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ _00395_ _00380_ _00381_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__nand3_1
X_14072_ _04240_ _04244_ _04252_ vssd1 vssd1 vccd1 vccd1 _09382_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11284_ _01337_ _01366_ _01367_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__nor3_2
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ _03100_ _03115_ _03080_ vssd1 vssd1 vccd1 vccd1 _03116_ sky130_fd_sc_hd__mux2_2
X_17900_ _08018_ _08415_ _08417_ vssd1 vssd1 vccd1 vccd1 _08418_ sky130_fd_sc_hd__o21a_1
X_10235_ _08822_ _08908_ vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__and2_1
X_18880_ clknet_4_15_0_clk net317 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__dfxtp_1
X_17831_ _06421_ _08335_ _08336_ _08342_ vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__a31o_1
X_10166_ _00216_ _00220_ vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__or2_1
X_17762_ _07130_ _07487_ _07593_ _07143_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__o22ai_1
X_14974_ _05229_ _05236_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__nand2_1
X_10097_ _00189_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__clkbuf_4
X_16713_ _06871_ _07032_ _00213_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a21bo_2
X_13925_ _03934_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__and3_1
X_17693_ _07630_ _07621_ vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__nor2_1
X_13856_ _00204_ _01866_ _04015_ vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__a21o_1
X_16644_ _06876_ _06885_ _06964_ vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _00887_ _00867_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__xor2_2
XFILLER_0_147_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13787_ _03782_ _05693_ _05606_ _03848_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16575_ _06973_ _06974_ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__or2_1
X_10999_ _01086_ _01091_ vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__xnor2_2
X_18314_ _08795_ _08842_ _08867_ vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15526_ _02998_ _03153_ _05743_ _05742_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__a31o_1
X_12738_ _02830_ _02800_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15457_ _05762_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18245_ _08791_ _08792_ vssd1 vssd1 vccd1 vccd1 _08793_ sky130_fd_sc_hd__and2_1
X_12669_ _02753_ _02761_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14408_ _04616_ _04618_ _04612_ vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15388_ _05530_ _05676_ _05687_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__nor3_1
X_18176_ _07608_ _07741_ _07859_ _07394_ vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14339_ _04542_ _04543_ _04423_ _04424_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__o211a_2
X_17127_ _06331_ _06790_ _07575_ _00558_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17058_ _07018_ _07106_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__nor2_1
X_16009_ _06356_ _06357_ _06358_ vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_148_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _07820_ _08191_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__and2b_1
XFILLER_0_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10020_ _09350_ _07570_ _07602_ _00112_ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__a22o_1
X_11971_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__xnor2_1
X_13710_ _03447_ _03710_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__or2_1
X_10922_ _00998_ _00999_ _01013_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__nand3_2
X_14690_ _04882_ _04883_ _04926_ _04927_ vssd1 vssd1 vccd1 vccd1 _04928_ sky130_fd_sc_hd__and4_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _03775_ _03780_ vssd1 vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__xor2_2
X_10853_ _00944_ _00945_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__and2b_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _06470_ _06740_ vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13572_ _09352_ _00398_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__nand2_1
X_10784_ _00203_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__buf_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15311_ _05503_ _05506_ _05603_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__and3_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _02561_ _02615_ vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _06563_ _06665_ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15242_ _05318_ _05438_ _05434_ vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__a21oi_2
X_18030_ _08473_ _08475_ _08558_ vssd1 vssd1 vccd1 vccd1 _08559_ sky130_fd_sc_hd__o21ai_2
X_12454_ _05562_ _05584_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.mux.sel vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__and4_1
XFILLER_0_124_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11405_ _01422_ _01432_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__or2b_2
XFILLER_0_90_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15173_ _05452_ _05454_ vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12385_ _02402_ _02477_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14124_ _04302_ _04117_ _04308_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11336_ _01424_ _01428_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__xnor2_2
X_14055_ _04058_ _04059_ _04234_ vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__o21ai_4
X_18932_ clknet_4_12_0_clk _00086_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[18\] sky130_fd_sc_hd__dfxtp_1
X_11267_ _01359_ _01357_ _01110_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__a21oi_1
X_13006_ _03098_ vssd1 vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__buf_4
X_10218_ _05508_ _05366_ _06689_ _08757_ vssd1 vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__and4_1
X_18863_ clknet_4_4_0_clk net264 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__dfxtp_1
X_11198_ _01004_ _01006_ vssd1 vssd1 vccd1 vccd1 _01291_ sky130_fd_sc_hd__and2_1
X_17814_ _08253_ _08254_ _08323_ vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__a21o_1
XFILLER_0_118_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10149_ _00235_ _00241_ vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__xnor2_1
X_18794_ _03000_ net48 _09301_ vssd1 vssd1 vccd1 vccd1 _09305_ sky130_fd_sc_hd__mux2_1
X_17745_ _02321_ _02325_ vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__nand2_1
X_14957_ _05210_ _05218_ vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13908_ _03930_ _04072_ _04073_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__and3_1
X_17676_ _07394_ net146 _07604_ _07751_ vssd1 vssd1 vccd1 vccd1 _08174_ sky130_fd_sc_hd__a22o_1
X_14888_ _00362_ _06482_ _05003_ _05002_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16627_ _06945_ _07030_ vssd1 vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__xnor2_1
X_13839_ _03805_ _03807_ _03996_ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16558_ sel_op\[0\] _06804_ _06955_ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15509_ _05817_ _05818_ _05813_ vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16489_ _06522_ _06525_ _06880_ _00515_ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18228_ _02045_ _00789_ _07743_ _07387_ vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__or4_1
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18159_ _06366_ _07650_ _07596_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09932_ _05410_ _05366_ _08757_ _05246_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _07951_ _08006_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__nand2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _07232_ _07254_ _06722_ _05704_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__nand4_2
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _02258_ _02260_ vssd1 vssd1 vccd1 vccd1 _02263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11121_ _01129_ _01210_ _01213_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__a21o_1
XFILLER_0_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _01120_ _01144_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__xor2_1
X_10003_ net167 _06906_ _09005_ _09016_ vssd1 vssd1 vccd1 vccd1 _09346_ sky130_fd_sc_hd__o211ai_4
X_15860_ _03007_ vssd1 vssd1 vccd1 vccd1 _06200_ sky130_fd_sc_hd__clkbuf_4
X_14811_ _05056_ _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__a21oi_1
X_15791_ _06124_ _06125_ vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nand2_1
X_17530_ _07931_ _07932_ _08013_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__or3b_4
X_14742_ _04843_ _04848_ _04841_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a21bo_1
Xwb_buttons_leds_161 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_161/HI led_enb[10] sky130_fd_sc_hd__conb_1
X_11954_ _01964_ _02046_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10905_ _00942_ _00947_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__nand2_1
X_14673_ _00109_ _09349_ _05388_ _05497_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and4_1
X_17461_ _07828_ _07827_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__or2_1
X_11885_ _01890_ _01977_ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__nand2_1
X_13624_ _04078_ _01151_ _08746_ vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__and3_1
X_16412_ _06649_ _06778_ _06779_ _06797_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__a31o_1
X_10836_ _00927_ _00928_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17392_ _06581_ _07741_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13555_ _03685_ _03686_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__nand2_1
X_16343_ _06671_ _06694_ _06719_ _06723_ _06427_ vssd1 vssd1 vccd1 vccd1 _09408_ sky130_fd_sc_hd__o32a_1
X_10767_ _00140_ _00139_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__and2b_1
XFILLER_0_81_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _00832_ _00177_ _02551_ _02552_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__a22o_1
X_16274_ _01746_ _06464_ _06648_ vssd1 vssd1 vccd1 vccd1 _09397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _04351_ _04373_ cla_inst.in1\[24\] _05693_ vssd1 vssd1 vccd1 vccd1 _03612_
+ sky130_fd_sc_hd__nand4_2
X_10698_ _00786_ _00787_ _00789_ _00790_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15225_ _05510_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__or2_1
X_18013_ _08459_ _08460_ _08540_ vssd1 vssd1 vccd1 vccd1 _08541_ sky130_fd_sc_hd__a21oi_1
X_12437_ _02523_ _02525_ _02524_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__o21a_1
XFILLER_0_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15156_ _05318_ _05434_ _05435_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12368_ _02458_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__and2b_1
X_14107_ _04290_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11319_ _01409_ _01411_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__xor2_1
X_15087_ _05253_ _05248_ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__and2b_1
X_12299_ _02385_ net123 _02390_ _02391_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__o211a_1
X_14038_ _04171_ _04172_ _04214_ _04215_ vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__a211oi_2
X_18915_ clknet_4_8_0_clk _00069_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_18846_ clknet_4_1_0_clk net272 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__dfxtp_1
X_18777_ _02989_ net42 _09276_ vssd1 vssd1 vccd1 vccd1 _09291_ sky130_fd_sc_hd__mux2_1
X_15989_ _02977_ _01248_ vssd1 vssd1 vccd1 vccd1 _06337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17728_ _01678_ _07355_ _02987_ vssd1 vssd1 vccd1 vccd1 _08231_ sky130_fd_sc_hd__or3b_1
X_17659_ _08153_ _08154_ vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 net112 vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _00026_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 net83 vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 net84 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold154 op_code\[2\] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__clkbuf_2
X_09915_ _08561_ _08572_ vssd1 vssd1 vccd1 vccd1 _08583_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09846_ _07777_ _07820_ vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__and2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _07069_ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__clkbuf_4
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ _01217_ _01219_ _01227_ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__nor3_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _00712_ _00713_ vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ _06029_ _06051_ _00498_ _08169_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and4_1
X_10552_ _05366_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__buf_6
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13271_ net172 net234 cla_inst.in1\[16\] _03345_ vssd1 vssd1 vccd1 vccd1 _03376_
+ sky130_fd_sc_hd__a22o_4
X_10483_ _00555_ _00556_ _00575_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15010_ _05263_ _05171_ _05275_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12222_ _02154_ _02156_ _02157_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12153_ _02244_ _02245_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _00217_ vssd1 vssd1 vccd1 vccd1 _02246_ sky130_fd_sc_hd__and4b_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11104_ _01193_ _01194_ _01195_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__and3_1
X_12084_ _02093_ _02096_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__xor2_1
X_16961_ _02476_ _07105_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__and2_4
X_18700_ _09209_ _09230_ vssd1 vssd1 vccd1 vccd1 _09231_ sky130_fd_sc_hd__and2_1
X_11035_ _07254_ _05333_ _05039_ _07232_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__a22o_1
X_15912_ _06254_ _06255_ vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__and2_1
X_16892_ _06579_ _07318_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__or2_1
X_18631_ net34 net67 net68 vssd1 vssd1 vccd1 vccd1 _09178_ sky130_fd_sc_hd__nand3_2
X_15843_ _06180_ _06182_ vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__xor2_2
XFILLER_0_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18562_ salida\[3\] _09114_ _09118_ salida\[35\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09132_ sky130_fd_sc_hd__a221o_1
X_15774_ _06100_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__nand2_1
X_12986_ _02780_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17513_ _07851_ _07878_ _07996_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14725_ _04794_ _04796_ _04924_ _04925_ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__o211a_1
X_11937_ _01082_ _01081_ _03826_ _03388_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__and4_1
X_18493_ _02951_ _09060_ vssd1 vssd1 vccd1 vccd1 _09061_ sky130_fd_sc_hd__nor2_1
X_17444_ _02973_ _07920_ _07921_ _06484_ vssd1 vssd1 vccd1 vccd1 _07922_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14656_ _04887_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__xnor2_2
X_11868_ _01946_ _01959_ vssd1 vssd1 vccd1 vccd1 _01961_ sky130_fd_sc_hd__xnor2_1
X_10819_ _03465_ _00909_ _00910_ _00911_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__nand4_2
X_13607_ _03358_ _03360_ _03527_ _03528_ _03744_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__a41o_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17375_ _07039_ _07108_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14587_ net244 _04686_ _04815_ vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__or3_1
X_11799_ _01887_ _01890_ _01707_ _01891_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16326_ _06698_ _06704_ _03080_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__mux2_1
X_13538_ _03667_ _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13469_ _03629_ _03596_ _05333_ _00439_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__and4_1
X_16257_ _06617_ _06629_ _04247_ vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15208_ _05375_ _05376_ _05492_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__o21ai_2
X_16188_ _06516_ _06527_ _06542_ _06554_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15139_ _05407_ _05416_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09700_ _06202_ _06224_ _06213_ vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__a21o_1
X_09631_ _05028_ vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__buf_4
X_18829_ net69 _09116_ _09180_ vssd1 vssd1 vccd1 vccd1 _09331_ sky130_fd_sc_hd__or3_4
X_09562_ _04624_ _04733_ vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__xnor2_2
X_09493_ _03717_ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09829_ _07570_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__clkbuf_4
X_12840_ _00884_ _02921_ _02932_ vssd1 vssd1 vccd1 vccd1 _02933_ sky130_fd_sc_hd__o21a_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _02860_ _02861_ _02862_ vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__o21bai_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14510_ _04576_ _04577_ _04729_ vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11722_ _01813_ _01814_ _03990_ _09212_ vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__and4b_1
XFILLER_0_84_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ _02973_ _03583_ _05799_ vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__o21ai_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14441_ _00148_ _00149_ _08452_ _04700_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__and4_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _07646_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__clkbuf_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ _00694_ _00695_ _00491_ _00535_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__o211a_1
X_14372_ _04573_ net178 _04579_ vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__nand3_1
XFILLER_0_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17160_ _07609_ _07610_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__and2b_1
X_11584_ _00845_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__buf_4
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13323_ _03374_ _03264_ _03431_ _03433_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__o211a_2
X_16111_ _06467_ vssd1 vssd1 vccd1 vccd1 _06470_ sky130_fd_sc_hd__buf_2
X_10535_ _00623_ _00626_ _00627_ vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17091_ _07483_ _07430_ _07535_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13254_ _00759_ _00908_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__and2_1
X_16042_ _06393_ _06394_ _04887_ vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__a21bo_1
X_10466_ _00163_ _00558_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ net129 _02294_ _02230_ _02282_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ _03280_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__xor2_2
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10397_ _00486_ _00487_ _00488_ _00467_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12136_ _02198_ _02199_ _02202_ vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__a21oi_1
X_17993_ _07084_ _08517_ _08519_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__or3_1
X_12067_ _02154_ _02158_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02160_ sky130_fd_sc_hd__o211a_1
X_16944_ _06508_ _07361_ _07362_ _07376_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11018_ _01107_ _01109_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__nor2_1
X_16875_ _06762_ _06890_ _06947_ _07026_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__and4_1
X_18614_ salida\[24\] _09159_ _09160_ salida\[56\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09168_ sky130_fd_sc_hd__a221o_1
X_15826_ _06037_ _05652_ _02992_ vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__and3b_1
XFILLER_0_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18545_ net28 net148 vssd1 vssd1 vccd1 vccd1 _09116_ sky130_fd_sc_hd__nand2_1
X_15757_ _03012_ _03149_ _03067_ _03010_ vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__a22oi_1
X_12969_ _03061_ vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14708_ _04551_ _04691_ _04693_ _04818_ vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__or4_4
X_18476_ _08961_ _09036_ _09004_ vssd1 vssd1 vccd1 vccd1 _09042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15688_ _06013_ _06014_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__or2_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _07790_ _07794_ _07791_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__o21a_4
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14639_ _04870_ _05921_ _03014_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__and4b_1
XFILLER_0_117_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17358_ _00557_ _07825_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16309_ _06333_ _06334_ vssd1 vssd1 vccd1 vccd1 _06686_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17289_ _07207_ _07039_ _07751_ _06947_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09614_ cla_inst.in1\[19\] vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__buf_6
XFILLER_0_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09545_ _04548_ vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03804_ sky130_fd_sc_hd__buf_6
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire117 _05408_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__buf_2
XFILLER_0_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire139 _01406_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_1
XFILLER_0_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10320_ _00411_ _00401_ _00402_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ _07080_ cla_inst.in1\[28\] _07374_ _07047_ vssd1 vssd1 vccd1 vccd1 _00344_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10182_ _03629_ _03596_ _04482_ _03815_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__nand4_2
X_14990_ _05247_ _05254_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__xor2_1
X_13941_ _04001_ _07134_ _03941_ _03940_ _00309_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16660_ _07065_ _07063_ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__or2b_1
X_13872_ cla_inst.in2\[25\] _03750_ vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__nand2_1
X_15611_ _05892_ _05929_ _05930_ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__and3_1
X_12823_ _02895_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__xnor2_1
X_16591_ _06990_ _06991_ vssd1 vssd1 vccd1 vccd1 _06992_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ _07371_ _08141_ _08884_ _06721_ vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__o211a_1
X_15542_ _05848_ _05854_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__nand2_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _02462_ _02464_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__xor2_2
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _01791_ _01797_ vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18261_ _08736_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__xnor2_2
X_15473_ _05596_ _05699_ _05697_ vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__a21oi_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _02744_ _02752_ _02775_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__a21oi_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17212_ _07586_ _07587_ _07667_ vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__nor3_1
X_14424_ _04496_ _04631_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__nor3_1
XFILLER_0_71_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11636_ _01221_ _01693_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__nor2_1
X_18192_ _08660_ _08697_ _08734_ vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17143_ _04725_ _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__nand2_4
X_11567_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel _03903_ vssd1
+ vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14355_ _03164_ _03159_ _04561_ _03916_ vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13306_ _05747_ _00513_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__nand2_1
X_10518_ _00607_ _00608_ _00609_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__a21o_1
X_14286_ _04470_ _04472_ _04486_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17074_ _07514_ _07517_ vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11498_ _00806_ _06591_ _00210_ _04220_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__and4_1
X_13237_ _03337_ _03338_ _03297_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16025_ _06372_ _06375_ _06376_ vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__a21bo_1
X_10449_ _00385_ _00392_ _00541_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _00676_ _00689_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__or2_2
X_12119_ _05638_ _00774_ _00176_ _05562_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__a22o_1
X_17976_ _08499_ _08500_ vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__xor2_1
X_13099_ _03191_ vssd1 vssd1 vccd1 vccd1 _03192_ sky130_fd_sc_hd__inv_2
X_16927_ _07257_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__inv_2
X_16858_ _02099_ _06723_ _07255_ _07282_ vssd1 vssd1 vccd1 vccd1 _09417_ sky130_fd_sc_hd__o22a_2
X_15809_ _06145_ _03906_ _03907_ _03909_ _02980_ _02978_ vssd1 vssd1 vccd1 vccd1 _06146_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16789_ _07026_ vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__clkbuf_4
X_18528_ net68 _09096_ vssd1 vssd1 vccd1 vccd1 _09097_ sky130_fd_sc_hd__nor2_4
XFILLER_0_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18459_ _02938_ _09023_ _03930_ vssd1 vssd1 vccd1 vccd1 _09024_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _04362_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__buf_6
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _03607_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ _01113_ _02099_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11421_ _01508_ _01513_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__or2b_1
XFILLER_0_34_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14140_ _04325_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__and2_1
X_11352_ _01442_ _01443_ _01375_ _01376_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10303_ _00380_ _00381_ _00395_ vssd1 vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14071_ _03199_ _04251_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__nand2_1
X_11283_ _01267_ _01365_ vssd1 vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13022_ _03106_ _03114_ _03061_ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__mux2_1
X_10234_ _00306_ _00307_ _00325_ vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__nand3_1
X_17830_ _03197_ _05625_ _08338_ _08341_ vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__a211o_1
X_10165_ _00254_ _00257_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__xnor2_1
X_17761_ _07751_ net145 vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__nand2_1
X_14973_ _05229_ _05236_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__or2_1
X_10096_ _00173_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__buf_2
X_16712_ _06951_ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__buf_2
X_13924_ _03962_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__inv_2
X_17692_ _08189_ _08190_ vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__nand2_1
X_16643_ _07017_ _07048_ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ _00204_ _01866_ _04015_ vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__nand3_1
XFILLER_0_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12806_ _01465_ _01466_ _00854_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__a211o_1
X_16574_ _06749_ _06891_ _06970_ _06972_ vssd1 vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13786_ _03848_ _03782_ cla_inst.in1\[22\] vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__and3_1
X_10998_ _01089_ _01090_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18313_ _08864_ _08866_ vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__xnor2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15525_ _05836_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _02820_ _02828_ _02829_ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _08786_ _08790_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__nand2_1
X_15456_ _05761_ _01317_ _05449_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__and4b_1
XFILLER_0_72_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ _02759_ _02760_ vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ _04612_ _04616_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or3_2
XFILLER_0_53_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11619_ _01187_ _01188_ _01191_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__a21o_1
X_18175_ _07195_ _07861_ _07745_ _07604_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__o211a_1
X_15387_ _05530_ _05676_ _05687_ vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ _02683_ _02691_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ _02347_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14338_ _04423_ _04424_ _04542_ _04543_ vssd1 vssd1 vccd1 vccd1 _04544_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17057_ _07497_ _07498_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__xnor2_2
X_14269_ _04461_ _04462_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__nand3_4
XFILLER_0_150_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ _02476_ _00167_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__and2_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _08363_ _08450_ _08481_ vssd1 vssd1 vccd1 vccd1 _08482_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11970_ _02022_ _02016_ _02021_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__nor3_1
X_10921_ _00998_ _00999_ _01013_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__a21o_2
X_13640_ _03778_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__nor2_1
X_10852_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel net209 _03388_
+ _04493_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _03703_ _03704_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nor2_1
X_10783_ _00870_ _00875_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__and2b_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15310_ _05503_ _05506_ _05603_ vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__a21oi_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _02604_ _02613_ net137 _02614_ vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _06664_ vssd1 vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ _05320_ _05439_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__and2_1
X_12453_ _05638_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel _07581_
+ _05562_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11404_ _01494_ _01495_ _01451_ _01444_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15172_ _05444_ _05451_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12384_ _05834_ _00357_ _07657_ _02476_ vssd1 vssd1 vccd1 vccd1 _02477_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14123_ _04302_ _04117_ _04308_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o21a_1
X_11335_ _01426_ _01427_ vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__xnor2_2
X_18931_ clknet_4_12_0_clk _00085_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[17\] sky130_fd_sc_hd__dfxtp_2
X_11266_ _01356_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__clkbuf_8
X_14054_ _04061_ _04060_ vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__or2b_1
X_10217_ _08724_ _00309_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13005_ _02489_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__buf_4
X_18862_ clknet_4_5_0_clk net288 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__dfxtp_1
X_11197_ _00967_ _01274_ _01288_ _01289_ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__o211a_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17813_ _08253_ _08254_ _08323_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__nand3_1
X_10148_ _07624_ _00240_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__xnor2_1
X_18793_ _09304_ vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17744_ _08225_ _08229_ _08248_ _06723_ _01671_ vssd1 vssd1 vccd1 vccd1 _09395_ sky130_fd_sc_hd__o32a_1
X_14956_ _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__xor2_1
X_10079_ _00171_ vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__buf_4
X_13907_ _04068_ _04071_ vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__nand2_1
X_17675_ _08057_ _08058_ vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__or2_1
X_14887_ _05021_ _05023_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__nand2_1
X_16626_ _07028_ _07029_ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__xnor2_1
X_13838_ _03805_ _03807_ _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16557_ _04449_ _04471_ _03184_ vssd1 vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o21a_1
X_13769_ _03916_ _03917_ _03919_ _03921_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15508_ _05813_ _05817_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16488_ _06878_ _06879_ _00194_ vssd1 vssd1 vccd1 vccd1 _06880_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18227_ _08739_ _08749_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__and2b_1
X_15439_ _02998_ _03153_ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18158_ _07751_ _08150_ _08625_ _08540_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__a31o_1
X_17109_ _07554_ _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__xnor2_1
X_18089_ _00558_ _07390_ _08621_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09931_ _08746_ vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _06982_ _07962_ _07951_ _07995_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__nand4_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _07243_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__buf_4
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _05682_ _04700_ _01211_ _01212_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__a31o_1
X_11051_ _01134_ _01143_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _07482_ _07908_ _09339_ _09340_ vssd1 vssd1 vccd1 vccd1 _09345_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14810_ _05056_ _05057_ _05058_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__and3_1
X_15790_ _06097_ _06123_ vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or2_1
X_14741_ _04975_ _04976_ _04981_ vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__a21o_1
Xwb_buttons_leds_151 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_151/HI led_enb[0] sky130_fd_sc_hd__conb_1
X_11953_ _01106_ _00515_ _02044_ _02045_ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__or4_4
Xwb_buttons_leds_162 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_162/HI led_enb[11] sky130_fd_sc_hd__conb_1
XFILLER_0_98_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10904_ _00990_ _00996_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__and2_1
X_17460_ _07936_ _07937_ vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__xnor2_2
X_14672_ _00125_ _00443_ _05050_ _00151_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11884_ _01871_ _01888_ _01889_ _01887_ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16411_ _06508_ _06783_ _06784_ _06796_ vssd1 vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__a31o_1
X_13623_ _03758_ _03759_ net226 _03754_ vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__a211o_1
X_10835_ _03771_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel
+ cla_inst.in2\[16\] vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17391_ _07860_ _07862_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16342_ _06721_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__clkbuf_4
X_13554_ _03685_ _03686_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__or2_1
X_10766_ _00857_ _00858_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_335 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12505_ _02595_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16273_ _06559_ _06583_ _06584_ _06608_ _06647_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__o311a_1
X_13485_ _00294_ cla_inst.in1\[24\] _05693_ _04504_ vssd1 vssd1 vccd1 vccd1 _03611_
+ sky130_fd_sc_hd__a22o_1
X_10697_ _04548_ _04482_ vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__nand2_2
XFILLER_0_82_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18012_ _07035_ _07933_ _08538_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__or3b_2
X_15224_ _05428_ _05396_ _05509_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12436_ _02471_ _02528_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15155_ _02987_ _03456_ _00513_ _02985_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12367_ _02452_ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__or3_1
X_14106_ _04558_ _09248_ _04288_ _04289_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__and4_1
X_11318_ _01410_ _01329_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__or2_1
X_15086_ _05237_ _05359_ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__xnor2_1
X_12298_ _02295_ _02298_ _02297_ vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__o21ai_1
X_14037_ _04212_ _04213_ _03997_ _04173_ vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__a211oi_1
X_11249_ cla_inst.in2\[24\] _00174_ _00871_ _09179_ vssd1 vssd1 vccd1 vccd1 _01342_
+ sky130_fd_sc_hd__nand4_1
X_18914_ clknet_4_9_0_clk _00068_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_129_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18845_ clknet_4_1_0_clk net274 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__dfxtp_1
X_18776_ _09290_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__buf_1
X_15988_ _02977_ _00134_ vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__or2_2
X_17727_ _02987_ _06511_ _01671_ vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14939_ _05199_ _05077_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _02200_ _06891_ vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16609_ _02829_ _02820_ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__xor2_1
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17589_ _08065_ _08078_ vssd1 vssd1 vccd1 vccd1 _08079_ sky130_fd_sc_hd__xor2_1
XFILLER_0_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 net100 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold111 _00011_ vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold122 net88 vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _00004_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _00014_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 op_code\[3\] vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_2
X_09914_ _04438_ _05388_ _05497_ _04646_ vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _07788_ _07384_ _07810_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__and3_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07069_ sky130_fd_sc_hd__buf_6
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ _00700_ _00701_ _00711_ vssd1 vssd1 vccd1 vccd1 _00713_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10551_ _05453_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__buf_4
XFILLER_0_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13270_ _03224_ _03225_ _03236_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__nor3_1
X_10482_ _00559_ _00574_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _02302_ _02304_ _02305_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__nor3_1
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12152_ _05584_ net206 _00179_ _05562_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11103_ _01193_ _01194_ _01195_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12083_ _02175_ _01999_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__nor2_1
X_16960_ _06571_ _06653_ _07194_ _07290_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__or4_2
X_11034_ _07232_ _07254_ _05333_ _05039_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__nand4_2
X_15911_ _06244_ _06253_ vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__or2_1
X_16891_ _07218_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__clkbuf_4
X_18630_ net310 _09097_ _09177_ _09176_ vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__o211a_1
X_15842_ _06128_ _06131_ vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__nand2_1
X_18561_ net311 _09098_ _09130_ _09126_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__o211a_1
X_15773_ _06104_ _06106_ vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__and2_1
X_12985_ _03066_ _03076_ _03077_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17512_ _07970_ _07994_ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__xnor2_1
X_14724_ _04924_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__inv_2
X_11936_ _01081_ _03826_ _03399_ _01082_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__a22o_1
X_18492_ _02939_ net115 _02960_ vssd1 vssd1 vccd1 vccd1 _09060_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17443_ _03080_ _03062_ _06724_ _03536_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__a31o_1
X_14655_ _04888_ _04889_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11867_ _01946_ _01959_ vssd1 vssd1 vccd1 vccd1 _01960_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13606_ _03527_ _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nand2_1
X_10818_ cla_inst.in2\[17\] ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel
+ _00179_ _03520_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__a22o_1
X_17374_ _07042_ _07721_ _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__o21ba_1
X_14586_ _04812_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__xnor2_1
X_11798_ _01704_ _01705_ _01706_ _01642_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ _06701_ _06703_ _03060_ vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13537_ _03426_ _03428_ _03666_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__or3b_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10749_ _06971_ _06722_ _07951_ _07995_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16256_ _06621_ _06628_ _03099_ vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__mux2_1
X_13468_ _03589_ net225 _03588_ vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_140_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15207_ _05374_ _05373_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12419_ _02414_ _02511_ vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16187_ _06477_ _03029_ _06543_ _06546_ _06553_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__o32a_2
X_13399_ _03469_ _03470_ _03514_ _03515_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _05407_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__or2_1
X_15069_ _05339_ _05340_ vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09630_ _05322_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__buf_4
X_18828_ net27 net28 _09109_ _09330_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09561_ _04668_ _04722_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__and2b_1
X_18759_ _00644_ net36 _09276_ vssd1 vssd1 vccd1 vccd1 _09277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09492_ _03706_ _03957_ _03946_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09828_ _07537_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__clkbuf_4
X_09759_ _06526_ _06537_ _04973_ _06191_ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__o211ai_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _02860_ _02861_ _02862_ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__or3b_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _03782_ _09179_ _07581_ _03848_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _03321_ _04591_ _01005_ _00112_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _00204_ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__buf_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10603_ _00491_ _00535_ net164 _00695_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__a211oi_4
X_14371_ _04577_ _04578_ vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__nor2_2
XFILLER_0_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _01673_ _01675_ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _02983_ _02257_ _03181_ _06467_ _06468_ vssd1 vssd1 vccd1 vccd1 _06469_ sky130_fd_sc_hd__o311a_1
X_13322_ _03408_ _03409_ _03429_ _03430_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__nand4_4
XFILLER_0_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10534_ _05017_ _05964_ _00624_ _00625_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a22o_1
X_17090_ _07533_ _07534_ vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16041_ _02998_ _04647_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__or2_1
XFILLER_0_134_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ _03355_ _03357_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__and2_1
X_10465_ _00557_ vssd1 vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12204_ _02274_ _02296_ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__xor2_1
X_10396_ _00467_ _00486_ _00487_ _00488_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__nand4_2
X_13184_ _03282_ _03283_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__xor2_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12135_ _02224_ _02225_ _02227_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__or3_2
X_17992_ _04630_ _06392_ _06391_ vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__a21oi_1
X_16943_ _03198_ _04559_ _07365_ _07375_ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__a211o_1
X_12066_ _02136_ _02137_ _02154_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__a211oi_1
X_11017_ _01107_ _01109_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__and2_1
X_16874_ _07298_ _07299_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__nand2_1
X_15825_ _03016_ _03072_ _06091_ _06090_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__a31o_1
X_18613_ net281 _09157_ _09167_ _09162_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__o211a_1
X_18544_ net13 net2 net24 vssd1 vssd1 vccd1 vccd1 _09115_ sky130_fd_sc_hd__or3b_4
X_15756_ _03007_ _03142_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12968_ _03060_ vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14707_ _04691_ _04692_ _04816_ _04817_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__and4b_1
XFILLER_0_75_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11919_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ net207
+ _00179_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__and4_1
X_18475_ _09038_ _09040_ vssd1 vssd1 vccd1 vccd1 _09041_ sky130_fd_sc_hd__xnor2_1
X_15687_ _05938_ _05941_ _06012_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__a21oi_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__buf_2
XFILLER_0_129_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17426_ _07900_ _07901_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__and2b_1
X_14638_ _07515_ _01962_ _01575_ _03008_ vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__a22o_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17357_ _07657_ net168 _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__and3_1
X_14569_ _04775_ _04794_ _04795_ vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__nor3_2
XFILLER_0_83_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16308_ _02980_ _01503_ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17288_ _06871_ _07032_ _00213_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_70_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16239_ _03064_ _06609_ _03089_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09613_ _05290_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__buf_4
X_09544_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04548_ sky130_fd_sc_hd__buf_4
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09475_ _03782_ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10250_ _07232_ _07254_ cla_inst.in1\[28\] _07374_ vssd1 vssd1 vccd1 vccd1 _00343_
+ sky130_fd_sc_hd__and4_1
X_10181_ _09027_ _09341_ _09345_ _09343_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__or4b_4
XFILLER_0_100_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13940_ _04092_ _03945_ _04106_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__nor3_1
X_13871_ _04031_ _04032_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__nor2_2
XFILLER_0_69_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15610_ _05927_ _05928_ _05828_ _05893_ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__a211o_1
X_12822_ _02913_ _02914_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__and2_1
X_16590_ _06908_ _06910_ _06909_ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_96_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15541_ _05848_ _05854_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__or2_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12753_ _02529_ _02589_ _02844_ _02845_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__o31ai_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _01795_ _01796_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__and2_1
X_18260_ _08807_ _08808_ vssd1 vssd1 vccd1 vccd1 _08809_ sky130_fd_sc_hd__and2_1
X_15472_ _05778_ _05779_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__or2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12684_ _02710_ _02745_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__xor2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _07663_ _07666_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__xnor2_1
X_14423_ _04634_ _04636_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _07853_ _00461_ _01220_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18191_ _08655_ _08733_ vssd1 vssd1 vccd1 vccd1 _08734_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ _06889_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__buf_4
X_14354_ _03164_ _03163_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11566_ _06008_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13305_ _09311_ _03412_ _03413_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10517_ _00607_ _00608_ _00609_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__nand3_1
X_17073_ _06581_ _07516_ vssd1 vssd1 vccd1 vccd1 _07517_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14285_ _04484_ _04485_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__and2_1
XFILLER_0_150_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11497_ _06591_ _00210_ _03607_ _05399_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16024_ _06374_ _03107_ vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__nand2_1
X_13236_ _03297_ _03337_ _03338_ vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__nand3_4
X_10448_ _00386_ _00391_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13167_ _03263_ _03264_ _00634_ _00660_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__o211a_2
X_10379_ _08713_ _06732_ _00470_ _00471_ vssd1 vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__and4_2
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _05562_ _05584_ _04242_ net206 vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__and4_1
X_17975_ _08381_ _08396_ _08394_ vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__a21o_1
X_13098_ _03185_ _03190_ _02489_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__mux2_1
X_12049_ _02058_ _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__xnor2_1
X_16926_ _07289_ _00248_ _06673_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__or3_2
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16857_ _07256_ _07261_ _07262_ _07279_ _07281_ vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__a311o_1
X_15808_ _03054_ _03058_ _03050_ vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__mux2_1
X_16788_ _06652_ _06764_ _06944_ _07115_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15739_ _06068_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18527_ net34 net67 vssd1 vssd1 vccd1 vccd1 _09096_ sky130_fd_sc_hd__nand2_1
X_18458_ _02920_ _08985_ _02918_ vssd1 vssd1 vccd1 vccd1 _09023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17409_ _07881_ _07882_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18389_ _07743_ _08947_ vssd1 vssd1 vccd1 vccd1 _08948_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09527_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04362_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09458_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03607_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11420_ _01511_ _01512_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _01375_ _01376_ _01442_ _01443_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10302_ _00383_ _00394_ vssd1 vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14070_ _03539_ _04248_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__o21ai_1
X_11282_ _01362_ _01338_ _01363_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13021_ _03110_ _03113_ _03090_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__mux2_1
X_10233_ _00306_ _00307_ _00325_ vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__a21o_2
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10164_ _00255_ _00256_ vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__and2b_1
X_14972_ _05233_ _05234_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__xor2_1
X_10095_ _00186_ _00187_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__or2_1
X_17760_ _08263_ _08264_ vssd1 vssd1 vccd1 vccd1 _08265_ sky130_fd_sc_hd__xnor2_1
X_13923_ _03368_ _01678_ _04021_ vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__nand3_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16711_ _07119_ _07121_ vssd1 vssd1 vccd1 vccd1 _07122_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17691_ _07207_ _07649_ _07780_ _06947_ vssd1 vssd1 vccd1 vccd1 _08190_ sky130_fd_sc_hd__a22o_1
X_16642_ _07019_ _07046_ vssd1 vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__xnor2_1
X_13854_ _04013_ _04014_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__xnor2_1
X_12805_ _00824_ _00853_ _00852_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__a21oi_1
X_16573_ _06970_ _06972_ _06749_ _06891_ vssd1 vssd1 vccd1 vccd1 _06973_ sky130_fd_sc_hd__o211a_1
X_13785_ _03934_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__a21o_1
X_10997_ _06971_ _06689_ _01087_ _01088_ vssd1 vssd1 vccd1 vccd1 _01090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15524_ _02998_ _05652_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nand2_1
X_18312_ _08638_ _08787_ _07604_ _07859_ vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _02797_ _02795_ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18243_ _08786_ _08790_ vssd1 vssd1 vccd1 vccd1 _08791_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15455_ _07515_ _05758_ _05986_ _03008_ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__a22o_1
X_12667_ _02719_ _02725_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__xnor2_1
X_14406_ _03014_ _02124_ _04615_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ _01614_ _01616_ _01613_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__a21o_1
X_18174_ _07109_ _07859_ _08640_ _08639_ vssd1 vssd1 vccd1 vccd1 _08716_ sky130_fd_sc_hd__a31o_1
X_15386_ _05685_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ _02683_ _02684_ _02690_ vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__or3_1
XFILLER_0_41_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _00558_ _06437_ _07573_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__o21a_1
X_14337_ _04540_ _04541_ _04425_ _04382_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__o211a_1
X_11549_ _01564_ _01604_ _01640_ _01641_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17056_ _06764_ _07194_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__nor2_1
X_14268_ _04463_ _04466_ vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__xor2_2
XFILLER_0_122_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16007_ _02476_ _00167_ vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nor2_1
X_13219_ _00125_ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__clkbuf_4
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _04222_ _04225_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__and2b_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _08469_ _08480_ vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__xnor2_1
X_16909_ _07336_ _07337_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__and2_1
X_17889_ _08298_ _08309_ vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ _01007_ _01012_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel
+ net209 _03388_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__and4_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ _00148_ _00149_ _04154_ _00563_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__and4_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10782_ _00190_ _00192_ _00134_ _00108_ _00874_ vssd1 vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__a41o_1
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _02560_ _02562_ _02564_ _02558_ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__o31a_1
XFILLER_0_66_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15240_ _05443_ _05455_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__and2_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ _02494_ _02492_ _02493_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _01451_ _01444_ _01494_ _01495_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15171_ _05444_ _05451_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12383_ _00645_ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14122_ _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__xnor2_1
X_11334_ _00195_ _00702_ _00127_ _07559_ _01344_ vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__a41o_1
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14053_ _04230_ _04232_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__nor2_2
X_18930_ clknet_4_10_0_clk _00084_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[16\] sky130_fd_sc_hd__dfxtp_2
X_11265_ _01356_ _01357_ _01110_ vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13004_ _03093_ _03096_ _03090_ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__mux2_1
X_10216_ _00308_ vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18861_ clknet_4_7_0_clk net282 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__dfxtp_1
X_11196_ _01279_ _01287_ _01286_ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__o21ai_1
X_17812_ _08320_ _08321_ vssd1 vssd1 vccd1 vccd1 _08323_ sky130_fd_sc_hd__nand2_1
X_10147_ _00236_ _00239_ vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__xnor2_1
X_18792_ _09298_ _09302_ vssd1 vssd1 vccd1 vccd1 _09304_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14955_ _02985_ _02988_ _09311_ _08224_ _05105_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a41o_1
X_17743_ _07256_ _08234_ _08236_ _08247_ vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10078_ _04242_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__buf_4
X_13906_ _04068_ _04071_ vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__or2_1
X_14886_ _05032_ _05030_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__and2b_1
X_17674_ _08070_ _08072_ _08069_ vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__o21ai_1
X_13837_ _03792_ _03995_ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__xnor2_1
X_16625_ _06653_ _06874_ vssd1 vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__nor2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16556_ _06812_ _06529_ _06953_ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__or3_1
X_13768_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15507_ _00115_ _00339_ _05814_ _05815_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12719_ _02789_ _02811_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__or2b_1
XFILLER_0_72_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16487_ _06812_ _06529_ _06530_ vssd1 vssd1 vccd1 vccd1 _06879_ sky130_fd_sc_hd__or3_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13699_ _03843_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__xor2_1
X_15438_ _05741_ _05742_ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__nor2_1
X_18226_ _08750_ _08756_ _08772_ _06721_ _06776_ vssd1 vssd1 vccd1 vccd1 _09402_ sky130_fd_sc_hd__o32a_2
XFILLER_0_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15369_ _00591_ _05652_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__and3_1
X_18157_ _08662_ _08664_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__and2b_1
XFILLER_0_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17108_ _07443_ _07445_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__or2_1
X_18088_ _02259_ _07387_ _08621_ vssd1 vssd1 vccd1 vccd1 _08622_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ cla_inst.in1\[21\] vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17039_ _07458_ _07465_ _07479_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _07973_ cla_inst.in1\[23\] cla_inst.in1\[22\] _07984_ vssd1 vssd1 vccd1 vccd1
+ _07995_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07243_ sky130_fd_sc_hd__buf_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11050_ _01134_ _01135_ _01142_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__nand3_2
XFILLER_0_101_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10001_ _09027_ _09341_ _09342_ _09343_ vssd1 vssd1 vccd1 vccd1 _09344_ sky130_fd_sc_hd__and4bb_2
X_14740_ _04975_ _04976_ _04981_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__nand3_2
XFILLER_0_99_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11952_ _01575_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__clkinv_4
Xwb_buttons_leds_152 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_152/HI led_enb[1] sky130_fd_sc_hd__conb_1
Xwb_buttons_leds_163 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_163/HI o_wb_stall sky130_fd_sc_hd__conb_1
X_10903_ _00991_ _00995_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__xor2_2
X_14671_ _04747_ _04748_ _04746_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__o21ai_1
X_11883_ _01944_ _01973_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 _01976_ sky130_fd_sc_hd__or4_4
X_16410_ _02823_ _06785_ _06795_ vssd1 vssd1 vccd1 vccd1 _06796_ sky130_fd_sc_hd__o21ai_1
X_13622_ _03590_ _03754_ _03758_ net336 vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__o211ai_4
X_10834_ cla_inst.in2\[16\] ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _00927_ sky130_fd_sc_hd__and4_1
X_17390_ _06561_ _07124_ _07516_ _07861_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16341_ _06720_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13553_ _00203_ _01962_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10765_ _00162_ _00230_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12504_ _07352_ _00146_ _02595_ _02596_ vssd1 vssd1 vccd1 vccd1 _02597_ sky130_fd_sc_hd__nand4_2
XFILLER_0_137_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16272_ _03117_ _06630_ _06644_ _06645_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13484_ _03990_ _06062_ _03385_ _03384_ _00459_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__a32o_1
X_10696_ _00786_ _00787_ _00788_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15223_ _05428_ _05396_ _05509_ vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18011_ _07125_ _07706_ vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12435_ _02460_ _02472_ _02527_ vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15154_ _02985_ _03456_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__nand2_1
X_12366_ _02389_ _02457_ _02451_ _02456_ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__o211a_1
X_14105_ _04515_ _02188_ _00498_ _08169_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__nand4_1
XFILLER_0_22_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11317_ _01324_ _01326_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__and2b_1
X_15085_ _05350_ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ _02295_ _02297_ _02298_ vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__or3_1
X_14036_ _03997_ _04173_ _04212_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__o211a_1
X_18913_ clknet_4_8_0_clk _00067_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[31\] sky130_fd_sc_hd__dfxtp_1
X_11248_ _00203_ _01264_ vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18844_ clknet_4_0_0_clk net262 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__dfxtp_1
X_11179_ _01147_ _01148_ _01237_ vssd1 vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__a21oi_1
X_18775_ _09273_ _09289_ vssd1 vssd1 vccd1 vccd1 _09290_ sky130_fd_sc_hd__and2_1
X_15987_ _06332_ _06333_ _06334_ _02677_ vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__a31o_1
X_17726_ _02326_ _02467_ _08226_ _08228_ vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__a31oi_4
X_14938_ _04946_ vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17657_ _08151_ _08152_ vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__nand2_1
X_14869_ _05121_ _05122_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16608_ _06421_ _06996_ _06997_ _07005_ _07010_ vssd1 vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__a311o_1
X_17588_ _08076_ _08077_ vssd1 vssd1 vccd1 vccd1 _08078_ sky130_fd_sc_hd__or2_1
XFILLER_0_147_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _06826_ _06899_ vssd1 vssd1 vccd1 vccd1 _06935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18209_ _08676_ _08677_ _08675_ vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 _00029_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 net91 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _00018_ vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 net86 vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 net103 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _04646_ _04373_ _05333_ _05039_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _07799_ _07722_ vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__and2_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _07047_ vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__buf_4
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10550_ _00641_ _00642_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _00572_ _00573_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__and2_1
X_12220_ _02126_ _02128_ _02303_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__or3_1
XFILLER_0_60_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _05562_ _05584_ net206 _00179_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__and4_1
X_11102_ _01062_ _01067_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__xnor2_2
X_12082_ _02173_ _02174_ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__or2b_1
X_11033_ _01096_ _01124_ _01125_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__nand3_2
X_15910_ _06244_ _06253_ vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__nand2_1
X_16890_ _07315_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__nor2_1
X_15841_ _06178_ _06179_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__or2_2
XFILLER_0_99_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18560_ salida\[2\] _09114_ _09118_ salida\[34\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09130_ sky130_fd_sc_hd__a221o_1
X_15772_ _06026_ _06028_ _06103_ vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__or3_1
X_12984_ _02981_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__buf_4
X_17511_ _07974_ _07993_ vssd1 vssd1 vccd1 vccd1 _07994_ sky130_fd_sc_hd__xor2_1
X_14723_ _04934_ _04935_ vssd1 vssd1 vccd1 vccd1 _04964_ sky130_fd_sc_hd__and2_1
X_11935_ _01949_ _01957_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__xnor2_2
X_18491_ _06248_ _06413_ _06412_ _06328_ vssd1 vssd1 vccd1 vccd1 _09058_ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14654_ _00195_ _00702_ _06062_ _05257_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__and4_1
X_17442_ _06736_ _06729_ _06731_ _06726_ _02977_ _02981_ vssd1 vssd1 vccd1 vccd1 _07920_
+ sky130_fd_sc_hd__mux4_1
X_11866_ _01949_ net176 _01958_ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13605_ _03355_ _03528_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__or2b_1
XFILLER_0_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10817_ net227 net169 _04242_ _00179_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__nand4_2
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14585_ _03368_ _04647_ _04645_ _04813_ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__a31oi_2
X_17373_ _06957_ _07194_ _07290_ _06961_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__o22a_1
X_11797_ _01871_ _01887_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nand4_2
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13536_ _03426_ _03428_ _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__o21ba_1
X_16324_ _03152_ _06496_ _06702_ _06626_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__o211a_1
X_10748_ _08006_ _00837_ _00840_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16255_ _06627_ vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13467_ _03588_ _03589_ _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__or3_4
XFILLER_0_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00772_ sky130_fd_sc_hd__buf_6
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15206_ _05489_ _05490_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__xor2_2
XFILLER_0_125_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12418_ _02401_ _02413_ vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16186_ _03029_ _06420_ _06543_ _06552_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o31a_1
X_13398_ _03469_ _03470_ _03514_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__nand4_4
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15137_ _05411_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__nand2_2
X_12349_ _02372_ _02374_ _02375_ _02369_ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ _05331_ _05338_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__nand2_1
X_14019_ _04029_ _04037_ _04194_ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__a21o_1
X_18827_ net69 _09111_ net67 vssd1 vssd1 vccd1 vccd1 _09330_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _04668_ _04679_ _04711_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__or3_1
X_18758_ _09250_ vssd1 vssd1 vccd1 vccd1 _09276_ sky130_fd_sc_hd__buf_4
X_17709_ _08086_ _08096_ _08209_ vssd1 vssd1 vccd1 vccd1 _08210_ sky130_fd_sc_hd__a21bo_1
X_09491_ _03706_ _03946_ _03957_ vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__nand3_2
X_18689_ net44 _09189_ _09223_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09827_ _07515_ _07537_ _07570_ _07613_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__and4_1
X_09758_ _06819_ _06830_ _06852_ vssd1 vssd1 vccd1 vccd1 _06873_ sky130_fd_sc_hd__nand3_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _05997_ _06116_ vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__xnor2_4
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _03848_ _01151_ _09179_ _07581_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__and4_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11651_ _01743_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__inv_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ _00661_ net165 _00692_ _00693_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14370_ _04001_ _07733_ _04575_ _04576_ vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__o2bb2a_1
X_11582_ _07853_ _06482_ _01674_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__and3_2
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _03408_ _03409_ _03429_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10533_ _04558_ _05964_ _00624_ _00625_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__nand4_2
XFILLER_0_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _06391_ _06392_ _04630_ vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13252_ _03353_ _03354_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__nand2_1
X_10464_ _04012_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__buf_6
XFILLER_0_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _02277_ _02279_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13183_ _07091_ _00509_ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10395_ _00465_ _00466_ _00291_ _00431_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a211o_4
X_12134_ _02193_ _02226_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__nand2_1
X_17991_ _04630_ _06391_ _06392_ vssd1 vssd1 vccd1 vccd1 _08517_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16942_ _06680_ _07367_ _07369_ _07373_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__or4_1
X_12065_ _02154_ _02156_ _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__nor3_1
X_11016_ _07788_ _05975_ _01108_ vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__and3_2
X_16873_ _07200_ _07296_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__nand2_1
X_18612_ salida\[23\] _09159_ _09160_ salida\[55\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09167_ sky130_fd_sc_hd__a221o_1
X_15824_ _06115_ _06113_ vssd1 vssd1 vccd1 vccd1 _06162_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18543_ _09113_ vssd1 vssd1 vccd1 vccd1 _09114_ sky130_fd_sc_hd__buf_2
X_15755_ _06034_ _06058_ _06059_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__nand3_1
X_12967_ _02489_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14706_ _04942_ _04945_ vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__xor2_2
X_11918_ _01922_ _02010_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__xnor2_1
X_18474_ _03108_ _03760_ _08047_ _09039_ vssd1 vssd1 vccd1 vccd1 _09040_ sky130_fd_sc_hd__o31a_1
X_12898_ _00148_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__clkbuf_4
X_15686_ _05938_ _05941_ _06012_ vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17425_ _07821_ _07786_ _07899_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__or3b_2
XFILLER_0_27_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14637_ _03008_ _07515_ _01962_ _02124_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11849_ _01841_ _01882_ _01883_ _01881_ vssd1 vssd1 vccd1 vccd1 _01942_ sky130_fd_sc_hd__a22o_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14568_ _04776_ _04664_ _04793_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17356_ _04034_ _06889_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__and2_1
XFILLER_0_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16307_ _06332_ _06545_ _06681_ _01503_ _06683_ vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13519_ _03622_ _03623_ _03646_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__and3_1
X_14499_ _04712_ _04713_ _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__nand3_1
X_17287_ _07302_ _07303_ _07130_ _07126_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__or4_1
XFILLER_0_153_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16238_ _09263_ _03074_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16169_ _03184_ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09612_ ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05290_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09543_ _04406_ _04526_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__or2_4
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09474_ _03771_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwire119 _03888_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__buf_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ _09348_ _00270_ _00271_ _00272_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__nand4_4
X_13870_ cla_inst.in2\[27\] cla_inst.in2\[26\] _03903_ _03914_ vssd1 vssd1 vccd1 vccd1
+ _04032_ sky130_fd_sc_hd__and4_2
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12821_ _02911_ _02912_ _01492_ _01494_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__a211o_2
X_15540_ _05851_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _02528_ _02587_ _02471_ vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__o21ai_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _01764_ _01792_ _01794_ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__or3_1
X_15471_ _05776_ _05777_ _05674_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__o21a_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _02744_ _02752_ _02775_ vssd1 vssd1 vccd1 vccd1 _02776_ sky130_fd_sc_hd__and3_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _00253_ _00460_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__nand2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ _06750_ _07665_ _07543_ _07541_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__a31oi_2
X_11634_ _01221_ _01693_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18190_ _08731_ _08732_ vssd1 vssd1 vccd1 vccd1 _08733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ _03138_ _03147_ _03185_ _03190_ _03062_ _02979_ vssd1 vssd1 vccd1 vccd1 _04560_
+ sky130_fd_sc_hd__mux4_1
X_17141_ _06937_ _07314_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__nor2_1
X_11565_ _06982_ _01005_ _01656_ _01657_ vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13304_ _06051_ _09303_ _07733_ _06040_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ _00433_ _00434_ _00432_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__a21bo_1
X_17072_ _07410_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__clkbuf_4
X_14284_ _04309_ _04473_ _04483_ vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__or3_1
XFILLER_0_24_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11496_ _01587_ _01588_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13235_ _03335_ _03336_ _00690_ _00692_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_21_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16023_ _06374_ _03107_ vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__or2_1
X_10447_ _00383_ _00394_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _00634_ _00660_ _03263_ _03264_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a211oi_2
X_10378_ _05508_ _05464_ _00308_ _05964_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__nand4_1
X_12117_ _02181_ _02204_ _02209_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__or3_1
X_17974_ _08497_ _08498_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__and2_1
X_13097_ _03187_ _03189_ _03047_ vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__mux2_1
X_12048_ _01905_ _02060_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__nand2_1
X_16925_ _07289_ _07355_ _00248_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16856_ _02776_ _02834_ _07280_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15807_ _03034_ _06143_ _04247_ vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16787_ _07203_ _07204_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__nor2_1
X_13999_ _03985_ _03999_ vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18526_ _09074_ _09081_ _09095_ _06721_ _00516_ vssd1 vssd1 vccd1 vccd1 _09410_ sky130_fd_sc_hd__o32a_1
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _05994_ _06067_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18457_ _09020_ _09021_ vssd1 vssd1 vccd1 vccd1 _09022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15669_ _05920_ _05993_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17408_ _07731_ _07767_ _07880_ vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18388_ _03760_ _08047_ vssd1 vssd1 vccd1 vccd1 _08947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _04853_ _06371_ _06370_ vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19009_ clknet_4_1_0_clk _09376_ vssd1 vssd1 vccd1 vccd1 salida\[62\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _04340_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__buf_6
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _03366_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ _01440_ _01441_ _01337_ _01377_ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10301_ _00384_ _00393_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__xnor2_1
X_11281_ _01371_ _01372_ _01370_ _01373_ vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13020_ _03023_ _03112_ vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__nand2_1
X_10232_ _00316_ _00324_ vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10163_ _00175_ _03618_ _00218_ _00173_ vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _00362_ _05856_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__nand2_1
X_10094_ _00170_ _00172_ _00182_ _00185_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__a22oi_1
X_16710_ _07022_ _07027_ _07120_ vssd1 vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__a21oi_1
X_13922_ _04018_ _04020_ vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__or2b_1
X_17690_ _07302_ _07303_ _07516_ _07511_ vssd1 vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__or4_1
XFILLER_0_88_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16641_ _07021_ _07045_ vssd1 vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__xnor2_1
X_13853_ _03839_ _03842_ _03840_ vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16572_ _06882_ _06883_ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__and2b_1
X_13784_ _03934_ _03936_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__nand3_1
X_10996_ _06971_ _06689_ _01087_ _01088_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18311_ _08862_ _08863_ vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__nor2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15523_ _05832_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__nand2_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12735_ _02826_ _02827_ vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _08787_ _08788_ vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__xor2_1
X_15454_ _03008_ _07515_ _05758_ _05986_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _02754_ _02756_ _02757_ _02758_ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__or4_2
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14405_ _04614_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__inv_2
X_11617_ _01610_ _01619_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__o211ai_2
X_18173_ _08712_ _08714_ vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__or2_1
X_15385_ _05677_ _05684_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ _02687_ _02688_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17124_ _06424_ _06438_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nor2_1
X_14336_ _04425_ _04382_ _04540_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__a211oi_2
X_11548_ _01621_ _01639_ _01638_ vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17055_ _06657_ _07396_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ _08724_ _04067_ _01570_ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ _00681_ _00682_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__nor2_1
X_16006_ _06354_ _06355_ _01829_ vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14198_ _04387_ _04388_ _04389_ vssd1 vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__o21a_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _03245_ _03246_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__xor2_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _08470_ _08479_ vssd1 vssd1 vccd1 vccd1 _08480_ sky130_fd_sc_hd__xnor2_1
X_16908_ _06665_ _07332_ _07335_ vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__o21ai_1
X_17888_ _08403_ _08404_ vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__or2_1
X_16839_ _07259_ _07260_ vssd1 vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18509_ _00516_ _09076_ _06512_ vssd1 vssd1 vccd1 vccd1 _09077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10850_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _03903_ vssd1
+ vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09509_ _04099_ _04132_ _04143_ _04154_ vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__and4_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _00169_ _00180_ _00872_ _00873_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__and4_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _02605_ _02606_ _02612_ vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__or3_4
XFILLER_0_149_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12451_ _02498_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ _01492_ _01493_ _01452_ _01453_ vssd1 vssd1 vccd1 vccd1 _01495_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15170_ _05448_ _05450_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__or2_1
XFILLER_0_117_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12382_ _02425_ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_90 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14121_ _02533_ _03456_ _04134_ _04133_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11333_ _00874_ _01425_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14052_ _04228_ _04229_ _04089_ _04090_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__o211a_1
X_11264_ _09354_ vssd1 vssd1 vccd1 vccd1 _01357_ sky130_fd_sc_hd__buf_4
X_13003_ _03040_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__nand2_1
X_10215_ _05693_ vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18860_ clknet_4_7_0_clk net284 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__dfxtp_1
X_11195_ _01279_ _01286_ _01287_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17811_ _08318_ _08319_ vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__or2_1
X_10146_ _00237_ _00238_ vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__and2b_1
X_18791_ _03368_ net47 _09301_ vssd1 vssd1 vccd1 vccd1 _09302_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _06421_ _08237_ _08238_ _08240_ _08245_ vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__a311o_1
X_14954_ _05214_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__xnor2_1
X_10077_ _00169_ vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13905_ _03741_ _03746_ _03902_ _04070_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__o31a_1
X_17673_ _08167_ _08170_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__xor2_1
X_14885_ _04877_ _05029_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__and2b_1
X_16624_ _07022_ _07027_ vssd1 vssd1 vccd1 vccd1 _07028_ sky130_fd_sc_hd__xnor2_1
X_13836_ _03993_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16555_ _03804_ _03826_ _03399_ vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10979_ _01069_ _01070_ _01071_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__a21o_1
X_13767_ _02972_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__clkbuf_4
X_15506_ _05816_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__inv_2
X_12718_ _02786_ _02787_ _02788_ _02782_ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ _03184_ _06529_ net150 _03313_ vssd1 vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13698_ _00253_ _01575_ _03680_ _03679_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18225_ _06426_ _06447_ _08758_ _08771_ vssd1 vssd1 vccd1 vccd1 _08772_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_143_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15437_ _02993_ _02996_ _00495_ _00339_ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__and4_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12649_ _02733_ _02739_ _02740_ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18156_ _08695_ vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__inv_2
X_15368_ _05665_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17107_ _07552_ _07553_ vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__xnor2_1
X_14319_ _04514_ _04522_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__xnor2_1
X_18087_ _08619_ _08620_ vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__and2_1
X_15299_ _05590_ _05591_ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17038_ _03921_ _03120_ _04826_ _07468_ _07478_ vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09860_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07984_ sky130_fd_sc_hd__buf_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _07221_ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__buf_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ clknet_4_6_0_clk _09385_ vssd1 vssd1 vccd1 vccd1 salida\[42\] sky130_fd_sc_hd__dfxtp_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10000_ _09005_ _09016_ net166 _06906_ vssd1 vssd1 vccd1 vccd1 _09343_ sky130_fd_sc_hd__a211o_1
X_09989_ cla_inst.in1\[29\] vssd1 vssd1 vccd1 vccd1 _09303_ sky130_fd_sc_hd__clkbuf_4
X_11951_ _04700_ vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__clkinv_4
Xwb_buttons_leds_153 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_153/HI led_enb[2] sky130_fd_sc_hd__conb_1
X_10902_ _05497_ _00993_ _00994_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__a21bo_1
X_14670_ _00115_ _05888_ _04784_ _04783_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__a31o_1
X_11882_ _01943_ _01919_ _01941_ vssd1 vssd1 vccd1 vccd1 _01975_ sky130_fd_sc_hd__and3_1
X_13621_ _03755_ _03756_ _03757_ vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__a21o_1
X_10833_ _00918_ _00919_ _00924_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16340_ _02966_ _06459_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__or2_2
X_10764_ _00828_ _00851_ _00827_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__a21bo_2
X_13552_ _03682_ _03683_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _07973_ _00196_ _01031_ _07221_ vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__a22o_1
X_13483_ _03398_ _03400_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__nand2_1
X_16271_ _03036_ _02965_ _06422_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__or3_4
X_10695_ _04427_ _03739_ _03804_ _04635_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18010_ _08535_ _08536_ vssd1 vssd1 vccd1 vccd1 _08537_ sky130_fd_sc_hd__xnor2_1
X_15222_ _05506_ _05507_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__nand2_1
X_12434_ _02523_ _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15153_ _02987_ _00665_ _05317_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__and3_1
X_12365_ _02451_ _02456_ _02389_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_50_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14104_ _04438_ _07722_ _08169_ _04515_ vssd1 vssd1 vccd1 vccd1 _04288_ sky130_fd_sc_hd__a22o_1
X_11316_ _01407_ _01408_ vssd1 vssd1 vccd1 vccd1 _01409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15084_ _05351_ _05357_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _02385_ _02387_ _02388_ vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__nor3_1
X_14035_ _04210_ _04211_ _04191_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__o21ai_1
X_18912_ clknet_4_8_0_clk _00066_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[30\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11247_ _00204_ _01248_ _01259_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18843_ clknet_4_0_0_clk net253 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11178_ _01251_ _01270_ vssd1 vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__xnor2_1
X_10129_ _00220_ _00221_ vssd1 vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__or2_1
X_18774_ _06374_ net41 _09276_ vssd1 vssd1 vccd1 vccd1 _09289_ sky130_fd_sc_hd__mux2_1
X_15986_ _07711_ _00357_ _07657_ _02505_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_12 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17725_ _03930_ _08227_ vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__nand2_1
X_14937_ _05196_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _02044_ _06755_ _06764_ _07933_ vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__or4_1
X_14868_ _04992_ _04998_ vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__and2_1
X_16607_ _06543_ _06434_ _07006_ _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__a31o_1
X_13819_ _03974_ _03975_ vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__xor2_2
X_17587_ _08074_ _08075_ _08066_ vssd1 vssd1 vccd1 vccd1 _08077_ sky130_fd_sc_hd__o21a_1
X_14799_ _05045_ _05046_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16538_ _06898_ _06897_ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16469_ _03120_ _03565_ _06850_ _06859_ vssd1 vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18208_ _08751_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__and2b_1
XFILLER_0_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ _08675_ _08676_ _08677_ vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold102 net93 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _00021_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 net99 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _00016_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 _00032_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _04558_ _05486_ vssd1 vssd1 vccd1 vccd1 _08550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ ApproximateM_inst.lob_16.lob2.mux.sel vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__clkbuf_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _07036_ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__clkbuf_8
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ _00571_ _00560_ _00561_ vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12150_ _06993_ _00166_ _02241_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__a31o_1
X_11101_ _01175_ _01171_ vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__or2b_1
X_12081_ _02169_ _02081_ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _06971_ _05246_ _01094_ _01095_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__a22o_1
X_15840_ _06121_ _06124_ _06177_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__and3_1
X_15771_ _06026_ _06028_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12983_ _03070_ _03075_ _03050_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__mux2_1
X_17510_ _07991_ _07992_ vssd1 vssd1 vccd1 vccd1 _07993_ sky130_fd_sc_hd__and2b_1
X_14722_ _00592_ _04900_ _04899_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__and3_1
X_18490_ _06836_ _09055_ _09056_ vssd1 vssd1 vccd1 vccd1 _09057_ sky130_fd_sc_hd__or3_1
X_11934_ _02009_ _02024_ _02026_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17441_ _06375_ _06545_ _07917_ _03108_ vssd1 vssd1 vccd1 vccd1 _07918_ sky130_fd_sc_hd__a22o_1
X_14653_ _00191_ _06094_ _00460_ _00189_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11865_ _01953_ _01956_ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13604_ _03358_ _03359_ _03527_ _03528_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__and4_1
XFILLER_0_67_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10816_ _00772_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__buf_6
X_17372_ _07714_ _07715_ _07712_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__a21oi_1
X_14584_ _04643_ _04644_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__and2b_1
X_11796_ _01885_ _01886_ _01881_ _01884_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_28_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16323_ _03047_ _06499_ vssd1 vssd1 vccd1 vccd1 _06702_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ _03660_ _03665_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10747_ _05671_ _00459_ _00838_ _00839_ _05388_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__a32oi_2
XFILLER_0_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16254_ _03152_ _06622_ _06625_ _06626_ vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__o211a_1
X_13466_ _03520_ _03498_ _05311_ cla_inst.in1\[17\] vssd1 vssd1 vccd1 vccd1 _03590_
+ sky130_fd_sc_hd__and4_4
X_10678_ cla_inst.in2\[19\] cla_inst.in2\[17\] ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _00771_ sky130_fd_sc_hd__and4_2
XFILLER_0_36_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15205_ _02999_ _00339_ vssd1 vssd1 vccd1 vccd1 _05490_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12417_ _02484_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__xnor2_1
X_16185_ _03027_ _06420_ _06549_ _06551_ _02779_ vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__a2111o_1
X_13397_ _03512_ _03513_ _03333_ _03335_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ _04409_ _05409_ _05413_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__o211a_4
X_12348_ _02435_ _02440_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15067_ _05331_ _05338_ vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__or2_1
X_12279_ _02260_ _02371_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__nor2_1
X_14018_ _04030_ _04036_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18826_ _09329_ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__clkbuf_1
X_18757_ _09275_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__buf_1
X_15969_ _03920_ _05095_ _06316_ vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__a21oi_2
X_17708_ _08097_ _08084_ vssd1 vssd1 vccd1 vccd1 _08209_ sky130_fd_sc_hd__or2b_1
X_09490_ _03553_ _03563_ _03695_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18688_ _01671_ _09183_ _09191_ vssd1 vssd1 vccd1 vccd1 _09223_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _08132_ _08133_ _06589_ vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09826_ _07602_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__clkbuf_8
X_09757_ _06819_ _06830_ _06852_ vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__a21o_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _06073_ _06105_ vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__and2b_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ cla_inst.in2\[20\] _07646_ _09354_ _00877_ vssd1 vssd1 vccd1 vccd1 _01743_
+ sky130_fd_sc_hd__a22o_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10601_ _00661_ _00662_ _00692_ _00693_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_36_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11581_ _00515_ _01671_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nor2_4
XFILLER_0_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ _04646_ _04438_ _08757_ _05246_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__nand4_2
X_13320_ _03426_ _03427_ _03254_ _03256_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10463_ _00554_ _00539_ _00540_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13251_ _03353_ _03354_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__or2_4
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ _02230_ _02282_ net129 _02294_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__a211oi_4
X_13182_ _07058_ _00502_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand2_1
X_10394_ _00484_ _00485_ _00482_ _00483_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__o211ai_4
X_12133_ _02190_ _02192_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__nand2_1
X_17990_ _08512_ _08513_ _08514_ vssd1 vssd1 vccd1 vccd1 _08516_ sky130_fd_sc_hd__a21o_1
X_12064_ _02070_ _02153_ _02148_ _02152_ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__a211oi_1
X_16941_ _02973_ _07370_ _07372_ _06484_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__o211a_1
X_11015_ _07799_ _05715_ vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__and2_4
X_16872_ _07200_ _07296_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__or2_1
X_18611_ net283 _09157_ _09165_ _09162_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__o211a_1
X_15823_ _06153_ _06160_ vssd1 vssd1 vccd1 vccd1 _06161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18542_ net24 _09110_ _09111_ vssd1 vssd1 vccd1 vccd1 _09113_ sky130_fd_sc_hd__nor3_2
X_15754_ _06061_ _06063_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__or2b_1
XFILLER_0_99_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12966_ _03054_ _03058_ _03050_ vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14705_ _04943_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11917_ _01924_ _01923_ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__nand2_1
X_18473_ _08999_ _09002_ vssd1 vssd1 vccd1 vccd1 _09039_ sky130_fd_sc_hd__nand2_1
X_15685_ _06010_ _06011_ vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__or2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _02985_ _02987_ _02988_ _02989_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__or4_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17424_ _07821_ _07786_ _07899_ vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__o21ba_2
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _03006_ _00716_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _01938_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__or3_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _07091_ _06753_ _07780_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14567_ _04776_ _04664_ _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21oi_4
X_11779_ _01844_ _01871_ vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16306_ _06427_ _06429_ _06682_ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__a21oi_1
X_13518_ _03622_ _03623_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_125_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17286_ _07747_ _07748_ vssd1 vssd1 vccd1 vccd1 _07749_ sky130_fd_sc_hd__nand2_1
X_14498_ _04716_ _04717_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16237_ _03117_ _03035_ _03121_ _06590_ _06607_ vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__o311a_1
XFILLER_0_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13449_ _03570_ _03157_ _02983_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16168_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel sel_op\[0\] vssd1
+ vssd1 vccd1 vccd1 _06533_ sky130_fd_sc_hd__or2b_1
XFILLER_0_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15119_ _05310_ _05395_ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16099_ _06415_ _06416_ _06421_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__a31o_1
X_09611_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05279_ sky130_fd_sc_hd__buf_4
X_18809_ _01417_ net53 _09301_ vssd1 vssd1 vccd1 vccd1 _09316_ sky130_fd_sc_hd__mux2_1
X_09542_ _04438_ _04460_ _04482_ _04515_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09473_ ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel vssd1 vssd1 vccd1 vccd1
+ _03771_ sky130_fd_sc_hd__buf_6
XFILLER_0_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _07080_ _07406_ _07112_ _07047_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__a22o_1
X_12820_ _01492_ _01494_ _02911_ _02912_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _02633_ _02671_ _02842_ _02843_ _02590_ vssd1 vssd1 vccd1 vccd1 _02844_ sky130_fd_sc_hd__o32a_4
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _01764_ _01792_ _01794_ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__o21ai_2
X_15470_ _05674_ _05776_ _05777_ vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__nor3_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _02762_ _02773_ _02774_ vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _04632_ _04633_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__nor2_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _01722_ _01723_ _01724_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17140_ _07485_ _07491_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14352_ _03921_ _04557_ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__nor2_1
X_11564_ _01082_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _01657_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13303_ _06040_ _06051_ _07733_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__and3_1
X_10515_ _00604_ _00605_ _00606_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a21o_1
X_17071_ _07512_ _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__and2b_1
XFILLER_0_150_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14283_ _04309_ _04473_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__o21ai_1
X_11495_ _01571_ _01570_ vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16022_ _04034_ vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__clkbuf_4
X_10446_ _00384_ _00393_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__and2b_1
X_13234_ _00690_ _00692_ _03335_ _03336_ vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__a211o_2
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _05366_ _05704_ _05606_ _05410_ vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13165_ _03240_ _03241_ _03261_ _03262_ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__and4_2
X_12116_ _09219_ _02205_ _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__a21oi_1
X_17973_ _08449_ _08400_ _08495_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__or3_1
X_13096_ _01863_ _03188_ _03022_ vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__o21a_1
X_12047_ _02059_ _09354_ _02139_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__nand3_1
X_16924_ _06673_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16855_ _02776_ _02834_ _02968_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__a21oi_1
X_15806_ _03910_ _03924_ _02981_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__mux2_1
X_16786_ _07107_ _07202_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__and2_1
X_13998_ _04024_ _04041_ _04042_ vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18525_ _06421_ _09082_ _09083_ _09090_ _09094_ vssd1 vssd1 vccd1 vccd1 _09095_ sky130_fd_sc_hd__a311o_1
XFILLER_0_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15737_ _05994_ _06067_ vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ _03025_ _03041_ _01674_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18456_ _08980_ _08982_ _08979_ vssd1 vssd1 vccd1 vccd1 _09021_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15668_ _02994_ _05652_ _05992_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__and3_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_180 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17407_ _07731_ _07767_ _07880_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__o21ai_1
X_14619_ _04841_ _04843_ _04848_ vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18387_ _08909_ _08910_ vssd1 vssd1 vccd1 vccd1 _08946_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15599_ _05916_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17338_ _04853_ _06370_ _06371_ vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__nand3_1
XFILLER_0_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17269_ _07718_ _07728_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008_ clknet_4_5_0_clk _09375_ vssd1 vssd1 vccd1 vccd1 salida\[61\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09525_ ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04340_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09456_ _03574_ _03432_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10300_ _00385_ _00392_ vssd1 vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__xor2_1
X_11280_ _01368_ _01369_ _01238_ _01273_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10231_ _00321_ _00323_ vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10162_ _00184_ _00183_ _03618_ _00171_ vssd1 vssd1 vccd1 vccd1 _00255_ sky130_fd_sc_hd__and4_1
X_14970_ _05231_ _05232_ vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__nor2_1
X_10093_ _00170_ _00172_ _00182_ _00185_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__and4_1
X_13921_ _04087_ vssd1 vssd1 vccd1 vccd1 _09381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ _07031_ _07044_ vssd1 vssd1 vccd1 vccd1 _07045_ sky130_fd_sc_hd__xnor2_1
X_13852_ _04010_ _04011_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _01483_ _01469_ _01484_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16571_ _06527_ _06877_ _06969_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__and3_1
X_13783_ _03755_ _03757_ _03756_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__a21bo_1
X_10995_ _07973_ _08746_ _06613_ _07984_ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18310_ _08785_ _08791_ _08861_ vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__and3_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15522_ _05833_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12734_ _02803_ _02819_ vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _07608_ _07861_ _08638_ vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ _03006_ _03044_ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__nand2_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12665_ _02721_ _02755_ vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__and2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14404_ _04614_ _01575_ _07537_ _04615_ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and4b_1
X_11616_ _01166_ _01177_ _01176_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_93_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18172_ _08629_ _08711_ _08698_ vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__and3_1
X_15384_ _05677_ _05684_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__or2_1
X_12596_ _02647_ _02686_ vssd1 vssd1 vccd1 vccd1 _02689_ sky130_fd_sc_hd__and2_1
X_17123_ _00787_ _06331_ _06365_ _07084_ _07571_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_142_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14335_ _04538_ _04539_ _04426_ _04385_ vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__o211a_1
X_11547_ _01621_ _01638_ _01639_ vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__nor3_4
X_17054_ _07494_ _07495_ vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__or2_1
X_14266_ _00644_ _04125_ _04130_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11478_ _00806_ _05290_ _00949_ _03421_ vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16005_ _02533_ _00214_ vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__or2_2
XFILLER_0_150_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13217_ _01356_ _00213_ _00728_ _00727_ vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a31o_1
X_10429_ _07635_ _00193_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__nand2_1
X_14197_ _04387_ _04388_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__nor3_1
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _05747_ _09311_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _02685_ _03170_ _03023_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__o21ai_1
X_17956_ _08477_ _08478_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__and2_1
X_16907_ _06665_ _07332_ _07335_ vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__or3_4
X_17887_ _08292_ _08348_ _08402_ vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__nor3_1
XFILLER_0_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16838_ _07259_ _07260_ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ _03916_ _06503_ _07185_ _06645_ vssd1 vssd1 vccd1 vccd1 _07186_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18508_ _06303_ _06416_ vssd1 vssd1 vccd1 vccd1 _09076_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18439_ _06277_ _09000_ _04995_ _07592_ _09001_ vssd1 vssd1 vccd1 vccd1 _09002_ sky130_fd_sc_hd__o311a_1
XFILLER_0_29_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09508_ _03410_ vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__buf_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10780_ cla_inst.in2\[23\] _00129_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ cla_inst.in2\[24\] vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _03388_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__clkbuf_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12450_ _02491_ _02497_ _02496_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _01452_ _01453_ _01492_ _01493_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12381_ _05747_ _00193_ _02473_ _02424_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_80 _07766_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_91 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _04303_ _04304_ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or2_1
X_11332_ _00169_ _00146_ _00872_ _00873_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14051_ _04089_ _04090_ _04228_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__a211oi_2
X_11263_ _09353_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__clkbuf_8
X_13002_ _00167_ _03094_ _02505_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__mux2_1
X_10214_ _08605_ _08626_ vssd1 vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__nand2_1
X_11194_ _01278_ _01275_ _01276_ vssd1 vssd1 vccd1 vccd1 _01287_ sky130_fd_sc_hd__and3_1
X_17810_ _08318_ _08319_ vssd1 vssd1 vccd1 vccd1 _08320_ sky130_fd_sc_hd__nand2_1
X_10145_ _09349_ _00181_ _00197_ _00109_ vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__a22o_1
X_18790_ _09250_ vssd1 vssd1 vccd1 vccd1 _09301_ sky130_fd_sc_hd__clkbuf_4
X_17741_ _06462_ _08242_ _08244_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__or3_1
X_14953_ _02986_ _09311_ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nand2_1
X_10076_ cla_inst.in2\[22\] vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__buf_2
X_13904_ _03900_ _03901_ _04069_ vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17672_ _08054_ _08061_ _08168_ vssd1 vssd1 vccd1 vccd1 _08170_ sky130_fd_sc_hd__a21bo_1
X_14884_ _05034_ vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16623_ _07613_ _06541_ _07026_ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__and3_1
X_13835_ _03989_ _03992_ _03986_ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_140 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _06427_ _06651_ _06951_ vssd1 vssd1 vccd1 vccd1 _06952_ sky130_fd_sc_hd__or3_1
XFILLER_0_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13766_ _03913_ _03918_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__nor2_1
X_10978_ _00990_ _00996_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15505_ _00107_ _07744_ _05814_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12717_ _02489_ _02779_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__or3b_1
X_16485_ _06567_ _06570_ _06807_ _00357_ vssd1 vssd1 vccd1 vccd1 _06877_ sky130_fd_sc_hd__o211a_1
X_13697_ _03841_ _03842_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18224_ _08762_ _08765_ _08769_ _08770_ vssd1 vssd1 vccd1 vccd1 _08771_ sky130_fd_sc_hd__and4b_1
X_15436_ _02996_ _00495_ _00339_ _02993_ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12648_ _02701_ _02703_ _02702_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18155_ _08665_ _08666_ vssd1 vssd1 vccd1 vccd1 _08695_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15367_ _05653_ _05585_ _05664_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ _02644_ _02645_ _02651_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__nand3_1
XFILLER_0_81_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17106_ _07324_ _07326_ _07436_ _07438_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__o31ai_2
X_14318_ _04516_ _04521_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__xnor2_1
X_18086_ _07313_ _07410_ _07486_ _07593_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15298_ _00591_ _03154_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__nand2_2
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17037_ _06425_ _06437_ _07469_ _07473_ _07477_ vssd1 vssd1 vccd1 vccd1 _07478_ sky130_fd_sc_hd__o311a_1
X_14249_ _04442_ _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07221_ sky130_fd_sc_hd__buf_4
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ clknet_4_6_0_clk _09384_ vssd1 vssd1 vccd1 vccd1 salida\[41\] sky130_fd_sc_hd__dfxtp_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _07042_ _08260_ vssd1 vssd1 vccd1 vccd1 _08460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _09271_ _09279_ vssd1 vssd1 vccd1 vccd1 _09295_ sky130_fd_sc_hd__or2_1
X_11950_ _02028_ _02041_ vssd1 vssd1 vccd1 vccd1 _02043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xwb_buttons_leds_154 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_154/HI led_enb[3] sky130_fd_sc_hd__conb_1
X_10901_ _05638_ _05028_ _04569_ _00992_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ _01971_ _01972_ _01960_ _01968_ vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__o211a_1
X_13620_ _03755_ _03756_ _03757_ vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__nand3_2
X_10832_ _00918_ _00919_ _00924_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13551_ _00170_ _00715_ _03475_ _03474_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__a31o_1
X_10763_ _00823_ _00854_ _08311_ _00855_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__o211a_4
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12502_ _07036_ _07069_ _00130_ _00871_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__nand4_2
XFILLER_0_125_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16270_ _06636_ _06643_ _03538_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__o21a_1
X_13482_ _03603_ _03604_ _03605_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10694_ _04427_ _03804_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__nand2_4
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _05387_ _05505_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__or2_1
X_12433_ _02524_ _02523_ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__nor3_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ _05326_ _05328_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12364_ _02385_ _02388_ _02387_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14103_ _04103_ _04104_ _04102_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_50_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ net139 _01405_ _01306_ _01304_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__o211a_1
X_15083_ _05354_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12295_ _02282_ _02384_ _02352_ net323 vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_120_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14034_ _04191_ _04210_ _04211_ vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__or3_2
X_18911_ clknet_4_10_0_clk _00065_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[29\] sky130_fd_sc_hd__dfxtp_1
X_11246_ _01241_ _01258_ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18842_ clknet_4_0_0_clk net251 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__dfxtp_1
X_11177_ _01252_ _01269_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__xnor2_1
X_10128_ _00170_ _00206_ _00216_ _00219_ vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__o2bb2a_1
X_18773_ _09288_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__clkbuf_1
X_15985_ _07711_ _00357_ vssd1 vssd1 vccd1 vccd1 _06333_ sky130_fd_sc_hd__or2_2
X_10059_ _00149_ _00131_ _00127_ _00151_ vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a22o_1
X_14936_ _05194_ _05195_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__nand2_1
X_17724_ _02467_ _08226_ _02326_ vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__a21o_1
X_14867_ _05119_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__or2_1
X_17655_ _02977_ _06753_ _07859_ _08150_ _06762_ vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__a32o_1
X_13818_ _03796_ _03798_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__nand2_1
X_16606_ _03537_ _03197_ _04076_ _06680_ _07008_ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__a311o_1
X_17586_ _08066_ _08074_ _08075_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__nor3_1
X_14798_ _05044_ _05043_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__or2b_1
X_16537_ _06933_ vssd1 vssd1 vccd1 vccd1 _09413_ sky130_fd_sc_hd__inv_2
X_13749_ _03897_ _03899_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ _06425_ _06851_ _06853_ _06856_ _06858_ vssd1 vssd1 vccd1 vccd1 _06859_ sky130_fd_sc_hd__o311a_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15419_ _02991_ _08876_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__a21oi_1
X_18207_ _04900_ _08428_ _02994_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16399_ _06780_ _06781_ _06782_ vssd1 vssd1 vccd1 vccd1 _06784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18138_ _08609_ _08610_ _08607_ vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold103 _00023_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold114 net114 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18069_ _06394_ _06790_ _08601_ _04647_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold125 _00028_ vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 net87 vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 net107 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09911_ _06277_ _06288_ _06298_ vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_22_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _07700_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__clkbuf_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07036_ sky130_fd_sc_hd__buf_4
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11100_ _01167_ _01170_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__nand2_1
X_12080_ _02164_ _02166_ vssd1 vssd1 vccd1 vccd1 _02173_ sky130_fd_sc_hd__xnor2_2
X_11031_ _05671_ _04580_ _01122_ _01123_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__a31o_1
X_15770_ _06101_ _06102_ vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__xor2_1
X_12982_ _07810_ _03074_ _03024_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__o21ai_1
X_14721_ _04937_ _04936_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__and2b_2
XFILLER_0_99_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11933_ _01968_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__nand2_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ _06374_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__a21o_1
X_14652_ _00253_ _05975_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__nand2_4
X_11864_ _01953_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__xor2_2
XFILLER_0_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13603_ _03738_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nand2_1
X_10815_ _00906_ _00907_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__nor2_2
X_17371_ _07723_ _07725_ _07721_ _07018_ vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__o2bb2a_1
X_14583_ _04809_ _04811_ vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__xnor2_2
X_11795_ _01844_ _01870_ net199 _01869_ vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16322_ _02982_ _06500_ _06699_ _06466_ vssd1 vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13534_ _03661_ _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__xor2_1
X_10746_ _06019_ _08039_ _08049_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16253_ _06466_ vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__clkbuf_4
X_13465_ _03366_ _05311_ _05028_ _03345_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__a22oi_2
X_10677_ _04263_ _04253_ _04231_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15204_ _05485_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12416_ _02500_ _02508_ vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16184_ _06550_ vssd1 vssd1 vccd1 vccd1 _06551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13396_ _03333_ _03335_ _03512_ _03513_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__o211ai_4
X_15135_ _04950_ net117 vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__nand2_2
XFILLER_0_49_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12347_ _02437_ _02438_ _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15066_ _05335_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__or2_1
X_12278_ _07711_ _00247_ _02370_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14017_ _04028_ _04039_ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _00835_ _01321_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__and2b_1
X_18825_ _09125_ _09328_ vssd1 vssd1 vccd1 vccd1 _09329_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18756_ _09273_ _09274_ vssd1 vssd1 vccd1 vccd1 _09275_ sky130_fd_sc_hd__and2_1
X_15968_ _03920_ _05097_ vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__nor2_1
X_17707_ _08206_ _08207_ vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__nor2_1
X_14919_ _05176_ _05177_ vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__and2_1
X_18687_ _09222_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__clkbuf_1
X_15899_ _06211_ _06241_ vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17638_ _08023_ _08027_ vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17569_ _07944_ _08056_ vssd1 vssd1 vccd1 vccd1 _08057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09825_ _07591_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__clkbuf_8
X_09756_ _05551_ _05791_ _06841_ vssd1 vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__a21o_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _06084_ _06094_ _05257_ _06040_ vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a22o_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ _00690_ _00691_ _00507_ _00528_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__a211o_1
XFILLER_0_92_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11580_ _01106_ _01671_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__or3b_4
XFILLER_0_25_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10531_ _04373_ _05617_ _05246_ _04351_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _00752_ _00754_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ _00539_ _00540_ _00554_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12201_ _02287_ _02291_ _02292_ _02290_ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _00639_ _00642_ _00640_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10393_ _00482_ _00483_ _00484_ _00485_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12132_ _02223_ _02210_ _02221_ vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16940_ _02972_ _07371_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__nand2_1
X_12063_ _02135_ _02155_ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__nand2_1
X_11014_ _01106_ _00514_ _06776_ _00309_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__or4b_4
X_16871_ _07285_ _07295_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__xnor2_1
X_18610_ salida\[22\] _09159_ _09160_ salida\[54\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09165_ sky130_fd_sc_hd__a221o_1
X_15822_ _06157_ _06158_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__nor2_1
X_18541_ net13 net2 vssd1 vssd1 vccd1 vccd1 _09111_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15753_ _04823_ _06081_ _06082_ _06085_ vssd1 vssd1 vccd1 vccd1 _09370_ sky130_fd_sc_hd__a31o_1
X_12965_ _03024_ _03057_ vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14704_ _04814_ _04812_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__and2b_1
X_11916_ _02007_ _02008_ vssd1 vssd1 vccd1 vccd1 _02009_ sky130_fd_sc_hd__or2_1
X_15684_ _05955_ _06009_ vssd1 vssd1 vccd1 vccd1 _06011_ sky130_fd_sc_hd__and2_1
X_18472_ _03108_ _04853_ _08150_ vssd1 vssd1 vccd1 vccd1 _09038_ sky130_fd_sc_hd__and3_1
X_12896_ _04099_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__clkbuf_8
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _07896_ _07898_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__xnor2_1
X_14635_ _04865_ _04866_ _04737_ _04739_ vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__a211o_4
XFILLER_0_68_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11847_ _01917_ _01918_ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _04791_ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17354_ _07710_ _07716_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11778_ net199 _01869_ _01844_ _01870_ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13517_ _03644_ _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nor2_1
X_16305_ _06424_ _06430_ vssd1 vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__or2_1
X_10729_ _06149_ _06159_ _06170_ _05181_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__a22o_1
X_17285_ _06581_ _07621_ _07742_ _07746_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__a2bb2o_1
X_14497_ _04001_ _09248_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16236_ _06600_ _06604_ _06606_ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__and3_1
X_13448_ _03162_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _00217_ _00909_ vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__or2_1
X_13379_ _01356_ _00166_ _03326_ _03325_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__a31o_1
X_15118_ _05392_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16098_ _06426_ _06453_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__o21ai_1
X_15049_ _05317_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__xnor2_1
X_09610_ _05235_ _05257_ vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__nand2_1
X_18808_ _09315_ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__clkbuf_1
X_09541_ _04504_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__buf_4
X_18739_ _03117_ net61 _09251_ vssd1 vssd1 vccd1 vccd1 _09261_ sky130_fd_sc_hd__mux2_1
X_09472_ _03728_ _03750_ vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__nand2_4
XFILLER_0_148_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09808_ _07232_ _07254_ _07406_ _07102_ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__and4_1
X_09739_ _06646_ _06656_ vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12750_ _02669_ _02670_ _02632_ vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__o21a_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _01251_ _01793_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__nor2_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _02768_ _02772_ _02739_ _02763_ vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__o211a_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _00195_ _00702_ _05845_ _00443_ vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__and4_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _01722_ _01723_ _01724_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__nand3_1
XFILLER_0_139_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14351_ _03131_ _03178_ _03080_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ _01082_ vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _03226_ _03234_ _03233_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__a21o_1
X_10514_ _00604_ _00605_ _00606_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__nand3_1
X_17070_ net334 _07124_ _07126_ _07511_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__or4_1
X_14282_ _04480_ _04481_ vssd1 vssd1 vccd1 vccd1 _04483_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11494_ _05224_ _04056_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16021_ _06370_ _06371_ _04853_ vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__a21bo_1
X_13233_ _03333_ _03334_ _03314_ vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__o21a_1
X_10445_ _00396_ _00397_ _00415_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ _03240_ _03241_ _03261_ _03262_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__a22oi_2
X_10376_ _00299_ _00300_ vssd1 vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12115_ _08713_ _00131_ _02206_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__and4_1
X_17972_ _08449_ _08400_ _08495_ vssd1 vssd1 vccd1 vccd1 _08497_ sky130_fd_sc_hd__o21ai_1
X_13095_ _02505_ _01671_ vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__nor2_1
X_12046_ _02088_ _02138_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__and2_1
X_16923_ _02751_ _02836_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16854_ _03198_ _04414_ _07266_ _07278_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__a211o_1
X_15805_ _02976_ _04241_ _04415_ _03036_ vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__a31o_1
X_13997_ _04041_ vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16785_ _07107_ _07202_ vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__nor2_1
X_18524_ _03201_ _09092_ _09093_ vssd1 vssd1 vccd1 vccd1 _09094_ sky130_fd_sc_hd__and3_1
X_12948_ _01695_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__clkbuf_4
X_15736_ _06065_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18455_ _09018_ _09019_ vssd1 vssd1 vccd1 vccd1 _09020_ sky130_fd_sc_hd__or2b_1
X_12879_ _07058_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__buf_4
X_15667_ _02997_ _03154_ vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nand2_1
XANTENNA_170 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17406_ _07878_ _07879_ vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14618_ _04841_ _04843_ _04848_ vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nand3_1
X_15598_ _02994_ _02997_ _04125_ _03153_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__and4_1
X_18386_ _03068_ _06464_ _08924_ _08945_ vssd1 vssd1 vccd1 vccd1 _09405_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14549_ _01873_ _01112_ vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__nand2_1
X_17337_ _07801_ _07802_ _07803_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17268_ _07718_ _07728_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19007_ clknet_4_7_0_clk _09374_ vssd1 vssd1 vccd1 vccd1 salida\[60\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16219_ _06586_ _06587_ _06513_ vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17199_ _07652_ _07531_ _07653_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09524_ _04023_ _04110_ _04165_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _03454_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10230_ _08865_ _00322_ _00317_ _00320_ vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_14_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ _00253_ _00212_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10092_ _00183_ _00177_ _00146_ _00184_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13920_ _04074_ _04086_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__or2_1
X_13851_ _00170_ _04591_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ _00592_ _00881_ _01481_ _01479_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__a31o_1
X_13782_ _03574_ _00459_ _03932_ _03933_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__a22o_1
X_16570_ _06968_ vssd1 vssd1 vccd1 vccd1 _06969_ sky130_fd_sc_hd__clkbuf_4
X_10994_ _07036_ _07069_ _08746_ _06613_ vssd1 vssd1 vccd1 vccd1 _01087_ sky130_fd_sc_hd__nand4_1
XFILLER_0_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15521_ _02993_ _02996_ _00665_ _03071_ vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__and4_1
X_12733_ _02823_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__and2_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15452_ _05755_ _05756_ _05717_ _05718_ vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__o211ai_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18240_ _06368_ _07390_ _08700_ _08699_ vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__a31o_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _00845_ _00134_ _02720_ vssd1 vssd1 vccd1 vccd1 _02757_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _07504_ _03750_ _04012_ _00358_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11615_ _01166_ _01176_ _01177_ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__or3_4
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15383_ _05681_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18171_ _08629_ _08698_ _08711_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12595_ _07700_ _00194_ _02646_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ _04426_ _04385_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17122_ _00787_ _06331_ _06365_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ _01619_ _01620_ _01605_ _01606_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17053_ _07388_ _07492_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__and2_1
X_14265_ _04287_ _04291_ _04292_ _04294_ _04286_ vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__a32o_1
X_11477_ _06591_ _03476_ _00210_ _00806_ vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__a22o_1
X_16004_ _06338_ _06350_ _06353_ _06339_ vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ _01503_ _00511_ _00684_ _00686_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10428_ _00134_ _00359_ _00520_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14196_ _04214_ _04216_ vssd1 vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _07744_ _03243_ _03244_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _04427_ _06613_ _08049_ _04504_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _03026_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__and2_1
X_17955_ _08475_ _08476_ _08352_ _08471_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__o211ai_1
X_12029_ _02108_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__or2_1
X_16906_ _07333_ _07334_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__xor2_1
X_17886_ _08292_ _08348_ _08402_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16837_ _07168_ _07170_ _07165_ vssd1 vssd1 vccd1 vccd1 _07260_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16768_ _07183_ _07184_ _03920_ vssd1 vssd1 vccd1 vccd1 _07185_ sky130_fd_sc_hd__mux2_1
X_18507_ _03011_ _06512_ _03155_ vssd1 vssd1 vccd1 vccd1 _09075_ sky130_fd_sc_hd__a21boi_1
X_15719_ _06046_ _06047_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__xnor2_1
X_16699_ _07108_ vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__clkbuf_4
X_18438_ _09000_ _04995_ _06277_ vssd1 vssd1 vccd1 vccd1 _09001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18369_ _08925_ _08926_ vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09507_ _03914_ vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09438_ ApproximateM_inst.lob_16.lob1.genblk1\[10\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03388_ sky130_fd_sc_hd__buf_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11400_ _01490_ _01491_ _01415_ _01454_ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _02423_ vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__inv_2
XANTENNA_70 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _07810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11331_ cla_inst.in2\[21\] _00223_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__nand2_1
XANTENNA_92 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _04225_ _04226_ _04227_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _01353_ _01354_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__xor2_4
XFILLER_0_30_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13001_ _00214_ vssd1 vssd1 vccd1 vccd1 _03094_ sky130_fd_sc_hd__clkbuf_4
X_10213_ _08539_ _08594_ vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__or2b_1
X_11193_ _01284_ _01285_ vssd1 vssd1 vccd1 vccd1 _01286_ sky130_fd_sc_hd__nand2_1
X_10144_ _00109_ _09349_ _00146_ _00197_ vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17740_ _03119_ _05621_ _06705_ _08243_ vssd1 vssd1 vccd1 vccd1 _08244_ sky130_fd_sc_hd__a2bb2o_1
X_14952_ _05211_ _05212_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__nor2_1
X_10075_ _00164_ _00167_ vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__nand2_2
X_13903_ _03900_ _03901_ _03738_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__o21a_1
X_17671_ _08052_ _08053_ vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__nand2_1
X_14883_ _05136_ _05138_ vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__nor2_1
X_16622_ _07023_ _07024_ _06040_ vssd1 vssd1 vccd1 vccd1 _07026_ sky130_fd_sc_hd__o21a_2
X_13834_ _03986_ _03989_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__or3_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16553_ _06802_ _06806_ _03535_ vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a21o_2
X_13765_ _03164_ _03066_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nor2_2
X_10977_ _01044_ _01047_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ _03322_ _03321_ _08224_ _08158_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__nand4_4
XFILLER_0_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ _02785_ _02806_ _02808_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13696_ _00169_ _04700_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__nand2_1
X_16484_ _06563_ _06875_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18223_ _03198_ _06083_ _07184_ _08141_ vssd1 vssd1 vccd1 vccd1 _08770_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_127_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ _05659_ _05658_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__or2b_1
X_12647_ _02701_ _02702_ _02703_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15366_ _05653_ _05585_ _05664_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__a21oi_1
X_18154_ _03052_ _06463_ _08672_ _08694_ vssd1 vssd1 vccd1 vccd1 _09401_ sky130_fd_sc_hd__a22oi_2
X_12578_ _02669_ _02670_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17105_ _07549_ _07551_ vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__xnor2_1
X_14317_ _04519_ _04520_ vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__xnor2_1
X_11529_ _01185_ _01183_ _01184_ vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__nand3_1
X_15297_ _05588_ _05589_ vssd1 vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__nand2_1
X_18085_ _07649_ _07489_ _07596_ _07664_ vssd1 vssd1 vccd1 vccd1 _08619_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _04442_ _04443_ _04444_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__and3_2
X_17036_ _03920_ _07474_ _07476_ _06645_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14179_ _04158_ _04368_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__nand2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ clknet_4_6_0_clk _09383_ vssd1 vssd1 vccd1 vccd1 salida\[40\] sky130_fd_sc_hd__dfxtp_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _07130_ _07706_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17869_ _07302_ _07741_ vssd1 vssd1 vccd1 vccd1 _08384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09987_ _09271_ _09279_ vssd1 vssd1 vccd1 vccd1 _09287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10900_ _00992_ _05638_ _04569_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__and3_1
Xwb_buttons_leds_155 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_155/HI led_enb[4] sky130_fd_sc_hd__conb_1
X_11880_ _01960_ _01968_ net193 _01972_ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _00922_ _00923_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__xnor2_1
X_13550_ _03680_ _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__xor2_2
XFILLER_0_13_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10762_ _08278_ _08289_ _08300_ _06938_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_149_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12501_ _02550_ _02555_ _02554_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13481_ _03603_ _03604_ _03605_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__and3_2
X_10693_ _04635_ _03739_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__nand2_4
XFILLER_0_152_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15220_ _05387_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ _02456_ _02522_ _02515_ net122 vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _05223_ _05329_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _02450_ _02454_ _02455_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__or3_4
X_14102_ _04112_ _04113_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2_2
X_11314_ _01304_ _01306_ _01405_ net139 vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15082_ _09352_ _00309_ _05352_ _05353_ vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12294_ _02263_ _02386_ vssd1 vssd1 vccd1 vccd1 _02387_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14033_ _04192_ _04193_ _04207_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__and3_1
X_18910_ clknet_4_8_0_clk _00064_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[28\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_31_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ _01120_ _01144_ _01118_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18841_ clknet_4_0_0_clk net260 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__dfxtp_1
X_11176_ _01267_ _01268_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__nor2_1
X_10127_ _00216_ _00219_ _00170_ _00206_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__and4bb_1
X_18772_ _09273_ _09286_ vssd1 vssd1 vccd1 vccd1 _09288_ sky130_fd_sc_hd__and2_1
X_15984_ _06993_ _00108_ vssd1 vssd1 vccd1 vccd1 _06332_ sky130_fd_sc_hd__or2_1
X_17723_ _02849_ _02846_ vssd1 vssd1 vccd1 vccd1 _08226_ sky130_fd_sc_hd__or2b_1
X_10058_ cla_inst.in2\[27\] vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__clkbuf_4
X_14935_ _05194_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17654_ _07825_ vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__clkbuf_4
X_14866_ _04986_ _04990_ _05118_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ _06345_ _06545_ _07007_ _03169_ vssd1 vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a22o_1
X_13817_ _03972_ _03973_ vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__xnor2_2
X_17585_ _08067_ _07947_ _08073_ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__nor3_1
X_14797_ _05043_ _05044_ vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__or2b_1
X_16536_ _06904_ _06907_ _06932_ _06463_ _03086_ vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__a32o_2
X_13748_ _03368_ _03693_ _03692_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16467_ _06349_ _06338_ _06348_ _06598_ _06857_ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__a311o_1
X_13679_ _03817_ _03820_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__or3_2
XFILLER_0_73_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18206_ _02994_ _06511_ _06776_ vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15418_ _09350_ _07015_ vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16398_ _06780_ _06781_ _06782_ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__nand3_1
XFILLER_0_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _03052_ _08428_ _02997_ vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__or3b_1
X_15349_ _05644_ _05645_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold104 net102 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _00013_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18068_ _02998_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _08601_ sky130_fd_sc_hd__a21o_1
Xhold126 net90 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _00017_ vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 net105 vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09910_ _08496_ _08507_ _08518_ vssd1 vssd1 vccd1 vccd1 _08529_ sky130_fd_sc_hd__and3_2
X_17019_ _02968_ _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09841_ _07711_ _07744_ _07766_ vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__nand3_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _07015_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__clkbuf_8
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11030_ _00992_ _08039_ _04449_ _04471_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__and4_1
X_12981_ _03025_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__and2_1
X_14720_ _04953_ _04954_ _04956_ _03125_ _04960_ vssd1 vssd1 vccd1 vccd1 _09357_ sky130_fd_sc_hd__a221o_1
X_11932_ _01965_ _01966_ _01967_ _01961_ vssd1 vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__o31ai_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14651_ _04764_ _04765_ vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__nand2_1
X_11863_ _01954_ _01955_ vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13602_ _03736_ _03737_ vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nand2_1
X_10814_ _00761_ _00905_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__and2_1
X_17370_ _07823_ _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__xor2_1
X_14582_ _04678_ _04681_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__nor2_1
X_11794_ _01881_ _01884_ _01885_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__a211o_2
XFILLER_0_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16321_ _03047_ _06489_ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__or2_1
X_13533_ _02972_ _03456_ _03663_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__and3_1
X_10745_ _08039_ net230 net222 _06019_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13464_ _03454_ _05377_ vssd1 vssd1 vccd1 vccd1 _03588_ sky130_fd_sc_hd__nand2_8
X_16252_ _03048_ _06623_ vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _04263_ _04231_ _04253_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__nand3_1
X_15203_ _05370_ _05487_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__nor2_1
X_12415_ _02501_ _02507_ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__or2b_1
X_13395_ _03510_ _03511_ _03471_ _03472_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__a211o_1
X_16183_ _06459_ _03292_ _03217_ vssd1 vssd1 vccd1 vccd1 _06550_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15134_ _05198_ _05201_ _05302_ _05412_ vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__o31a_1
X_12346_ _02371_ _02436_ vssd1 vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15065_ _00362_ _00461_ _05336_ _05332_ vssd1 vssd1 vccd1 vccd1 _05337_ sky130_fd_sc_hd__o2bb2a_1
X_12277_ _00120_ _00398_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__and2_2
X_14016_ _03823_ _04038_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11228_ _06971_ _05704_ _00833_ _00834_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ _06200_ net59 _09250_ vssd1 vssd1 vccd1 vccd1 _09328_ sky130_fd_sc_hd__mux2_1
X_11159_ _01231_ _01233_ vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18755_ _02476_ net66 _09251_ vssd1 vssd1 vccd1 vccd1 _09274_ sky130_fd_sc_hd__mux2_1
X_15967_ _06314_ _03930_ vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__and2_4
X_17706_ _08203_ _08205_ vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__nor2_1
X_14918_ _00591_ _03142_ _05175_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__a21o_1
X_18686_ _09209_ _09221_ vssd1 vssd1 vccd1 vccd1 _09222_ sky130_fd_sc_hd__and2_1
X_15898_ _06238_ _06240_ vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17637_ _08129_ _08131_ vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__and2_1
X_14849_ _03596_ _07755_ cla_inst.in1\[27\] _03629_ vssd1 vssd1 vccd1 vccd1 _05101_
+ sky130_fd_sc_hd__a22o_1
X_17568_ _06969_ _07596_ vssd1 vssd1 vccd1 vccd1 _08056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16519_ _06616_ _06621_ _03099_ vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17499_ _07207_ net146 _07664_ _06947_ vssd1 vssd1 vccd1 vccd1 _07981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09824_ _07581_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__clkbuf_8
X_09755_ _05540_ _05442_ vssd1 vssd1 vccd1 vccd1 _06841_ sky130_fd_sc_hd__and2b_1
X_09686_ _06062_ vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__buf_4
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10530_ _04984_ _00443_ _00441_ _00440_ _04132_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10461_ _00542_ _00553_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12200_ _02287_ _02290_ _02291_ _02292_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__nor4_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13180_ _00669_ _00670_ vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__nand2_1
X_10392_ _00316_ _00324_ vssd1 vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12131_ _02210_ _02221_ _02223_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12062_ _02049_ _02107_ _02134_ vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__or3_1
X_11013_ _01105_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__buf_4
X_16870_ _07287_ _07294_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__xnor2_2
X_15821_ _03016_ _03154_ _06154_ _06156_ vssd1 vssd1 vccd1 vccd1 _06158_ sky130_fd_sc_hd__a22oi_1
X_18540_ net28 _09109_ net27 vssd1 vssd1 vccd1 vccd1 _09110_ sky130_fd_sc_hd__or3b_2
X_15752_ _04264_ _05623_ _06083_ _03124_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__a22o_1
X_12964_ _03027_ _03056_ _01114_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__a21o_1
X_14703_ _04811_ _04809_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__and2b_1
X_11915_ _01928_ _01931_ vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__xnor2_1
X_18471_ _09007_ vssd1 vssd1 vccd1 vccd1 _09036_ sky130_fd_sc_hd__inv_2
X_15683_ _05955_ _06009_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nor2_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _01520_ vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__clkbuf_8
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _06750_ _07780_ _07778_ _07776_ vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__a31oi_2
X_14634_ _04737_ _04739_ _04865_ _04866_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__o211ai_4
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _01936_ _01937_ net341 _01932_ vssd1 vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__a211oi_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _07705_ _07717_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__or2b_1
X_14565_ _04778_ _04779_ _04790_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__or3_1
X_11777_ _01843_ _01842_ _01841_ _01828_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__o211a_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16304_ _02981_ _06592_ _06550_ vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__a21o_1
X_13516_ _03642_ _03643_ _03422_ _03424_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__o211a_1
X_10728_ _00797_ _00819_ _00820_ vssd1 vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__nor3_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17284_ _06581_ _07621_ _07742_ _07746_ vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__or4bb_2
X_14496_ _04714_ _04715_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16235_ _02806_ _02968_ _06605_ vssd1 vssd1 vccd1 vccd1 _06606_ sky130_fd_sc_hd__or3b_1
XFILLER_0_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10659_ _00585_ _00599_ _00750_ _00751_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__o211a_2
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ _03567_ _03568_ _03098_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13378_ _03319_ _03329_ _03493_ vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16166_ _00211_ _06529_ _06530_ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__or3_2
XFILLER_0_140_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15117_ _05243_ _05287_ _05393_ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__o21ba_1
X_12329_ _02419_ _02421_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _03038_ _06454_ _06455_ _03120_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__o22a_1
X_15048_ _02987_ _00513_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__nand2_1
X_18807_ _09298_ _09314_ vssd1 vssd1 vccd1 vccd1 _09315_ sky130_fd_sc_hd__and2_1
X_16999_ _07316_ _07320_ _07315_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__o21ba_1
X_09540_ _04493_ vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__buf_6
X_18738_ _09260_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__buf_1
X_09471_ _03739_ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__buf_6
X_18669_ net36 _03101_ _09193_ vssd1 vssd1 vccd1 vccd1 _09210_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_506 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09807_ cla_inst.in1\[26\] vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__clkbuf_4
X_09738_ _05235_ _05257_ _05421_ _05344_ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__a31o_1
X_09669_ _05410_ _05366_ _05497_ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__and3_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _01226_ _01250_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__nor2_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _02739_ _02763_ _02768_ _02772_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _01685_ _01686_ _01684_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__a21bo_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _01646_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14350_ _03125_ _04414_ _04419_ _03199_ _04556_ vssd1 vssd1 vccd1 vccd1 _09384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10513_ _03465_ _04460_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__and2_1
X_13301_ _03406_ _03407_ _03224_ _03375_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a211o_2
XFILLER_0_64_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14281_ _04477_ _04479_ _04474_ vssd1 vssd1 vccd1 vccd1 _04481_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11493_ _01581_ _01584_ _01583_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13232_ _03314_ _03333_ _03334_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nor3_4
X_16020_ _02200_ _03311_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__or2_1
X_10444_ net186 _00375_ _00535_ _00536_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__o211a_2
XFILLER_0_134_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13163_ _03258_ _03259_ _00651_ _00653_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__o211ai_2
X_10375_ _00292_ _00298_ vssd1 vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ _05301_ _09212_ _09188_ _05279_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13094_ _02125_ _03186_ _03022_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__o21a_1
X_17971_ _08484_ _08494_ vssd1 vssd1 vccd1 vccd1 _08495_ sky130_fd_sc_hd__xnor2_1
X_12045_ _02083_ _02087_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__nand2_1
X_16922_ _02751_ _02836_ vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__or2_1
X_16853_ _06462_ _07271_ _07273_ _07277_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15804_ _06137_ _06139_ vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16784_ _07200_ _07201_ vssd1 vssd1 vccd1 vccd1 _07202_ sky130_fd_sc_hd__nand2_1
X_13996_ _04166_ _04167_ _04168_ vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__a21oi_1
X_18523_ _02949_ _09061_ _02956_ vssd1 vssd1 vccd1 vccd1 _09093_ sky130_fd_sc_hd__o21ai_1
X_15735_ _06023_ _06064_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__and2_1
X_12947_ _03022_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__clkbuf_4
X_18454_ _03073_ _08428_ _03013_ vssd1 vssd1 vccd1 vccd1 _09019_ sky130_fd_sc_hd__or3b_1
X_15666_ _05989_ _05990_ vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__nand2_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _00759_ _02964_ _02970_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__o21ai_2
XANTENNA_160 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17405_ _07854_ _07877_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__and2_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14617_ _04846_ _04847_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__xnor2_1
X_18385_ _07256_ _08929_ _08931_ _08944_ vssd1 vssd1 vccd1 vccd1 _08945_ sky130_fd_sc_hd__a31o_1
X_11829_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel _03607_ vssd1
+ vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__and2_1
X_15597_ _02997_ _04125_ _03153_ _02994_ vssd1 vssd1 vccd1 vccd1 _05916_ sky130_fd_sc_hd__a22oi_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17336_ _07801_ _07802_ _07803_ vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14548_ _04771_ _04772_ vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__nor2_1
X_17267_ _07719_ _07727_ vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14479_ _03125_ _04559_ _04563_ _03199_ _04697_ vssd1 vssd1 vccd1 vccd1 _09385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19006_ clknet_4_5_0_clk _09373_ vssd1 vssd1 vccd1 vccd1 salida\[59\] sky130_fd_sc_hd__dfxtp_1
X_16218_ _01106_ _07646_ _06585_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__or3_1
XFILLER_0_140_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17198_ _06581_ _07516_ _07512_ _07513_ vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__o31a_1
X_16149_ _06511_ vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09523_ _03968_ _03979_ _04307_ vssd1 vssd1 vccd1 vccd1 _04318_ sky130_fd_sc_hd__nand3_4
XFILLER_0_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09454_ _03443_ _03542_ _03487_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10160_ _00169_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__buf_4
X_10091_ cla_inst.in2\[24\] vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__clkbuf_4
X_13850_ _04008_ _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12801_ _02892_ _02888_ _02889_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__o22ai_4
X_13781_ _03574_ _00459_ _03932_ _03933_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nand4_2
X_10993_ _06471_ _00993_ _00991_ _00995_ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15520_ _02996_ _03153_ _03071_ _02993_ vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__a22o_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12732_ _02818_ _02824_ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _05717_ _05718_ _05755_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__a211o_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _02721_ _02755_ vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14402_ _00358_ _07504_ _03750_ _04012_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__and4_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11614_ _01642_ _01704_ _01705_ _01706_ vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__nor4_2
X_18170_ _08709_ _08710_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__nand2_1
X_15382_ _03015_ _01112_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__nand2_1
X_12594_ _02647_ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__nor2_1
X_17121_ _07565_ _07566_ _07567_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14333_ _04489_ _04490_ _04535_ _04536_ vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11545_ _01636_ _01637_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17052_ _07388_ _07492_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__nor2_1
X_14264_ _04305_ _04306_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__or2b_1
X_11476_ _01565_ _01567_ _01566_ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a21o_1
X_16003_ _06341_ _06345_ _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__and3_1
X_13215_ _00724_ _00731_ _03316_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__a21o_1
X_10427_ _07504_ _00131_ _09219_ _00358_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__a22o_1
X_14195_ _04385_ _04386_ _04169_ net120 vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13146_ _06051_ _00498_ _07384_ _06029_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a22o_1
X_10358_ _04351_ _00294_ _05246_ _05322_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__nand4_2
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _00878_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__clkbuf_4
X_17954_ _08352_ _08471_ _08475_ _08476_ vssd1 vssd1 vccd1 vccd1 _08477_ sky130_fd_sc_hd__a211o_1
X_10289_ _00241_ _00235_ vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__and2b_1
X_12028_ _02111_ _02119_ _02120_ vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a21oi_1
X_16905_ _07220_ _07222_ _07219_ vssd1 vssd1 vccd1 vccd1 _07334_ sky130_fd_sc_hd__o21ai_2
X_17885_ _08400_ _08401_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__nor2_1
X_16836_ _07257_ _07258_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16767_ _02979_ _06494_ vssd1 vssd1 vccd1 vccd1 _07184_ sky130_fd_sc_hd__or2_1
X_13979_ _03005_ _00213_ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__nand2_1
X_18506_ _09044_ _09047_ _09073_ _06649_ vssd1 vssd1 vccd1 vccd1 _09074_ sky130_fd_sc_hd__o31a_1
X_15718_ _05972_ _05982_ _05980_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__a21oi_1
X_16698_ _02533_ _07104_ _07105_ vssd1 vssd1 vccd1 vccd1 _07108_ sky130_fd_sc_hd__and3_2
X_18437_ _06374_ _03311_ vssd1 vssd1 vccd1 vccd1 _09000_ sky130_fd_sc_hd__nand2_1
X_15649_ _01359_ _03071_ _05900_ _05898_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18368_ _03068_ _08428_ _02992_ vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17319_ _07783_ _07784_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ _07314_ _08260_ _08777_ _04023_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__or4b_1
XFILLER_0_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ _04121_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_67_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ net172 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__buf_6
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_60 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _05845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ cla_inst.in2\[21\] _00193_ _01349_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__and3_1
XANTENNA_82 _07810_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_93 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ _00163_ _00223_ vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__nand2_2
X_10212_ _08529_ _08659_ _00303_ _00304_ vssd1 vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__o211a_1
X_13000_ _03040_ _03092_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11192_ _01283_ _01280_ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__or2b_1
X_10143_ _00106_ _00194_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14951_ _02984_ _01520_ _09256_ _00498_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__and4_2
X_10074_ _00166_ vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__buf_4
X_13902_ _04065_ _04066_ vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__nand2_1
X_17670_ _08165_ _08166_ vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__nor2_1
X_14882_ _05100_ _05013_ _05135_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nor3_1
X_16621_ _04132_ _03184_ _03313_ net150 vssd1 vssd1 vccd1 vccd1 _07024_ sky130_fd_sc_hd__a211oi_2
X_13833_ _07537_ _00247_ _03988_ _03991_ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16552_ _06945_ _06948_ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13764_ _03054_ _03058_ _03070_ _03075_ _03050_ _03061_ vssd1 vssd1 vccd1 vccd1 _03917_
+ sky130_fd_sc_hd__mux4_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _01040_ _01043_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _03321_ _07384_ _08158_ _03322_ vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12715_ _02783_ _02784_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__a21oi_1
X_16483_ _06874_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13695_ _03839_ _03840_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18222_ _06776_ _08766_ _08767_ _06721_ vssd1 vssd1 vccd1 vccd1 _08769_ sky130_fd_sc_hd__o211a_1
X_15434_ _05737_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12646_ _02733_ _02737_ _02738_ vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__nand3_2
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18153_ _02969_ _08674_ _08693_ vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15365_ _05662_ _05663_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12577_ _02592_ _02631_ vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17104_ _07432_ _07433_ _07550_ vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__o21ai_1
X_14316_ _00107_ _04591_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _01605_ _01606_ _01619_ _01620_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__a211oi_4
X_18084_ _08541_ _08542_ _08543_ _08537_ vssd1 vssd1 vccd1 vccd1 _08618_ sky130_fd_sc_hd__or4b_1
X_15296_ _05575_ _05576_ _05587_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__nand3_1
XFILLER_0_150_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17035_ _02973_ _07475_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__nor2_1
X_14247_ _04275_ _04281_ _04273_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__a21o_1
X_11459_ _03717_ _00177_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _04158_ _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__or2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13129_ _03221_ _03222_ _03223_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__a21oi_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ clknet_4_1_0_clk _09382_ vssd1 vssd1 vccd1 vccd1 salida\[39\] sky130_fd_sc_hd__dfxtp_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _08456_ _08457_ vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17868_ _07303_ _07621_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16819_ _07231_ _07239_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__xor2_1
X_17799_ _07038_ _07859_ _08306_ vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09986_ _07700_ _07733_ _07766_ vssd1 vssd1 vccd1 vccd1 _09279_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwb_buttons_leds_156 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_156/HI led_enb[5] sky130_fd_sc_hd__conb_1
X_10830_ _03717_ _03476_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10761_ _00824_ _00852_ _00853_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__and3_2
XFILLER_0_82_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _02576_ _02577_ vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__xnor2_1
X_13480_ _03383_ _03389_ _03382_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__a21bo_1
X_10692_ _00783_ _00784_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__or2_1
X_12431_ _02439_ _02518_ vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15150_ _05345_ _05346_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ net128 _02449_ _02416_ _02448_ vssd1 vssd1 vccd1 vccd1 _02455_ sky130_fd_sc_hd__o211a_1
X_14101_ _04267_ _04268_ _04282_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__nor3_1
XFILLER_0_105_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11313_ _01396_ _01404_ _01397_ _01398_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor4_1
X_15081_ _05352_ _05353_ _00106_ _00309_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__and4bb_1
X_12293_ _02378_ _02380_ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14032_ _04208_ vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__inv_2
X_11244_ _01079_ _01147_ _01335_ _01336_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_31_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11175_ _01141_ _01266_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__and2_1
X_18840_ clknet_4_1_0_clk net312 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__dfxtp_1
X_10126_ _00175_ _00218_ _00178_ _00173_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__a22oi_1
X_18771_ _02200_ net40 _09276_ vssd1 vssd1 vccd1 vccd1 _09286_ sky130_fd_sc_hd__mux2_1
X_15983_ _02347_ _00558_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__or2_1
X_17722_ _06516_ _08222_ _08223_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__and3_1
X_10057_ _00148_ _00149_ _00131_ _00127_ vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__nand4_2
X_14934_ _05069_ _05071_ vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17653_ _08065_ _08078_ vssd1 vssd1 vccd1 vccd1 _08149_ sky130_fd_sc_hd__nor2_1
X_14865_ _04986_ _04990_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16604_ _02728_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _07007_ sky130_fd_sc_hd__a21o_1
X_13816_ _05224_ _09256_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17584_ _08067_ _07947_ _08073_ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__o21a_1
X_14796_ _04887_ _04888_ _04889_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__o21ba_1
X_16535_ _06836_ _06911_ _06912_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__o31a_1
X_13747_ _03687_ _03688_ _03691_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__and3_1
X_10959_ _00941_ _00954_ _00953_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16466_ _06349_ _06348_ _06338_ vssd1 vssd1 vccd1 vccd1 _06857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13678_ _07526_ _00165_ _03819_ _03821_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18205_ _08748_ _08749_ vssd1 vssd1 vccd1 vccd1 _08750_ sky130_fd_sc_hd__and2b_1
X_15417_ _05449_ _01112_ _05678_ _05680_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__a31o_1
X_12629_ _02686_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__and2_1
X_16397_ _06674_ _06675_ _06672_ vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_115_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18136_ _02997_ _06512_ _03052_ vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__a21boi_1
X_15348_ _05563_ _05630_ _05643_ vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18067_ _04647_ _06445_ vssd1 vssd1 vccd1 vccd1 _08600_ sky130_fd_sc_hd__or2_1
Xhold105 _00031_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15279_ _05567_ _05569_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold116 net95 vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _00020_ vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 net94 vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _00006_ vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17018_ _07455_ _07456_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ ApproximateM_inst.lob_16.lob2.mux.sel _07755_ vssd1 vssd1 vccd1 vccd1 _07766_
+ sky130_fd_sc_hd__and2_4
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _07004_ vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__buf_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ clknet_4_5_0_clk _09400_ vssd1 vssd1 vccd1 vccd1 salida\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09969_ _09037_ _09048_ _09145_ vssd1 vssd1 vccd1 vccd1 _09152_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ _03072_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__buf_4
X_11931_ _02023_ vssd1 vssd1 vccd1 vccd1 _02024_ sky130_fd_sc_hd__inv_2
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _04603_ _04752_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__and2b_1
X_11862_ _01847_ _01846_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ _03736_ _03737_ vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__or2_1
X_10813_ _00761_ _00905_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__nor2_1
X_14581_ _04807_ _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__xor2_2
XFILLER_0_83_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11793_ _01601_ _01602_ _01603_ _01564_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ _03061_ _06696_ _06697_ vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__a21bo_1
X_13532_ _03453_ _03457_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__or2b_1
X_10744_ _07352_ _06722_ _07951_ _07995_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16251_ _03026_ _03041_ _01696_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__a21o_1
X_13463_ _03393_ _03394_ _03405_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10675_ _00766_ _00767_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__xor2_2
XFILLER_0_152_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15202_ _01505_ _00322_ _05371_ vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__and3_1
XFILLER_0_153_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ _02503_ _02504_ _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__and3_1
X_16182_ _03200_ _06547_ _06477_ vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__o21a_1
X_13394_ _03471_ _03472_ _03510_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15133_ _05196_ _05299_ _05300_ vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__o21ba_1
X_12345_ _00846_ _00248_ _02370_ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ _05334_ vssd1 vssd1 vccd1 vccd1 _05336_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12276_ _02353_ _02367_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14015_ _04189_ _04190_ vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__xor2_4
X_11227_ _05050_ _01009_ _01008_ _01011_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__o2bb2a_1
X_18823_ _09327_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__buf_1
X_11158_ _01226_ _01250_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__and2_1
X_10109_ _00188_ _00201_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__and2b_1
X_11089_ _08713_ _00715_ _01054_ _01055_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__a22o_2
X_18754_ _09125_ vssd1 vssd1 vccd1 vccd1 _09273_ sky130_fd_sc_hd__buf_2
X_15966_ _06299_ _06301_ _06312_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17705_ _08203_ _08205_ vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__and2_1
X_14917_ _00591_ _03142_ _05175_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__nand3_1
X_18685_ net43 _03111_ _09193_ vssd1 vssd1 vccd1 vccd1 _09221_ sky130_fd_sc_hd__mux2_1
X_15897_ _06194_ _06195_ _06197_ _06239_ vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__a31oi_2
X_14848_ _04862_ _04969_ _04997_ _04998_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__o211a_1
X_17636_ _08130_ vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17567_ _06961_ _07487_ _07593_ _07018_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__o22a_1
XFILLER_0_147_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14779_ _05019_ _05023_ _05024_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16518_ _02981_ _06611_ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17498_ _07302_ _07115_ _07218_ _07313_ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16449_ _03535_ _06673_ _01264_ vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18119_ _08488_ _08556_ _08559_ vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09823_ ApproximateM_inst.lob_16.lob1.mux.sel vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__clkbuf_4
X_09754_ _06558_ _06569_ _06808_ vssd1 vssd1 vccd1 vccd1 _06830_ sky130_fd_sc_hd__nand3_1
X_09685_ _05649_ vssd1 vssd1 vccd1 vccd1 _06084_ sky130_fd_sc_hd__buf_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10460_ _00543_ _00552_ vssd1 vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10391_ _00314_ _00315_ vssd1 vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12130_ _02187_ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12061_ _02148_ _02152_ _02070_ _02153_ vssd1 vssd1 vccd1 vccd1 _02154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11012_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _01105_ sky130_fd_sc_hd__inv_2
X_15820_ _03016_ _03154_ _06154_ _06156_ vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__and4_1
X_15751_ _04256_ _04261_ _03537_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__mux2_1
X_12963_ _03055_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ _04939_ _04940_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or2_4
X_11914_ _02001_ _02004_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__o21ai_1
X_18470_ _03073_ _06464_ _09017_ _09035_ vssd1 vssd1 vccd1 vccd1 _09407_ sky130_fd_sc_hd__o2bb2a_1
X_15682_ _06006_ _06007_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__or2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _02986_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__buf_4
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _07893_ _07895_ vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__xor2_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _04862_ _04863_ _04730_ _04833_ vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__o211ai_4
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ net341 _01932_ _01936_ _01937_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__o211a_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _07783_ _07784_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14564_ _04778_ _04779_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ _01861_ _01865_ _01867_ _01868_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__or4_4
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _06461_ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13515_ _03422_ _03424_ _03642_ _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__a211oi_4
X_10727_ _00795_ _00796_ _00779_ _00794_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__o211a_1
X_17283_ _07038_ _07665_ _07745_ _06527_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__a22o_1
X_14495_ _03859_ _03793_ cla_inst.in1\[28\] _07374_ vssd1 vssd1 vccd1 vccd1 _04715_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16234_ _03161_ _03029_ _02805_ vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13446_ _03145_ _03151_ _03089_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__mux2_1
X_10658_ _00747_ _00748_ _00749_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16165_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel net208 ApproximateM_inst.lob_16.lob1.genblk1\[10\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _06530_ sky130_fd_sc_hd__or4_4
X_13377_ _03320_ _03328_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ _00680_ _00681_ _07537_ _00194_ vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__and4bb_1
X_15116_ _05240_ _05242_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__and2b_1
X_12328_ _02419_ _02420_ _00832_ _03618_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__and4bb_1
X_16096_ _05419_ _05422_ _02974_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15047_ _05315_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__nor2_1
X_12259_ _02228_ _02350_ _02351_ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__and3_1
X_18806_ _01359_ net52 _09301_ vssd1 vssd1 vccd1 vccd1 _09314_ sky130_fd_sc_hd__mux2_1
X_16998_ _07324_ _07326_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__nor2_1
X_18737_ _09245_ _09259_ vssd1 vssd1 vccd1 vccd1 _09260_ sky130_fd_sc_hd__and2_1
X_15949_ _03121_ _06295_ vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__nand2_1
X_09470_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03739_ sky130_fd_sc_hd__buf_6
X_18668_ _09125_ vssd1 vssd1 vccd1 vccd1 _09209_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17619_ _07999_ _08007_ _07997_ vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__a21o_1
X_18599_ salida\[19\] _09141_ _09142_ salida\[51\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09156_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09806_ _07363_ _07384_ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__nand2_1
X_09737_ _06580_ _06635_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__xnor2_1
X_09668_ _05366_ _05497_ _04580_ _05410_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__a22o_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09599_ _04941_ _04952_ _04962_ vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__a21o_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _01215_ _01214_ _01209_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__a21o_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11561_ _01652_ _01653_ vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_835 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13300_ _03224_ net135 _03406_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _03651_ _03662_ _04580_ _04482_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__nand4_2
XFILLER_0_52_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _04474_ _04477_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__or3_2
X_11492_ _01581_ _01583_ _01584_ vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nand3_4
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13231_ _03315_ _00735_ _03332_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10443_ _00532_ _00533_ _00534_ _00491_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__a22o_1
X_13162_ _00651_ _00653_ _03258_ _03259_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__a211o_1
X_10374_ _00291_ _00431_ _00465_ _00466_ vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ _00127_ _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__nand2_1
X_13093_ _02505_ _01862_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__nor2_1
X_17970_ _08391_ _08493_ vssd1 vssd1 vccd1 vccd1 _08494_ sky130_fd_sc_hd__xor2_1
X_12044_ _02073_ _02076_ _02075_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__o21ai_1
X_16921_ _07349_ _07350_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor2_2
X_16852_ _06357_ _07274_ _07275_ _00167_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__a2bb2o_1
X_15803_ _06137_ _06139_ vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__or2_1
X_16783_ _06937_ _07143_ _07198_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__o21ai_1
X_13995_ _04166_ _04167_ _04168_ vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__and3_4
XFILLER_0_99_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15734_ _06023_ _06064_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__nor2_1
X_18522_ _02949_ _02956_ _09061_ vssd1 vssd1 vccd1 vccd1 _09092_ sky130_fd_sc_hd__or3_1
XFILLER_0_99_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ _03038_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__clkbuf_4
X_15665_ _05970_ _05971_ _05988_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__or3_1
X_18453_ _03013_ _06512_ _03073_ vssd1 vssd1 vccd1 vccd1 _09018_ sky130_fd_sc_hd__a21boi_1
X_12877_ _00759_ _02964_ _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__a21oi_1
XANTENNA_150 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _07854_ _07877_ vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__nor2_1
X_14616_ _04001_ _00502_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__nand2_1
XANTENNA_172 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18384_ _04238_ _08934_ _08943_ vssd1 vssd1 vccd1 vccd1 _08944_ sky130_fd_sc_hd__o21ai_1
X_11828_ _01831_ _01830_ _01829_ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__a21oi_1
X_15596_ _05838_ _05839_ vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__nand2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _07681_ _07682_ _07680_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__a21bo_1
X_14547_ _04639_ _04641_ _04770_ vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__nor3_1
X_11759_ _01849_ _01851_ vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__or2_4
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17266_ _07720_ _07726_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__xor2_1
X_14478_ _04695_ _04696_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16217_ _01106_ _06585_ _07646_ vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19005_ clknet_4_7_0_clk _09372_ vssd1 vssd1 vccd1 vccd1 salida\[58\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13429_ _03096_ _03103_ _03047_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__mux2_1
X_17197_ _07651_ vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16148_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16079_ _00167_ _00214_ _06435_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__and3_1
XFILLER_0_11_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput1 buttons vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_4
X_09522_ _04187_ _04285_ _04296_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09453_ _03443_ _03487_ _03542_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__nand3_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _00174_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__buf_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12800_ _02869_ _02880_ _02879_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__a21o_1
X_13780_ _03531_ _03509_ _08746_ _08049_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__nand4_2
X_10992_ _07058_ _07091_ _00460_ _05856_ _01084_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__a41o_1
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12731_ _02814_ _02817_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__and2_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _05739_ _05754_ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _07788_ _00120_ _00132_ _09219_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__and4_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _03005_ _00399_ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__nand2_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _01640_ _01641_ _01564_ _01604_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15381_ _05679_ _05680_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12593_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel _00180_ _02685_
+ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _07565_ _07566_ _07567_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__nand3_1
X_14332_ _04489_ _04490_ _04535_ _04536_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and4_2
X_11544_ _01633_ _01634_ _01635_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17051_ _07485_ _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _04283_ _04429_ _04459_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__or3_2
XFILLER_0_123_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11475_ _01565_ _01566_ _01567_ vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__nand3_1
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16002_ _07058_ _00193_ _06346_ _02358_ _02215_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__a311o_1
XFILLER_0_122_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ _00725_ _00730_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10426_ _00512_ _00518_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14194_ _04169_ net120 _04385_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__o211a_4
XFILLER_0_104_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ _06029_ _06051_ _07384_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10357_ _00447_ _00448_ _00449_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__and3_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _03023_ _03167_ vssd1 vssd1 vccd1 vccd1 _03168_ sky130_fd_sc_hd__nand2_1
X_17953_ _07106_ _07621_ _08472_ _08473_ vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__o22a_1
X_10288_ _00233_ _00243_ vssd1 vssd1 vccd1 vccd1 _00381_ sky130_fd_sc_hd__or2_1
X_12027_ _02115_ net187 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__and2b_1
X_16904_ _07224_ _07226_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__nand2_1
X_17884_ _08380_ _08399_ vssd1 vssd1 vccd1 vccd1 _08401_ sky130_fd_sc_hd__nor2_1
X_16835_ _02476_ _02099_ _06510_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__and3_1
X_13978_ _03965_ _03978_ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16766_ _03912_ _06474_ vssd1 vssd1 vccd1 vccd1 _07183_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18505_ _03108_ _08150_ _09072_ _09042_ _09041_ vssd1 vssd1 vccd1 vccd1 _09073_ sky130_fd_sc_hd__a32o_1
X_15717_ _05966_ _06045_ vssd1 vssd1 vccd1 vccd1 _06046_ sky130_fd_sc_hd__xnor2_1
X_12929_ _03002_ _03021_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__nor2_2
X_16697_ _06563_ _06937_ _06961_ _07106_ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18436_ _08950_ _08952_ _08949_ vssd1 vssd1 vccd1 vccd1 _08999_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_8_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ _05909_ _05908_ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__and2b_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15579_ _00112_ _07384_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__and2_1
X_18367_ _02992_ _06512_ _03068_ vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17318_ _07647_ _07660_ _07645_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18298_ _02200_ _07780_ _08150_ _07650_ vssd1 vssd1 vccd1 vccd1 _08850_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17249_ _02059_ _07592_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__and2_2
XFILLER_0_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09505_ _03771_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__buf_6
XFILLER_0_94_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ cla_inst.in2\[17\] vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__buf_8
XFILLER_0_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_50 _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_61 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _06326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_83 _08345_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_94 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11260_ _01351_ _01352_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__nor2_2
X_10211_ _00291_ _00302_ _00301_ vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__o21ai_1
X_11191_ _01280_ _01283_ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__or2b_1
X_10142_ _00150_ _00153_ vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__nand2_1
X_10073_ _00165_ vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__buf_8
X_14950_ _01520_ _00502_ _07733_ _02984_ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__a22oi_4
X_13901_ _04062_ _04064_ vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__nand2_1
X_14881_ _05100_ _05013_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__o21a_1
X_13832_ _03987_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__inv_2
X_16620_ _06812_ _03003_ net211 vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__nor3_1
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ _06571_ _06874_ _06947_ _06542_ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__a2bb2o_1
X_13763_ _03913_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ _01062_ _01067_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _03014_ _01317_ _05762_ _05761_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__a31o_1
X_12714_ _02785_ _02806_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__and2_1
X_16482_ _06869_ _06872_ _05736_ vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__a21bo_2
X_13694_ cla_inst.in2\[24\] _00174_ _04471_ _03739_ vssd1 vssd1 vccd1 vccd1 _03840_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _05719_ _05644_ _05735_ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__nor3_1
X_18221_ _06399_ _06546_ vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12645_ _02700_ _02732_ _02731_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15364_ _02999_ _03153_ _05661_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__a21o_1
X_18152_ _06836_ _08678_ _08680_ _08685_ _08691_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__o311a_1
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12576_ _02634_ _02668_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__nand2_1
X_14315_ _04517_ _04518_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__nor2_1
X_17103_ _07434_ _07441_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11527_ _01610_ _01618_ _01617_ vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__o21a_1
X_18083_ _08459_ _08460_ _08540_ vssd1 vssd1 vccd1 vccd1 _08617_ sky130_fd_sc_hd__nand3_1
X_15295_ _05575_ _05576_ _05587_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__a21o_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17034_ _06739_ _06733_ _02978_ vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__mux2_1
X_14246_ _04434_ _04435_ _04441_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _01518_ _01523_ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10409_ cla_inst.in1\[30\] vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14177_ _04359_ _04367_ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _01474_ _01481_ vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__xnor2_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _03221_ _03222_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__and3_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ clknet_4_0_0_clk _09381_ vssd1 vssd1 vccd1 vccd1 salida\[38\] sky130_fd_sc_hd__dfxtp_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _08180_ _03150_ _03023_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__o21ai_1
X_17936_ _07664_ net145 vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__nand2_1
X_17867_ _08285_ _08280_ vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16818_ _07237_ _07238_ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__or2_1
X_17798_ _07038_ _07859_ _08306_ vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16749_ _07162_ _02831_ _07163_ vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18419_ _08979_ _08980_ vssd1 vssd1 vccd1 vccd1 _08981_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _07788_ _09248_ _09263_ vssd1 vssd1 vccd1 vccd1 _09271_ sky130_fd_sc_hd__nand3_1
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_157 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_157/HI led_enb[6] sky130_fd_sc_hd__conb_1
X_10760_ _06181_ _00822_ _00797_ _00821_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ sel_op\[2\] vssd1 vssd1 vccd1 vccd1 _03184_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10691_ _04722_ _00782_ _00780_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12430_ _02515_ net122 _02456_ _02522_ vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12361_ _02452_ _02453_ vssd1 vssd1 vccd1 vccd1 _02454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14100_ _04267_ _04268_ _04282_ vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__o21a_2
X_11312_ _01396_ _01397_ _01398_ _01404_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__o31a_1
X_15080_ _00151_ _00125_ _05964_ _06062_ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__and4_1
X_12292_ _02352_ net323 _02282_ _02384_ vssd1 vssd1 vccd1 vccd1 _02385_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14031_ _04192_ _04193_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__a21o_1
X_11243_ _01332_ _01333_ _01334_ _01312_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_30_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11174_ _01141_ _01266_ vssd1 vssd1 vccd1 vccd1 _01267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _00217_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__clkbuf_8
X_18770_ _09285_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__buf_1
X_15982_ _02992_ _03068_ vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nand2_1
X_17721_ _08220_ _08221_ _08218_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__o21ai_1
X_10056_ cla_inst.in2\[26\] vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__clkbuf_4
X_14933_ _05190_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__xor2_1
X_17652_ _08147_ vssd1 vssd1 vccd1 vccd1 _09394_ sky130_fd_sc_hd__inv_2
X_14864_ _05116_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16603_ _03169_ _06432_ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__or2_1
X_13815_ _03970_ _03971_ vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14795_ _05041_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__xnor2_1
X_17583_ _08070_ _08072_ vssd1 vssd1 vccd1 vccd1 _08073_ sky130_fd_sc_hd__xor2_1
X_13746_ _03895_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__xnor2_4
X_16534_ _02975_ _03120_ _03927_ _06919_ _06930_ vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10958_ _00941_ _00953_ _00954_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__or3_4
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13677_ _03818_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__inv_2
X_16465_ _06680_ _06855_ vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10889_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _00982_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18204_ _08745_ _08747_ _08741_ vssd1 vssd1 vccd1 vccd1 _08749_ sky130_fd_sc_hd__a21o_1
X_15416_ _05545_ _05642_ vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__and2b_1
X_12628_ _07700_ _00131_ _02720_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__nand3_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16396_ _02780_ _01248_ _06673_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15347_ _05563_ _05630_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18135_ _01998_ _08673_ vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_124_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12559_ _02644_ _02645_ _02651_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15278_ _05463_ _05471_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__a21oi_1
X_18066_ _04647_ _06445_ vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__nand2_1
Xhold106 net101 vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold117 _00024_ vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold128 net89 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _04387_ _04388_ _04389_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__or3_4
Xhold139 _00005_ vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _02840_ _07353_ vssd1 vssd1 vccd1 vccd1 _07456_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ cla_inst.in1\[26\] vssd1 vssd1 vccd1 vccd1 _07004_ sky130_fd_sc_hd__clkbuf_4
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18968_ clknet_4_4_0_clk _09399_ vssd1 vssd1 vccd1 vccd1 salida\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _04337_ _06389_ _06390_ _08438_ vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ clknet_4_12_0_clk _00053_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09968_ _09070_ _09137_ vssd1 vssd1 vccd1 vccd1 _09145_ sky130_fd_sc_hd__xnor2_2
X_09899_ _04395_ vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__buf_6
X_11930_ _02016_ _02021_ _02022_ vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__o21a_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _00832_ _04482_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13600_ _03523_ _03525_ vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__nor2_2
X_10812_ _00900_ _00904_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__nor2_1
X_14580_ _04672_ _04674_ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2_2
X_11792_ _01564_ _01601_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13531_ _08865_ _00665_ _03413_ _03412_ _00495_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__a32o_1
XFILLER_0_83_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10743_ _07058_ _07091_ _05975_ _06094_ _00835_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__a41o_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16250_ _03027_ _03111_ _01674_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__a21o_1
X_13462_ _03434_ _03435_ _03466_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__nor3_1
XFILLER_0_152_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _03728_ _04143_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ _05483_ _05484_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__xnor2_2
X_12413_ _02505_ _00247_ _00166_ _00845_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16181_ _06419_ _06459_ vssd1 vssd1 vccd1 vccd1 _06547_ sky130_fd_sc_hd__nor2_2
X_13393_ _03507_ _03508_ _03490_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15132_ _02959_ _02962_ _04403_ _05409_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__a211o_4
X_12344_ _02436_ _02371_ vssd1 vssd1 vccd1 vccd1 _02437_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15063_ _05332_ _00461_ _00362_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__and4b_1
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12275_ _02353_ _02367_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14014_ _00164_ _01695_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__nand2_2
X_11226_ _07058_ _07091_ _06094_ _00460_ _01089_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__a41o_1
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18822_ _09125_ _09325_ vssd1 vssd1 vccd1 vccd1 _09327_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ _01247_ _01249_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__xnor2_4
X_10108_ _00190_ _00192_ _00193_ _00132_ _00200_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__a41o_1
X_18753_ _09272_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__clkbuf_1
X_11088_ _01166_ net144 _01179_ _01180_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__o211ai_4
X_15965_ _06299_ _06301_ _06312_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__nand3_1
X_17704_ _08083_ _08098_ _08204_ vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__a21o_1
X_14916_ _05173_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__xnor2_1
X_10039_ _00131_ vssd1 vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__clkbuf_8
X_18684_ net42 _09189_ _09220_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__o21a_1
X_15896_ _06195_ _06199_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17635_ _01866_ _06510_ _02988_ vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__and3b_1
X_14847_ _03539_ _04241_ _04079_ _05098_ vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17566_ _08052_ _08053_ vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__xor2_1
X_14778_ _09353_ _04336_ _05020_ _05021_ vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16517_ _06908_ _06909_ _06910_ vssd1 vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__nor3_1
X_13729_ _03875_ _03876_ _03856_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17497_ _07977_ _07978_ vssd1 vssd1 vccd1 vccd1 _07979_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16448_ _01264_ _06673_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16379_ _06758_ _06761_ _00134_ vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__o21a_2
XFILLER_0_53_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18118_ _08556_ _08559_ _08488_ vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18049_ _08391_ _08493_ _08579_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09822_ _07559_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__buf_4
X_09753_ _06558_ _06569_ _06808_ vssd1 vssd1 vccd1 vccd1 _06819_ sky130_fd_sc_hd__a21o_2
X_09684_ _06040_ _06051_ _06062_ _05257_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__and4_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10390_ _00468_ _00469_ _00481_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__nand3_2
XFILLER_0_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ _02052_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__o21ai_1
X_11011_ _01093_ _01103_ vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__xor2_1
X_12962_ _00119_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__clkbuf_4
X_15750_ _06074_ _06080_ vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__nand2_1
X_14701_ _04938_ _04832_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__and2b_1
X_11913_ _01911_ _02005_ vssd1 vssd1 vccd1 vccd1 _02006_ sky130_fd_sc_hd__xnor2_1
X_12893_ _03574_ vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__clkbuf_8
X_15681_ _06004_ _06005_ _05956_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__o21a_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _07771_ _07782_ _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__a21bo_1
X_14632_ _04730_ _04833_ _04862_ _04863_ vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11844_ _01933_ _01934_ _01935_ vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__nand3_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _04619_ _04789_ vssd1 vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__xor2_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _07796_ _07800_ _07819_ _06723_ _02045_ vssd1 vssd1 vccd1 vccd1 _09391_ sky130_fd_sc_hd__o32a_1
X_11775_ _01675_ _01864_ vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__nor2_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16302_ _03077_ _03029_ _02809_ vssd1 vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__a21o_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13514_ _03639_ _03641_ _03624_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__a21oi_2
X_10726_ _00817_ _00818_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__nand2_1
X_14494_ _03793_ _07722_ _08169_ _03859_ vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__a22oi_1
X_17282_ _02045_ _07743_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__nor2_4
XFILLER_0_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16233_ _06462_ _06603_ vssd1 vssd1 vccd1 vccd1 _06604_ sky130_fd_sc_hd__nor2_1
X_13445_ _03090_ _03137_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10657_ _00747_ _00748_ _00749_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__or3_4
XFILLER_0_35_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ _03317_ _03331_ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16164_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__buf_4
X_10588_ _00358_ _07504_ _00147_ _00131_ vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__and4_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15115_ _05390_ _05391_ vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__nor2_1
X_12327_ _07069_ _00774_ _00909_ _07036_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16095_ _03921_ _05420_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15046_ _02984_ _02988_ _00509_ _09248_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__and4_2
X_12258_ _02224_ _02225_ _02227_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__o21ai_1
X_11209_ _01300_ _01301_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__xor2_2
X_12189_ _02231_ _02279_ _02280_ _02281_ vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__or4_4
X_18805_ _09313_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__buf_1
X_16997_ _07432_ _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__xnor2_1
X_18736_ _04241_ net60 _09251_ vssd1 vssd1 vccd1 vccd1 _09259_ sky130_fd_sc_hd__mux2_1
X_15948_ _03921_ _06292_ _06294_ vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__a21o_1
X_18667_ net66 _09189_ _09208_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15879_ _06219_ _06220_ vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _08103_ _08110_ vssd1 vssd1 vccd1 vccd1 _08111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18598_ net255 _09140_ _09155_ _09144_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17549_ _03536_ _06483_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__nand2_2
XFILLER_0_129_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09805_ _07374_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09736_ _06602_ _06624_ vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__and2b_1
X_09667_ _05878_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09598_ _05115_ _05126_ vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__xnor2_2
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11560_ _01649_ _01651_ _01650_ vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10511_ _03596_ _00439_ _04395_ _03629_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11491_ _01573_ _01574_ _01580_ vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13230_ _03315_ _00735_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_107_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _00491_ _00532_ _00533_ _00534_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__nand4_4
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13161_ _03256_ _03257_ _03242_ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a21oi_1
X_10373_ _00450_ _00464_ _00463_ vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12112_ _05399_ _05355_ _07548_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__and3_1
X_13092_ _01677_ _03180_ _03183_ vssd1 vssd1 vccd1 vccd1 _03185_ sky130_fd_sc_hd__o21ai_1
X_12043_ _02073_ _02075_ _02076_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__or3_1
X_16920_ _07347_ _07348_ _06649_ vssd1 vssd1 vccd1 vccd1 _07350_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16851_ _02476_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__a21o_1
X_15802_ _06071_ _06082_ vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__nand2_1
X_16782_ _06937_ _07143_ _07198_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__or3_1
X_13994_ _03984_ _04002_ vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__or2_1
X_18521_ _06543_ _06453_ _09084_ _09089_ vssd1 vssd1 vccd1 vccd1 _09090_ sky130_fd_sc_hd__a31o_1
X_15733_ _06061_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__xor2_1
X_12945_ _03036_ _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18452_ _06649_ _09014_ _09015_ vssd1 vssd1 vccd1 vccd1 _09017_ sky130_fd_sc_hd__and3_1
X_15664_ _05970_ _05971_ _05988_ vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__o21ai_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 _06765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__buf_8
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_151 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _07855_ _07876_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_162 _08934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14615_ _04844_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_173 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18383_ _06426_ _06449_ _08935_ _08939_ _08942_ vssd1 vssd1 vccd1 vccd1 _08943_ sky130_fd_sc_hd__o311a_1
X_11827_ _01831_ _01829_ _01830_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__and3_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15595_ _05912_ _05913_ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _03311_ _07355_ _02200_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__or3b_1
X_14546_ _04639_ _04641_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__o21a_1
X_11758_ _01849_ _01850_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03914_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and4b_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _06138_ _00800_ _00799_ vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17265_ _07724_ _07725_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__xnor2_1
X_14477_ _04691_ _04694_ _02969_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__a21o_1
X_11689_ _01771_ _01780_ _01779_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19004_ clknet_4_7_0_clk _09371_ vssd1 vssd1 vccd1 vccd1 salida\[57\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16216_ op_code\[0\] op_code\[3\] op_code\[2\] op_code\[1\] vssd1 vssd1 vccd1 vccd1
+ _06585_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_11_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13428_ _03088_ _03093_ _03047_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__mux2_1
X_17196_ _07510_ _07529_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13359_ _00183_ _04864_ _04143_ _00184_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a22oi_1
X_16147_ _06509_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16078_ _02214_ _06434_ vssd1 vssd1 vccd1 vccd1 _06435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15029_ _05296_ _05297_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2_1
Xinput2 i_wb_addr[0] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_09521_ _04198_ _04209_ _04274_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__nand3_1
XFILLER_0_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18719_ _09125_ vssd1 vssd1 vccd1 vccd1 _09245_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09452_ _03509_ _03410_ _03432_ _03531_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__a22o_1
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _06384_ _06439_ vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__xnor2_2
X_10991_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _05617_ _01080_
+ _01083_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__and4_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _02807_ _02822_ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__and2_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _02713_ _02715_ vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _04463_ _04466_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__nor2_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11612_ _01702_ _01703_ _01669_ _01681_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _03009_ _07668_ _01139_ _01223_ vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12592_ ApproximateM_inst.lob_16.lob2.mux.sel net185 vssd1 vssd1 vccd1 vccd1 _02685_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14331_ _04533_ _04534_ _04491_ _04378_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__a211o_1
X_11543_ _01633_ _01634_ _01635_ vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__nand3_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14262_ _04283_ _04429_ _04459_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__o21ai_4
X_17050_ _07488_ _07490_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__nand2_1
X_11474_ _05464_ _04056_ _00563_ _05508_ vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13213_ _00733_ vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__inv_2
X_16001_ _06342_ _06347_ _06348_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_ sky130_fd_sc_hd__and4b_1
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10425_ _07853_ _00513_ _00517_ _00353_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__a31oi_2
X_14193_ _04382_ _04383_ _04334_ vssd1 vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ _00622_ _00629_ _00628_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__a21o_1
X_10356_ _00286_ _00287_ _00281_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_131_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _03166_ _01248_ _03028_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__mux2_1
X_17952_ _08472_ _08473_ _07109_ _07623_ vssd1 vssd1 vccd1 vccd1 _08475_ sky130_fd_sc_hd__and4bb_1
X_10287_ _00234_ _00242_ vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12026_ _02115_ _02118_ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__xnor2_1
X_16903_ _07126_ vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__clkbuf_4
X_17883_ _08380_ _08399_ vssd1 vssd1 vccd1 vccd1 _08400_ sky130_fd_sc_hd__and2_1
X_16834_ _02476_ _06510_ _02099_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16765_ _06680_ _07175_ _07177_ _07181_ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__or4b_2
X_13977_ _03967_ _03977_ vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18504_ _04853_ _09039_ vssd1 vssd1 vccd1 vccd1 _09072_ sky130_fd_sc_hd__nand2_1
X_15716_ _06035_ _06044_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__xor2_1
X_12928_ _03003_ net212 _03017_ _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__or4_4
XFILLER_0_87_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16696_ _02533_ _07104_ _07105_ vssd1 vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__nand3_4
XFILLER_0_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18435_ _06408_ _06463_ _08998_ vssd1 vssd1 vccd1 vccd1 _09406_ sky130_fd_sc_hd__a21oi_1
X_15647_ _05855_ _05907_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__and2b_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _02942_ _02947_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__or2b_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18366_ _06649_ _08922_ _08923_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__and3_1
X_15578_ _05449_ _00119_ _05850_ _05849_ vssd1 vssd1 vccd1 vccd1 _05895_ sky130_fd_sc_hd__a31o_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17317_ _07771_ _07782_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__xnor2_1
X_14529_ _04750_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18297_ _07665_ _07650_ _07708_ _08150_ _08848_ vssd1 vssd1 vccd1 vccd1 _08849_ sky130_fd_sc_hd__a41o_1
XFILLER_0_43_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17248_ _06562_ _06756_ _07410_ _07706_ vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__or4_4
XFILLER_0_114_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17179_ _07631_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _04034_ _04045_ _04067_ _04099_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_154_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09435_ _03345_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__clkbuf_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_40 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_62 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_73 _06482_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_84 _08615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_95 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _00291_ _00301_ _00302_ vssd1 vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__or3_4
X_11190_ _01281_ _01282_ vssd1 vssd1 vccd1 vccd1 _01283_ sky130_fd_sc_hd__xnor2_1
X_10141_ _07690_ _07842_ _07864_ _07831_ vssd1 vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10072_ _03673_ vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__buf_6
XFILLER_0_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13900_ _04062_ _04064_ vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__or2_1
X_14880_ _05123_ _05134_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__xnor2_1
X_13831_ _03987_ _04154_ _07526_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__and4b_1
X_16550_ _06946_ vssd1 vssd1 vccd1 vccd1 _06947_ sky130_fd_sc_hd__clkbuf_4
X_10974_ _01063_ _01066_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__xor2_2
X_13762_ _03908_ _03911_ _03913_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__mux2_1
X_15501_ _01356_ _09059_ _05724_ _05723_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__a31o_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12713_ _07788_ _07613_ _02805_ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__and3_1
X_16481_ _03184_ _06575_ _06871_ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__a21o_1
X_13693_ _00174_ _04395_ _04657_ _00184_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__a22oi_1
X_18220_ _02994_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__a21oi_1
X_15432_ _05719_ _05644_ _05735_ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__o21a_1
X_12644_ _02735_ _02736_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18151_ _03120_ _06021_ _08687_ _08690_ vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15363_ _02999_ _03153_ _05661_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__nand3_1
X_12575_ _02655_ _02666_ _02667_ vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17102_ _07546_ _07547_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__nand2_1
X_14314_ _00112_ _09350_ _01005_ _08409_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11526_ _01610_ _01617_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nor3_4
XFILLER_0_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18082_ _08563_ _08564_ vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15294_ _05585_ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _04247_ _06727_ vssd1 vssd1 vccd1 vccd1 _07474_ sky130_fd_sc_hd__nand2_1
X_14245_ _04434_ _04435_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__nand3_1
X_11457_ _01548_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10408_ _00499_ _00500_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__nor2_1
X_14176_ _04360_ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__xnor2_1
X_11388_ _01479_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__nor2_2
XFILLER_0_110_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _03651_ _03662_ _04460_ _04657_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__nand4_2
X_13127_ _00611_ _00616_ _00610_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a21bo_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ clknet_4_3_0_clk _09380_ vssd1 vssd1 vccd1 vccd1 salida\[37\] sky130_fd_sc_hd__dfxtp_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _03025_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__and2_1
X_17935_ _08454_ _08455_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12009_ _02092_ _02097_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__or2b_1
X_17866_ _08304_ _08305_ _08307_ vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16817_ _07235_ _07236_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__nor2_1
X_17797_ _08304_ _08305_ vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__xor2_1
X_16748_ _07162_ _02831_ _04238_ vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16679_ _07087_ vssd1 vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18418_ _06408_ _08428_ _03016_ vssd1 vssd1 vccd1 vccd1 _08980_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18349_ _08904_ _08852_ _08851_ vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput60 i_wb_data[3] vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__buf_2
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09984_ _07799_ _09256_ vssd1 vssd1 vccd1 vccd1 _09263_ sky130_fd_sc_hd__and2_4
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_158 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_158/HI led_enb[7] sky130_fd_sc_hd__conb_1
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _04722_ _00780_ _00782_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12360_ _02375_ _02443_ _02445_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__or3_1
XFILLER_0_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11311_ _01401_ _01403_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__xor2_1
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _02279_ _02280_ _02281_ _02231_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_121_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14030_ _04195_ _04206_ vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11242_ _01312_ _01332_ _01333_ _01334_ vssd1 vssd1 vccd1 vccd1 _01335_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11173_ _01263_ _01265_ vssd1 vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__xor2_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10124_ _04242_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__clkbuf_4
X_15981_ _03013_ _03073_ vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _08218_ _08220_ _08221_ vssd1 vssd1 vccd1 vccd1 _08222_ sky130_fd_sc_hd__or3_1
X_10055_ cla_inst.in2\[27\] vssd1 vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__clkbuf_4
X_14932_ _05191_ _05054_ _05051_ vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__o21ai_1
X_17651_ _08124_ _08128_ _08146_ _06463_ _03111_ vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__a32o_1
X_14863_ _04977_ _04980_ _04978_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__o21ba_1
X_16602_ _03921_ _06998_ _07003_ _06484_ vssd1 vssd1 vccd1 vccd1 _07005_ sky130_fd_sc_hd__o211a_1
X_13814_ _05279_ _05355_ cla_inst.in1\[29\] cla_inst.in1\[28\] vssd1 vssd1 vccd1 vccd1
+ _03971_ sky130_fd_sc_hd__and4_1
X_17582_ _07109_ net146 vssd1 vssd1 vccd1 vccd1 _08072_ sky130_fd_sc_hd__nand2_1
X_14794_ _01505_ _05758_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__nand2_1
X_16533_ _06923_ _06925_ _06929_ _06720_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__and4b_1
X_13745_ _03725_ _03726_ _03724_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__o21ba_2
X_10957_ _01039_ _01048_ _01049_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__nor3_1
XFILLER_0_85_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16464_ _06348_ _06545_ _06854_ _03166_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__a22o_1
X_13676_ _03818_ _00563_ cla_inst.in2\[28\] _03819_ vssd1 vssd1 vccd1 vccd1 _03820_
+ sky130_fd_sc_hd__and4b_1
X_10888_ _05213_ _04460_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__nand2_1
X_18203_ _08741_ _08745_ _08747_ _03195_ vssd1 vssd1 vccd1 vccd1 _08748_ sky130_fd_sc_hd__a31o_1
X_15415_ _05651_ _05670_ vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ _07799_ _00181_ vssd1 vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__and2_2
XFILLER_0_54_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16395_ _02780_ _06673_ _01248_ vssd1 vssd1 vccd1 vccd1 _06780_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18134_ _01997_ _08593_ _01995_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__o21a_1
X_15346_ _05545_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12558_ _02648_ _02649_ _02650_ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18065_ _04887_ _06394_ _06393_ vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__a21o_1
X_11509_ _01593_ _01600_ _01585_ _01586_ vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__o211ai_4
X_15277_ _05470_ _05465_ vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ _02574_ _02580_ _02581_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__nor3_1
Xhold107 _00030_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 net98 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _02839_ _07454_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__nor2_1
Xhold129 _00019_ vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14228_ _04387_ vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _01745_ _01695_ _04346_ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__a21o_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ clknet_4_4_0_clk _09398_ vssd1 vssd1 vccd1 vccd1 salida\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _06420_ _08437_ vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18898_ clknet_4_12_0_clk _00052_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[16\] sky130_fd_sc_hd__dfxtp_2
X_17849_ _08356_ _08361_ vssd1 vssd1 vccd1 vccd1 _08362_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09967_ _09080_ _09131_ vssd1 vssd1 vccd1 vccd1 _09137_ sky130_fd_sc_hd__xor2_2
X_09898_ _08365_ _08376_ _08387_ vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__nand3_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _01950_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _00900_ _00902_ _00903_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__nor3_1
X_11791_ _01841_ _01881_ _01882_ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__nand4_2
XFILLER_0_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13530_ _03653_ _03659_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__xor2_2
XFILLER_0_94_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10742_ _00832_ _05704_ _00833_ _00834_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10673_ _03673_ _00764_ _00765_ vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__a21bo_1
X_13461_ _03573_ _03583_ _02976_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _01505_ _09059_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__nand2_1
X_12412_ _00120_ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__buf_4
X_16180_ _06545_ vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__buf_4
X_13392_ _03490_ _03507_ _03508_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__nand3b_4
XFILLER_0_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15131_ _04947_ net117 vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ _07788_ _00120_ _04067_ _00166_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__and4_2
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15062_ _07504_ _05845_ _05878_ _00679_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__a22o_1
X_12274_ _02356_ _02365_ _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14013_ _04186_ _04188_ vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__nor2_2
X_11225_ _00846_ _01317_ _00861_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__a21oi_2
X_11156_ cla_inst.in2\[20\] _01248_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nand2_2
X_18821_ _03011_ net58 _09250_ vssd1 vssd1 vccd1 vccd1 _09325_ sky130_fd_sc_hd__mux2_1
X_10107_ _00170_ _00194_ _00198_ _00199_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__and4_1
X_18752_ _09245_ _09270_ vssd1 vssd1 vccd1 vccd1 _09272_ sky130_fd_sc_hd__and2_1
X_11087_ _01039_ _01049_ _01048_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__o21ai_2
X_15964_ _06308_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__xnor2_1
X_17703_ _08079_ _08081_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__and2_1
X_14915_ _05047_ _05048_ _05046_ vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__o21ai_1
X_10038_ _00130_ vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__clkbuf_8
X_18683_ _01862_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09220_ sky130_fd_sc_hd__a21oi_1
X_15895_ _06237_ _06208_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__nand2_1
X_17634_ _02988_ _06510_ _03111_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__a21bo_1
X_14846_ _03117_ _05097_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17565_ _07935_ _07937_ _07934_ _06800_ vssd1 vssd1 vccd1 vccd1 _08053_ sky130_fd_sc_hd__a2bb2o_1
X_14777_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11989_ _05017_ _00131_ vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16516_ _06908_ _06909_ _06910_ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ _03856_ _03875_ _03876_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__or3_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _06579_ _07124_ _07511_ _07861_ vssd1 vssd1 vccd1 vccd1 _07978_ sky130_fd_sc_hd__or4_4
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16447_ _06589_ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13659_ _03797_ _03798_ _03799_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16378_ _03313_ _06760_ vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18117_ _08652_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15329_ _03534_ _03556_ _03536_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18048_ _08486_ _08492_ vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09821_ _07548_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__clkbuf_8
X_09752_ _06667_ _06798_ vssd1 vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__xnor2_1
X_09683_ _05617_ vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__buf_4
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11010_ _01097_ _01101_ _01102_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12961_ _03024_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__nand2_1
X_14700_ _04832_ _04938_ vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__and2b_1
X_11912_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _00180_ vssd1
+ vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__nand2_1
X_15680_ _05956_ _06004_ _06005_ vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nor3_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _02984_ vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__buf_4
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ _04860_ _04861_ _04723_ _04834_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__a211oi_4
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _01933_ _01934_ _01935_ vssd1 vssd1 vccd1 vccd1 _01936_ sky130_fd_sc_hd__a21o_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _07256_ _07804_ _07805_ _07818_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__a31o_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _04780_ _04787_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _00846_ _01866_ _01674_ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__a21oi_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16301_ _06672_ _06674_ _06675_ vssd1 vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__nand3_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _03624_ _03639_ _03641_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__and3_2
X_10725_ _00810_ _00816_ _00801_ _00802_ vssd1 vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__o211ai_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17281_ _06814_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__clkbuf_4
X_14493_ _04709_ _04710_ _04705_ _04706_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_634 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16232_ _06543_ _06429_ _06601_ _06546_ _06333_ vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__a32o_1
XFILLER_0_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13444_ _02982_ _03141_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__or2_1
X_10656_ _00578_ _00580_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16163_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _06528_ sky130_fd_sc_hd__or3_4
X_13375_ _03318_ _03330_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10587_ _00678_ _00147_ _00132_ _00679_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15114_ _05387_ _05389_ _05347_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__o21a_1
X_12326_ _07221_ _07243_ _04242_ _00176_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__and4_1
X_16094_ _06246_ _06452_ vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15045_ _02988_ _03455_ _09311_ _02984_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _02346_ _02349_ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11208_ _05878_ _00839_ _00838_ vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__a21bo_1
X_12188_ _02203_ _02229_ _02228_ vssd1 vssd1 vccd1 vccd1 _02281_ sky130_fd_sc_hd__o21a_1
X_18804_ _09298_ _09312_ vssd1 vssd1 vccd1 vccd1 _09313_ sky130_fd_sc_hd__and2_1
X_11139_ _01143_ _01230_ _01229_ _01196_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__a211oi_2
X_16996_ _07300_ _07327_ _07298_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__o21a_1
X_18735_ _09258_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__clkbuf_1
X_15947_ _03537_ _06293_ _03123_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a21o_1
X_18666_ _02099_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09208_ sky130_fd_sc_hd__a21oi_1
X_15878_ _06193_ _06175_ _06218_ vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__or3_1
X_17617_ _08108_ _08109_ vssd1 vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__nor2_1
X_14829_ _05077_ _05079_ vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18597_ salida\[18\] _09141_ _09142_ salida\[50\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09155_ sky130_fd_sc_hd__a221o_1
X_17548_ _06378_ _06546_ _08034_ _03693_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17479_ _07957_ _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09804_ cla_inst.in1\[27\] vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__clkbuf_4
X_09735_ _05355_ _06613_ net231 _05399_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09666_ _05388_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _04526_ _04602_ _04406_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ _00450_ _00463_ _00464_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__nor3_1
XFILLER_0_108_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11490_ _01582_ _01538_ _01534_ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _00489_ _00490_ net184 net340 vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__a211o_2
XFILLER_0_135_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _00450_ _00463_ _00464_ vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__or3_4
X_13160_ _03242_ _03256_ _03257_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ _05235_ _00147_ _02179_ _02180_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__a22oi_2
X_13091_ _03047_ _03182_ vssd1 vssd1 vccd1 vccd1 _03183_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12042_ _02107_ _02134_ _02049_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__o21ai_2
X_16850_ _06422_ _06459_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__or2_2
X_15801_ _06135_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__nor2_1
X_16781_ _07196_ _07197_ vssd1 vssd1 vccd1 vccd1 _07198_ sky130_fd_sc_hd__xnor2_1
X_13993_ _04146_ _04147_ _04164_ vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or3_1
X_18520_ _03120_ _06325_ _09088_ vssd1 vssd1 vccd1 vccd1 _09089_ sky130_fd_sc_hd__o21ai_1
X_15732_ _06000_ _06002_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__nand2_1
X_12944_ _02728_ _02965_ _03292_ _03217_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18451_ _08969_ _08978_ _09013_ vssd1 vssd1 vccd1 vccd1 _09015_ sky130_fd_sc_hd__o21ai_1
X_15663_ _05985_ _05987_ vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__nor2_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 _04132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _02967_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_141 _07091_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _07858_ _07874_ vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__xnor2_1
XANTENNA_152 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _03859_ _03793_ _07755_ cla_inst.in1\[28\] vssd1 vssd1 vccd1 vccd1 _04845_
+ sky130_fd_sc_hd__and4_4
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _05896_ _06407_ _06421_ _08940_ vssd1 vssd1 vccd1 vccd1 _08942_ sky130_fd_sc_hd__o211ai_1
XANTENNA_163 _08934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _01917_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__nand2_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _05894_ _05825_ _05911_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__nor3_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _02200_ _06510_ _02045_ vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__a21o_1
X_14545_ _04768_ _04769_ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__and2_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _05584_ _03388_ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ _06008_ vssd1 vssd1 vccd1 vccd1 _01850_ sky130_fd_sc_hd__a22o_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10708_ _06138_ _00799_ _00800_ vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__nand3_2
X_17264_ _07042_ _07106_ vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__nor2_1
X_14476_ _04691_ _04694_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11688_ _01771_ _01779_ _01780_ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__nor3_4
XFILLER_0_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19003_ clknet_4_5_0_clk _09370_ vssd1 vssd1 vccd1 vccd1 salida\[56\] sky130_fd_sc_hd__dfxtp_1
X_16215_ _06561_ _06572_ _06581_ _06563_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__o22a_1
X_13427_ _03544_ _03546_ _03547_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__mux2_1
X_10639_ _00724_ _00731_ vssd1 vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17195_ _07649_ vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16146_ _03239_ op_code\[3\] op_code\[2\] _03217_ vssd1 vssd1 vccd1 vccd1 _06509_
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13358_ _03267_ _03290_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12309_ _00645_ _05235_ _07570_ _07602_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__and4_2
X_16077_ _06433_ vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__inv_2
X_13289_ _03728_ _00459_ _03216_ _03215_ _05845_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__a32o_1
X_15028_ _05207_ _05176_ _05295_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__and3_1
XFILLER_0_20_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 i_wb_addr[10] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16979_ _06579_ _07313_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__or2_1
X_09520_ _04198_ _04209_ _04274_ vssd1 vssd1 vccd1 vccd1 _04285_ sky130_fd_sc_hd__a21o_1
X_18718_ _09244_ vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__clkbuf_1
X_09451_ _03520_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__buf_8
X_18649_ _09176_ _09194_ vssd1 vssd1 vccd1 vccd1 _09195_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _06395_ _06428_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__xnor2_2
X_10990_ _01081_ cla_inst.in1\[20\] net233 _01082_ vssd1 vssd1 vccd1 vccd1 _01083_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09649_ cla_inst.in1\[23\] vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _02724_ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__inv_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _01669_ _01681_ _01702_ _01703_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12591_ _02674_ _02682_ _02681_ vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14330_ _04491_ _04378_ _04533_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _01573_ _01581_ vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14261_ _04457_ _04458_ vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__nor2_2
X_11473_ _05224_ _04143_ vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16000_ _02972_ _01264_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__nand2_1
X_13212_ _03310_ _03312_ vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__xor2_2
XFILLER_0_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10424_ _00515_ _00516_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__nor2_4
XFILLER_0_123_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14192_ _04334_ _04382_ _04383_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__nand3_4
XFILLER_0_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13143_ _03237_ _03238_ _00620_ net136 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a211o_1
X_10355_ _00438_ _00446_ _00445_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__a21o_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _09339_ vssd1 vssd1 vccd1 vccd1 _00379_ sky130_fd_sc_hd__inv_2
X_13074_ _01264_ vssd1 vssd1 vccd1 vccd1 _03166_ sky130_fd_sc_hd__clkbuf_4
X_17951_ _07394_ _07604_ _07649_ _07780_ vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__and4_1
X_12025_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__xnor2_2
X_16902_ _07328_ _07329_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__xnor2_1
X_17882_ _08397_ vssd1 vssd1 vccd1 vccd1 _08399_ sky130_fd_sc_hd__inv_2
X_16833_ _06508_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__buf_4
X_16764_ _06424_ _07179_ _07180_ vssd1 vssd1 vccd1 vccd1 _07181_ sky130_fd_sc_hd__or3_1
X_13976_ _03792_ _03995_ vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15715_ _06036_ _06043_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__xnor2_1
X_18503_ _09051_ _09057_ _09071_ _06463_ _03155_ vssd1 vssd1 vccd1 vccd1 _09409_ sky130_fd_sc_hd__a32oi_2
X_12927_ _03018_ _03019_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__or2_1
X_16695_ _06812_ _06575_ _06871_ vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__o21ai_4
X_15646_ _05914_ _05926_ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and2_1
X_18434_ _06559_ _08977_ _08978_ _08997_ vssd1 vssd1 vccd1 vccd1 _08998_ sky130_fd_sc_hd__o31a_1
X_12858_ _02949_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__or2_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _01900_ _01899_ _01812_ _01811_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__o211ai_1
X_18365_ _08873_ _08893_ _08921_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__o21ai_1
X_15577_ _05767_ _05822_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12789_ _02871_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _07779_ _07781_ vssd1 vssd1 vccd1 vccd1 _07782_ sky130_fd_sc_hd__xnor2_2
X_14528_ _04743_ _04749_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18296_ _04023_ _07516_ _08260_ vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__or3_2
XFILLER_0_126_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17247_ _02059_ _06889_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__nand2_4
X_14459_ _04628_ _04629_ _04674_ _04675_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17178_ _06944_ _06957_ _07115_ _07035_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16129_ _08180_ _03144_ vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _04088_ vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09434_ cla_inst.in2\[19\] vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__buf_6
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_30 _01225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_41 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_63 _04414_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_74 _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_85 _08750_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_96 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10140_ _00144_ _00155_ vssd1 vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__nand2_1
X_10071_ _00163_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__clkbuf_8
X_13830_ _09172_ _03673_ _00211_ _09166_ vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13761_ _03912_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__buf_4
X_10973_ _00439_ _01064_ _01065_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__a21bo_1
X_15500_ _05734_ _05733_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12712_ _00120_ _07559_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__and2_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16480_ _06870_ vssd1 vssd1 vccd1 vccd1 _06871_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13692_ _03669_ _03652_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15431_ _05733_ _05734_ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__xnor2_1
X_12643_ _02689_ _02734_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18150_ _07089_ _08141_ _08689_ _06721_ vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15362_ _05658_ _05659_ vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12574_ _02656_ _02665_ vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__and2b_1
X_17101_ _07536_ _07538_ _07545_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14313_ _03321_ _01005_ _01575_ _03322_ vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11525_ _01607_ _01608_ _01609_ vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18081_ _08502_ _08585_ vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15293_ _02999_ _03071_ _05583_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__a21o_1
X_17032_ _06680_ _07471_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14244_ _04439_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11456_ _01527_ _01529_ vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10407_ _07047_ _07080_ _09303_ _07722_ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__and4_1
X_14175_ _04364_ _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11387_ _01478_ _01475_ _01476_ vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__nor3_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13126_ _03213_ _03214_ _03220_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a21o_1
X_10338_ _00291_ _00301_ _00302_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__nor3_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ clknet_4_1_0_clk _09379_ vssd1 vssd1 vccd1 vccd1 salida\[36\] sky130_fd_sc_hd__dfxtp_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _00339_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__buf_4
X_17934_ _07751_ _07595_ _08453_ vssd1 vssd1 vccd1 vccd1 _08455_ sky130_fd_sc_hd__and3_1
X_10269_ _07526_ vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12008_ _02034_ _02100_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__nor2_1
X_17865_ _08378_ _08379_ vssd1 vssd1 vccd1 vccd1 _08380_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16816_ _07235_ _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__and2_1
X_17796_ _08190_ _08193_ _08189_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13959_ _03951_ _03959_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nand2_1
X_16747_ _02832_ _02801_ vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__and2b_1
X_16678_ _06726_ _06729_ _03098_ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18417_ _03016_ _06512_ _06408_ vssd1 vssd1 vccd1 vccd1 _08979_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15629_ _05796_ _05949_ _05950_ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_57_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18348_ _08847_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ _04238_ _08820_ _08824_ _08829_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 i_wb_data[23] vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_1
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 i_wb_data[4] vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_2
XFILLER_0_114_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ cla_inst.in1\[30\] vssd1 vssd1 vccd1 vccd1 _09256_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwb_buttons_leds_159 vssd1 vssd1 vccd1 vccd1 wb_buttons_leds_159/HI led_enb[8] sky130_fd_sc_hd__conb_1
XFILLER_0_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11310_ _01319_ _01323_ _01402_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12290_ _02352_ _02380_ _02381_ _02382_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__nor4_2
XFILLER_0_133_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11241_ _01310_ _01311_ net220 _01020_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__a211o_2
X_11172_ _00163_ _01264_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__nand2_2
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10123_ _00184_ _00183_ _00171_ _00177_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__and4_1
XFILLER_0_100_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15980_ _00908_ _02963_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14931_ _05036_ _05037_ _05049_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__and3_1
X_10054_ _00146_ vssd1 vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__buf_4
X_14862_ _05113_ _05114_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17650_ _08135_ _08138_ _08145_ vssd1 vssd1 vccd1 vccd1 _08146_ sky130_fd_sc_hd__and3_1
X_13813_ _05301_ _07755_ cla_inst.in1\[28\] _05410_ vssd1 vssd1 vccd1 vccd1 _03970_
+ sky130_fd_sc_hd__a22oi_1
X_16601_ _03921_ _07002_ vssd1 vssd1 vccd1 vccd1 _07003_ sky130_fd_sc_hd__nand2_1
X_17581_ _08068_ _08069_ vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__nand2_1
X_14793_ _05038_ _05040_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__nor2_1
X_16532_ _06344_ _06346_ _06926_ _06927_ _06598_ vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__a311o_1
X_13744_ _03893_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10956_ _01022_ _01023_ _01038_ vssd1 vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_57_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16463_ _02972_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__a21o_1
X_13675_ cla_inst.in2\[29\] _03432_ _00205_ cla_inst.in2\[30\] vssd1 vssd1 vccd1 vccd1
+ _03819_ sky130_fd_sc_hd__a22o_1
X_10887_ net195 _00955_ _00978_ _00979_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__o211a_1
X_15414_ _05646_ _05650_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__nand2_1
X_18202_ _08018_ _08415_ _08743_ vssd1 vssd1 vccd1 vccd1 _08747_ sky130_fd_sc_hd__or3_4
XFILLER_0_72_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12626_ _02716_ _02718_ vssd1 vssd1 vccd1 vccd1 _02719_ sky130_fd_sc_hd__xnor2_2
X_16394_ _06582_ _06665_ _06774_ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__or3b_4
X_18133_ _08669_ _08671_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__nand2_1
X_15345_ _05631_ _05641_ vssd1 vssd1 vccd1 vccd1 _05642_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12557_ _02608_ _02647_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18064_ _04887_ _06393_ _06394_ vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__nand3_1
X_11508_ _01585_ _01586_ _01593_ _01600_ vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15276_ _05452_ _05566_ vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _02521_ _02579_ _02570_ _02578_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__o211a_1
Xhold108 net113 vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17015_ _02837_ _02838_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__nor2_1
X_14227_ _04421_ _04353_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__nand2_1
Xhold119 _00027_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11439_ _03717_ _00197_ _01510_ _01531_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__a31o_1
X_14158_ _02999_ _01695_ _04346_ vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _00747_ _00748_ _00749_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__nor3_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _02986_ _05975_ _04269_ _04270_ vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__nand4_4
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ clknet_4_5_0_clk _09396_ vssd1 vssd1 vccd1 vccd1 salida\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _04337_ _06390_ _06389_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__a21o_1
X_18897_ clknet_4_11_0_clk _00051_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17848_ _08358_ _08359_ _08360_ vssd1 vssd1 vccd1 vccd1 _08361_ sky130_fd_sc_hd__or3_1
X_17779_ _08280_ _08285_ vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09966_ _09091_ _09123_ vssd1 vssd1 vccd1 vccd1 _09131_ sky130_fd_sc_hd__xnor2_2
X_09897_ _06213_ _06224_ _06202_ vssd1 vssd1 vccd1 vccd1 _08387_ sky130_fd_sc_hd__a21bo_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10810_ _00430_ _00899_ _00893_ _00898_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__o211a_1
X_11790_ _01540_ _01880_ _01879_ vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10741_ _07973_ cla_inst.in1\[22\] _08746_ _07984_ vssd1 vssd1 vccd1 vccd1 _00834_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13460_ _03577_ _03582_ _03079_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__mux2_1
X_10672_ _03782_ _03399_ _03476_ _03848_ vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12411_ _02436_ _02502_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__or2_1
X_13391_ _03491_ _03492_ _03506_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__nand3_2
XFILLER_0_152_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15130_ _05199_ _05077_ _05198_ _05302_ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__nor4_1
X_12342_ _02433_ _02434_ vssd1 vssd1 vccd1 vccd1 _02435_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ _03008_ _07515_ _05856_ _05878_ vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _02361_ _02364_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__and2b_1
X_14012_ _04174_ _04016_ _04185_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__and3_1
X_11224_ _00318_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__buf_4
X_18820_ _09324_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__buf_1
X_11155_ _00134_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__clkbuf_8
X_10106_ _00183_ _00181_ _00197_ _00173_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__a22o_1
X_18751_ _02533_ net65 _09251_ vssd1 vssd1 vccd1 vccd1 _09270_ sky130_fd_sc_hd__mux2_1
X_11086_ _01039_ _01048_ _01049_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__or3_4
X_15963_ _06282_ _06310_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or2_1
X_17702_ _08185_ _08201_ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__xor2_1
X_14914_ _05171_ _05172_ vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__nand2_1
X_10037_ _00129_ vssd1 vssd1 vccd1 vccd1 _00130_ sky130_fd_sc_hd__buf_6
X_18682_ net41 _09189_ _09218_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__o21a_1
X_15894_ _06156_ _06204_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__or2_1
X_17633_ _02848_ _08125_ _08127_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__a21o_2
X_14845_ _04077_ _04083_ _02978_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14776_ _09352_ _00460_ _05020_ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__and4_1
X_17564_ _08050_ _08051_ vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11988_ _01990_ _02000_ _02080_ vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _03857_ _03858_ _03874_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16515_ _06839_ _06840_ _06838_ vssd1 vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__a21oi_2
X_10939_ _03454_ _01031_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__and2_1
X_17495_ _07124_ _07511_ _07861_ _06581_ vssd1 vssd1 vccd1 vccd1 _07977_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13658_ _03797_ _03798_ _03799_ vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__nand3_2
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16446_ _06649_ _06834_ vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12609_ _02650_ net203 vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__xnor2_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16377_ _06529_ _06565_ _06759_ _06520_ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13589_ _03722_ _03723_ _03469_ _03516_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__o211a_1
XFILLER_0_81_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15328_ _03538_ _03121_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__nor2_2
XFILLER_0_124_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18116_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15259_ _05536_ _05547_ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__xor2_1
X_18047_ _08576_ _08577_ vssd1 vssd1 vccd1 vccd1 _08578_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09820_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07548_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09751_ _06743_ _06787_ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__nor2_1
X_18949_ clknet_4_5_0_clk _09408_ vssd1 vssd1 vccd1 vccd1 salida\[2\] sky130_fd_sc_hd__dfxtp_2
X_09682_ _05649_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _06646_ _06656_ vssd1 vssd1 vccd1 vccd1 _08951_ sky130_fd_sc_hd__and2_1
X_12960_ _03027_ _03052_ _01224_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21o_1
X_11911_ _04548_ _00197_ _02003_ vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__and3_1
X_12891_ _03629_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__buf_4
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _04723_ _04834_ _04860_ _04861_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__o211a_4
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _01837_ _01838_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__xnor2_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _04781_ _04786_ vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__xnor2_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11773_ _06482_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__clkbuf_8
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _03637_ _03638_ _03630_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__a21o_1
X_16300_ _06672_ _06674_ _06675_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__a21o_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10724_ _00801_ _00802_ _00810_ _00816_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17280_ _06561_ _07124_ _07314_ _07741_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__or4_4
X_14492_ _04705_ _04706_ _04709_ _04710_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__o211ai_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16231_ _01746_ _03029_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__or2_1
X_13443_ _03538_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10655_ _00745_ _00746_ _00537_ net124 vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_153_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16162_ _06522_ _06525_ _01113_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__a21oi_4
X_13374_ _03488_ _03489_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__xor2_2
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10586_ _09166_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ _05347_ _05387_ _05389_ vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__nor3_2
X_12325_ _02356_ _02365_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16093_ _03155_ _06451_ vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__and2_1
X_15044_ _02987_ _00495_ _05214_ vssd1 vssd1 vccd1 vccd1 _05314_ sky130_fd_sc_hd__and3_1
X_12256_ _02190_ _02348_ vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _06711_ _00460_ vssd1 vssd1 vccd1 vccd1 _01300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12187_ _02277_ _02278_ _02254_ _02264_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__o211a_1
X_18803_ _02994_ net51 _09301_ vssd1 vssd1 vccd1 vccd1 _09312_ sky130_fd_sc_hd__mux2_1
X_11138_ _01196_ _01229_ _01230_ _01143_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__o211a_1
X_16995_ _07430_ _07431_ vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__or2_1
X_18734_ _09245_ _09257_ vssd1 vssd1 vccd1 vccd1 _09258_ sky130_fd_sc_hd__and2_1
X_11069_ _01159_ _01160_ _01161_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__o21a_1
X_15946_ _03917_ _03908_ _02979_ vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__mux2_1
X_18665_ _09207_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__buf_1
X_15877_ _06193_ _06175_ _06218_ vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__o21ai_1
X_17616_ _08106_ _08107_ vssd1 vssd1 vccd1 vccd1 _08109_ sky130_fd_sc_hd__and2_1
X_14828_ _05078_ _04953_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__and2_1
X_18596_ net275 _09140_ _09154_ _09144_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ _02989_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__a21o_1
X_14759_ _00678_ _08452_ _01005_ _00679_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17478_ _06957_ _07035_ _07195_ _07608_ vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_698 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16429_ _06815_ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__buf_2
XFILLER_0_116_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09803_ _07352_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ cla_inst.in1\[20\] vssd1 vssd1 vccd1 vccd1 _06613_ sky130_fd_sc_hd__buf_6
X_09665_ _05834_ _05856_ _05475_ _05519_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09596_ _05006_ _05104_ vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__xnor2_2
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ _00349_ _00531_ _00529_ _00530_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10371_ _00447_ _00448_ _00449_ vssd1 vssd1 vccd1 vccd1 _00464_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12110_ _02198_ _02199_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__and3_1
X_13090_ _02370_ _03181_ _03022_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12041_ _02122_ _02132_ _02107_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__a211oi_2
X_15800_ _06065_ _06068_ _06133_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__nor3_1
X_13992_ _04146_ _04147_ _04164_ vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__o21ai_1
X_16780_ _06572_ _07106_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15731_ _06034_ _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__xor2_1
X_12943_ _08865_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__clkbuf_4
X_18450_ _08969_ _08978_ _09013_ vssd1 vssd1 vccd1 vccd1 _09014_ sky130_fd_sc_hd__or3_1
X_15662_ _05903_ _05905_ _05984_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__nor3_1
XANTENNA_120 _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ _02965_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__or2_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 _04132_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _07866_ _07873_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__xnor2_1
XANTENNA_142 _08180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _03793_ _09303_ _00498_ _03859_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__a22oi_1
X_11825_ _01877_ _01878_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__xor2_1
XANTENNA_153 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15593_ _05894_ _05825_ _05911_ vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__o21a_1
X_18381_ _06330_ _06405_ _06404_ vssd1 vssd1 vccd1 vccd1 _08940_ sky130_fd_sc_hd__a21o_1
XANTENNA_164 _08934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _01745_ _01139_ _04767_ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__a21o_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17332_ _07797_ _03930_ _07798_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__and3_2
X_11756_ _06008_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel _03388_
+ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _01849_ sky130_fd_sc_hd__and4_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10707_ _05943_ _05954_ _06127_ vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14475_ _04410_ _04692_ _04693_ _04551_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o2bb2a_1
X_17263_ _07018_ _07721_ _07723_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__o21a_1
X_11687_ net198 _01770_ _01721_ _01739_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ clknet_4_7_0_clk _09369_ vssd1 vssd1 vccd1 vccd1 salida\[55\] sky130_fd_sc_hd__dfxtp_1
X_16214_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__inv_2
X_13426_ _03081_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__clkbuf_4
X_10638_ _00725_ _00730_ vssd1 vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17194_ _00399_ _07311_ vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__and2_2
XFILLER_0_141_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16145_ _06507_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__buf_4
X_13357_ _03289_ _03268_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__and2b_1
X_10569_ _00659_ _00660_ _00601_ _00602_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a211oi_2
X_12308_ _08615_ _01357_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__nand2_1
X_16076_ _03169_ _06432_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__and2_1
X_13288_ _03230_ _03231_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__nand2_1
X_15027_ _05207_ _05176_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12239_ _07591_ _02205_ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__nand2_1
X_16978_ _07411_ _07412_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__or2b_1
Xinput4 i_wb_addr[11] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18717_ _09209_ _09243_ vssd1 vssd1 vccd1 vccd1 _09244_ sky130_fd_sc_hd__and2_1
X_15929_ _06195_ _06199_ vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__and2b_1
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09450_ cla_inst.in2\[19\] vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__buf_6
X_18648_ net60 _03083_ _09193_ vssd1 vssd1 vccd1 vccd1 _09194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18579_ salida\[10\] _09141_ _09142_ salida\[42\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09143_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09717_ _06406_ _06417_ vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09648_ _05671_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__buf_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _04810_ _04821_ _04831_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__a21o_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _01701_ _01700_ _01602_ _01585_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12590_ _02674_ _02681_ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _01630_ _01632_ _01631_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14260_ _04445_ _04446_ _04456_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__nor3_4
XFILLER_0_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11472_ _05453_ _05464_ _04154_ _00563_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__nand4_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _00164_ _03311_ vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10423_ _00509_ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__inv_4
XFILLER_0_33_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14191_ _04380_ _04381_ _04208_ _04212_ vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o211ai_4
X_13142_ _00620_ net136 _03237_ _03238_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__o211ai_2
X_10354_ _00438_ _00445_ _00446_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__nand3_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _03139_ _03148_ _03160_ _03163_ _03164_ _03081_ vssd1 vssd1 vccd1 vccd1 _03165_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_130_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17950_ _07608_ _07410_ _07511_ _07195_ vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__o22a_1
X_10285_ _09346_ _00274_ net338 _00377_ vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__a211oi_4
X_12024_ _02030_ _02029_ vssd1 vssd1 vccd1 vccd1 _02117_ sky130_fd_sc_hd__and2b_1
X_16901_ _07205_ _07227_ _07203_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__a21o_1
X_17881_ _08381_ _08396_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__xnor2_1
X_16832_ _07250_ _07252_ _07253_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16763_ _03094_ _06435_ vssd1 vssd1 vccd1 vccd1 _07180_ sky130_fd_sc_hd__nor2_1
X_13975_ _04144_ _04145_ _03963_ _03982_ vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18502_ _06414_ _07084_ _09058_ _09062_ _09069_ vssd1 vssd1 vccd1 vccd1 _09071_ sky130_fd_sc_hd__o311a_1
X_15714_ _06041_ _06042_ vssd1 vssd1 vccd1 vccd1 _06043_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ _00806_ _06591_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__or2_1
X_16694_ _02347_ _06871_ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18433_ _06836_ _08983_ _08987_ _08996_ vssd1 vssd1 vccd1 vccd1 _08997_ sky130_fd_sc_hd__o211a_1
X_15645_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__and2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _02948_ _02941_ _02933_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nor3_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _01811_ _01812_ _01899_ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a211o_1
X_18364_ _08873_ _08893_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__or3_1
X_15576_ _05830_ _05843_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__and2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _02879_ _02880_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__and2b_2
XFILLER_0_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17315_ _06750_ _07780_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__nand2_1
X_14527_ _04743_ _04749_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11739_ _01829_ _01830_ _01831_ vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18295_ _08845_ _08846_ vssd1 vssd1 vccd1 vccd1 _08847_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ _07590_ _07600_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _04672_ _04673_ _04529_ _04531_ vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ _03525_ _03526_ _03349_ _03365_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_141_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14389_ _04596_ _04597_ _04445_ net335 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17177_ _06875_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16128_ _00861_ _03140_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16059_ _06328_ _06412_ _06413_ _06248_ vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_20_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09502_ _04078_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__buf_6
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09433_ _03324_ _03206_ _03228_ _03292_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 _01225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_42 _02188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_64 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_75 _06693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_86 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_97 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10070_ cla_inst.in2\[20\] vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _02978_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__buf_4
X_10972_ _05584_ cla_inst.in1\[16\] ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel
+ _05562_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12711_ _02755_ _02785_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__nor2_1
X_13691_ _03697_ _03698_ _03712_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ _05631_ _05641_ _05639_ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__a21oi_1
X_12642_ _02689_ _02734_ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__and2_1
X_15361_ _05577_ _05580_ _05578_ vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_65_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ _02656_ _02665_ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17100_ _07536_ _07538_ _07545_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__or3_1
X_14312_ _04320_ _04322_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__nor2_1
X_11524_ _01615_ _01616_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__xnor2_2
X_15292_ _03000_ _03071_ _05583_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__nand3_1
X_18080_ _08592_ _08596_ _08613_ _06721_ _01136_ vssd1 vssd1 vccd1 vccd1 _09400_ sky130_fd_sc_hd__o32a_2
XFILLER_0_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14243_ _02059_ _08224_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__nand2_1
X_17031_ _06364_ _06545_ _07470_ _00593_ vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__a22o_1
X_11455_ _01546_ _01547_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ _07080_ _09303_ _00498_ _07058_ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14174_ _09352_ _01962_ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11386_ _01475_ _01476_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ _03213_ _03214_ _03220_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10337_ _00428_ _00270_ _00427_ _00429_ vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a211oi_4
X_18982_ clknet_4_0_0_clk _09377_ vssd1 vssd1 vccd1 vccd1 salida\[35\] sky130_fd_sc_hd__dfxtp_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _03147_ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__inv_2
X_17933_ _07751_ _07596_ _08453_ vssd1 vssd1 vccd1 vccd1 _08454_ sky130_fd_sc_hd__a21oi_1
X_10268_ _00357_ _00359_ _00360_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__a21bo_1
X_12007_ _06765_ _02099_ _02032_ _02033_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__o22a_1
X_17864_ _08277_ _08290_ _08275_ vssd1 vssd1 vccd1 vccd1 _08379_ sky130_fd_sc_hd__a21o_1
X_10199_ _08420_ _08463_ _08431_ vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16815_ _06665_ _07130_ vssd1 vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__nor2_1
X_17795_ _08302_ _08303_ vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16746_ _07158_ _07159_ _03195_ vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13958_ _03952_ _03958_ vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__or2_1
X_12909_ _02990_ _02995_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__or3_2
X_16677_ _03062_ _06724_ vssd1 vssd1 vccd1 vccd1 _07086_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13889_ _04050_ _04051_ _03834_ net321 vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__a211oi_1
X_18416_ _08971_ _08976_ vssd1 vssd1 vccd1 vccd1 _08978_ sky130_fd_sc_hd__nor2_4
X_15628_ _05876_ _05873_ _05874_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__o21ai_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18347_ _08901_ _08902_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__and2_1
X_15559_ _05873_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__or2b_1
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18278_ _03036_ _06148_ _06426_ _08825_ _08828_ vssd1 vssd1 vccd1 vccd1 _08829_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput40 i_wb_data[14] vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__buf_2
X_17229_ _04247_ _06914_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput51 i_wb_data[24] vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput62 i_wb_data[5] vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_2
XFILLER_0_71_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09982_ _07755_ vssd1 vssd1 vccd1 vccd1 _09248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11240_ _01330_ _01331_ _01313_ _01314_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11171_ _00193_ vssd1 vssd1 vccd1 vccd1 _01264_ sky130_fd_sc_hd__buf_4
XFILLER_0_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10122_ _00203_ _00214_ vssd1 vssd1 vccd1 vccd1 _00215_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14930_ _05188_ _05189_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__nand2_1
X_10053_ _00145_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__buf_4
X_14861_ _04975_ _04982_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__nand2_2
X_16600_ _06999_ _07001_ _03080_ vssd1 vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__mux2_1
X_13812_ _03790_ _03455_ vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__nand2_1
X_17580_ _07130_ _07126_ _07195_ _07608_ vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__or4_1
X_14792_ _00190_ _00192_ _05986_ _01223_ vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__and4_1
X_16531_ _06344_ _06346_ _06926_ vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a21oi_1
X_13743_ net119 _03889_ _03891_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__o21a_1
X_10955_ _01044_ _01047_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16462_ _03166_ _06431_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13674_ cla_inst.in2\[30\] cla_inst.in2\[29\] _03432_ _00205_ vssd1 vssd1 vccd1 vccd1
+ _03818_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ _00967_ _00977_ _00976_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ _08588_ _08742_ _08743_ _08417_ _08744_ vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__o221a_1
X_15413_ _05691_ _05690_ vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__or2b_1
XFILLER_0_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12625_ _02681_ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__or2_2
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16393_ _06583_ _06750_ _06775_ _06777_ vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _08614_ _08590_ _08668_ _06516_ vssd1 vssd1 vccd1 vccd1 _08671_ sky130_fd_sc_hd__o31a_1
X_15344_ _05639_ _05640_ vssd1 vssd1 vccd1 vccd1 _05641_ sky130_fd_sc_hd__nor2_1
X_12556_ _07788_ _00878_ _02607_ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11507_ _01594_ _01599_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__and2_1
X_18063_ _01997_ _08593_ _08595_ vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_108_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15275_ _05556_ _05565_ vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__xor2_1
X_12487_ _02570_ _02578_ _02521_ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a211oi_2
Xhold109 _00012_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _03195_ _07451_ _07452_ vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__or3b_2
X_14226_ _00592_ _04336_ vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__and2_1
X_11438_ _04078_ _01151_ _01031_ _09179_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14157_ _04344_ _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__xnor2_1
X_11369_ _01460_ _01461_ vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__or2_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__buf_6
X_14088_ _03651_ _03662_ _00308_ _08757_ vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__nand4_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ clknet_4_7_0_clk _09395_ vssd1 vssd1 vccd1 vccd1 salida\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _06425_ _06444_ _08435_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__or3_1
X_13039_ _00494_ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__or2_1
X_18896_ clknet_4_11_0_clk _00050_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_17847_ _07143_ _07706_ _08260_ _06961_ vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__o22a_1
X_17778_ _08283_ _08284_ vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16729_ _07140_ _07141_ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09965_ _09101_ _09112_ vssd1 vssd1 vccd1 vccd1 _09123_ sky130_fd_sc_hd__and2b_1
X_09896_ _08333_ _08354_ _08344_ vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__a21o_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10740_ _07036_ _07069_ cla_inst.in1\[22\] _08746_ vssd1 vssd1 vccd1 vccd1 _00833_
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ _03848_ _03782_ _03399_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12410_ _02436_ _02502_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ _03491_ _03492_ _03506_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__a21o_2
XFILLER_0_105_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12341_ _02418_ _02432_ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15060_ _03006_ _01866_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12272_ _02361_ _02364_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__xnor2_1
X_14011_ _04174_ _04016_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11223_ _00862_ _01107_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__and2_1
X_11154_ _01240_ _01246_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__xnor2_4
X_10105_ _00195_ _00175_ _00181_ _00197_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__nand4_1
X_18750_ _09269_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__buf_1
X_11085_ _01166_ _01176_ _01177_ vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__nor3_1
X_15962_ _06258_ _06284_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__nor2_1
X_17701_ _08187_ _08200_ vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__xnor2_1
X_14913_ _02999_ _03055_ _05169_ vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__a21o_1
X_10036_ ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00129_ sky130_fd_sc_hd__buf_6
X_18681_ _02044_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09218_ sky130_fd_sc_hd__a21oi_1
X_15893_ _06171_ _06214_ _06216_ vssd1 vssd1 vccd1 vccd1 _06236_ sky130_fd_sc_hd__a21oi_1
X_17632_ _02848_ _08125_ _03201_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__o21ai_1
X_14844_ _02974_ _05095_ vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17563_ _06766_ _07706_ vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__nor2_1
X_14775_ _03322_ _03321_ _05486_ _05878_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__nand4_1
XFILLER_0_98_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11987_ _02053_ _02078_ _02079_ vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16514_ _08865_ _06509_ _00223_ vssd1 vssd1 vccd1 vccd1 _06909_ sky130_fd_sc_hd__a21boi_1
X_13726_ _03857_ _03858_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__a21oi_1
X_10938_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _01031_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17494_ _07841_ _07848_ vssd1 vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16445_ _06775_ _06779_ _06832_ vssd1 vssd1 vccd1 vccd1 _06834_ sky130_fd_sc_hd__a21o_1
X_13657_ _03632_ _03634_ _03633_ vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a21bo_1
X_10869_ _03465_ _00171_ _00771_ _00773_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12608_ _02662_ _02695_ _02700_ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__or3b_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _04384_ _03281_ vssd1 vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__and2_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _03469_ _03516_ _03722_ _03723_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18115_ _08650_ _08651_ vssd1 vssd1 vccd1 vccd1 _08652_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15327_ _05619_ _05620_ _05622_ vssd1 vssd1 vccd1 vccd1 _09363_ sky130_fd_sc_hd__a21bo_1
X_12539_ _02592_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _08482_ _08531_ _08575_ vssd1 vssd1 vccd1 vccd1 _08577_ sky130_fd_sc_hd__and3_1
X_15258_ _05545_ _05546_ vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14209_ _03742_ _04402_ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15189_ _05463_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _06754_ _06700_ _06765_ _06776_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__o2bb2a_1
X_18948_ clknet_4_5_0_clk _09397_ vssd1 vssd1 vccd1 vccd1 salida\[1\] sky130_fd_sc_hd__dfxtp_2
X_09681_ _06029_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__buf_4
X_18879_ clknet_4_15_0_clk net247 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ _08692_ _08702_ _08919_ vssd1 vssd1 vccd1 vccd1 _08941_ sky130_fd_sc_hd__nand3_2
X_09879_ _07700_ _08158_ _08180_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__and3_1
X_11910_ _02001_ _02002_ vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12890_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__clkbuf_4
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _01908_ _01912_ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__or2b_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560_ _04784_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__xnor2_1
X_11772_ _01675_ _01864_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__and2_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13511_ _03630_ _03637_ _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__nand3_1
X_10723_ _00811_ _00815_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__and2_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _01521_ _07156_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16230_ _01746_ _06595_ _06596_ _06599_ vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o2bb2a_1
X_10654_ _00537_ _00600_ _00745_ _00746_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__o211a_2
X_13442_ _02979_ _03562_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13373_ _01873_ _03107_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__nand2_1
X_16161_ _06051_ _05682_ _07047_ _06524_ vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__or4_4
XFILLER_0_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10585_ _09172_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__buf_2
XFILLER_0_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15112_ _05260_ _05283_ _05386_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12324_ _02414_ _02415_ vssd1 vssd1 vccd1 vccd1 _02417_ sky130_fd_sc_hd__xor2_1
XFILLER_0_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16092_ _03073_ _06408_ _06449_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15043_ _05210_ _05218_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ _08615_ _01746_ _01357_ _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__a22o_1
X_11206_ _01297_ _01298_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12186_ _02254_ _02264_ _02277_ _02278_ vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__a211oi_2
X_11137_ _01138_ _01140_ _01141_ _01135_ _01134_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__a32o_1
X_18802_ _09310_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__clkbuf_1
X_16994_ _07427_ _07429_ _07407_ vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__a21oi_1
X_18733_ _03077_ net57 _09251_ vssd1 vssd1 vccd1 vccd1 _09257_ sky130_fd_sc_hd__mux2_1
X_11068_ _03509_ _00871_ _07581_ _03345_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__a22o_1
X_15945_ _03911_ _03926_ _03912_ vssd1 vssd1 vccd1 vccd1 _06292_ sky130_fd_sc_hd__mux2_1
X_10019_ _00109_ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__clkbuf_4
X_18664_ _09176_ _09206_ vssd1 vssd1 vccd1 vccd1 _09207_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15876_ _06216_ _06217_ vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__nor2_1
X_17615_ _08106_ _08107_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14827_ _04942_ _04945_ vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18595_ salida\[17\] _09141_ _09142_ salida\[49\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17546_ _03693_ _06441_ _08032_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__o21a_1
X_14758_ _00679_ _00678_ _04591_ _01005_ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _03854_ _03855_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17477_ _07130_ _07195_ _07608_ _07042_ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__o22a_1
X_14689_ _04924_ _04925_ _04794_ _04796_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ _06811_ _06814_ _00181_ vssd1 vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__or3b_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16359_ _00881_ _03094_ _00167_ _03101_ _06477_ _03161_ vssd1 vssd1 vccd1 vccd1 _06740_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18029_ _08556_ _08557_ vssd1 vssd1 vccd1 vccd1 _08558_ sky130_fd_sc_hd__and2_1
X_09802_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07352_ sky130_fd_sc_hd__buf_4
X_09733_ _05399_ _06591_ cla_inst.in1\[20\] net233 vssd1 vssd1 vccd1 vccd1 _06602_
+ sky130_fd_sc_hd__and4_1
X_09664_ _05845_ vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__buf_4
X_09595_ _05061_ _05093_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__xnor2_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _00458_ _00462_ vssd1 vssd1 vccd1 vccd1 _00463_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12040_ _02050_ _02106_ _02105_ _02090_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_130_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13991_ _04148_ _04163_ vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__xnor2_1
X_15730_ _06058_ _06059_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__nand2_1
X_12942_ _02979_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__or2_4
XFILLER_0_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15661_ _05903_ _05905_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__o21a_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ _03239_ _03217_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__or2_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 _02476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_132 _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _07871_ _07872_ vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__xnor2_1
X_14612_ _04839_ _04840_ _04835_ _04836_ vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__a211o_1
XANTENNA_143 _08180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _01913_ _01916_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__and2b_1
X_18380_ _03120_ _06229_ _08938_ vssd1 vssd1 vccd1 vccd1 _08939_ sky130_fd_sc_hd__o21a_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _05908_ _05909_ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__xnor2_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 _09380_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17331_ _02589_ _02844_ vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__nand2_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14543_ _01745_ _01139_ _04767_ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__nand3_2
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _07363_ _01575_ _01846_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__a31o_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10706_ _00798_ _00791_ _00784_ vssd1 vssd1 vccd1 vccd1 _00799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17262_ _06969_ _07394_ _07396_ _06891_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__a22o_1
X_14474_ _04399_ _04400_ _04549_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11686_ _01748_ _01778_ vssd1 vssd1 vccd1 vccd1 _01779_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19001_ clknet_4_7_0_clk _09368_ vssd1 vssd1 vccd1 vccd1 salida\[54\] sky130_fd_sc_hd__dfxtp_1
X_16213_ _06561_ _06563_ _06572_ _06581_ vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__or4_2
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13425_ _03164_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10637_ _00728_ _00729_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17193_ _07645_ _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16144_ _03239_ _06418_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__nor2_1
X_10568_ _00601_ _00602_ _00659_ _00660_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__o211a_2
X_13356_ _03467_ _03468_ net131 _03373_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ _02395_ _02399_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__or2_1
X_16075_ _03086_ _01264_ _06431_ vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__and3_1
X_13287_ _03390_ _03391_ _03392_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__a21oi_1
X_10499_ _00591_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _05292_ _05294_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__xor2_2
X_12238_ _08724_ _00132_ _02206_ _02207_ vssd1 vssd1 vccd1 vccd1 _02331_ sky130_fd_sc_hd__a22oi_2
X_12169_ _00846_ _00557_ _02257_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__a21oi_2
X_16977_ net237 _06951_ _07035_ _07410_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__or4_1
Xinput5 i_wb_addr[12] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18716_ net56 _03073_ _09182_ vssd1 vssd1 vccd1 vccd1 _09243_ sky130_fd_sc_hd__mux2_1
X_15928_ _06237_ _06208_ _06240_ vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__a21o_1
X_18647_ _09182_ vssd1 vssd1 vccd1 vccd1 _09193_ sky130_fd_sc_hd__clkbuf_4
X_15859_ _03007_ _03149_ _06198_ vssd1 vssd1 vccd1 vccd1 _06199_ sky130_fd_sc_hd__and3_1
X_18578_ _09117_ vssd1 vssd1 vccd1 vccd1 _09142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17529_ _07931_ _07932_ _08013_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09716_ _04362_ _05028_ _04569_ _04635_ vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05671_ sky130_fd_sc_hd__buf_4
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _04853_ _04908_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__xnor2_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11540_ _01630_ _01631_ _01632_ vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nand3_2
XFILLER_0_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _01525_ _01540_ _01562_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__a211o_2
XFILLER_0_151_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13210_ _02124_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__buf_4
X_10422_ _00514_ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _04208_ _04212_ _04380_ _04381_ vssd1 vssd1 vccd1 vccd1 _04382_ sky130_fd_sc_hd__a211o_2
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10353_ _00435_ _00436_ _00437_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__a21o_1
X_13141_ _03224_ _03225_ _03236_ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _03062_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__clkbuf_4
X_10284_ _00372_ _00373_ _00376_ _00336_ vssd1 vssd1 vccd1 vccd1 _00377_ sky130_fd_sc_hd__o2bb2a_1
X_12023_ _00832_ _03815_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__nand2_1
X_16900_ _07300_ _07327_ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__xnor2_1
X_17880_ _08394_ _08395_ vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__nor2_1
X_16831_ _07250_ _07252_ _06559_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__a21oi_1
X_16762_ _03094_ _06435_ vssd1 vssd1 vccd1 vccd1 _07179_ sky130_fd_sc_hd__and2_1
X_13974_ _03963_ _03982_ _04144_ _04145_ vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__a211oi_2
X_18501_ _06426_ _06452_ _09063_ _09068_ vssd1 vssd1 vccd1 vccd1 _09069_ sky130_fd_sc_hd__o31a_1
X_15713_ _01359_ _04125_ _06038_ _06039_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__a22oi_1
X_12925_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel _06008_ vssd1
+ vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__or2_1
X_16693_ _07019_ _07046_ vssd1 vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18432_ _06410_ _07084_ _08988_ _08990_ _08994_ vssd1 vssd1 vccd1 vccd1 _08996_ sky130_fd_sc_hd__o311a_1
X_15644_ _05958_ _05965_ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__nand2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _02941_ _02933_ _02948_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11807_ _01897_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__inv_2
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _08917_ _08920_ vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__xnor2_1
X_15575_ _05890_ _05891_ vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__and2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _02863_ _02872_ _02878_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _02259_ _06814_ vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__nor2_4
XFILLER_0_139_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14526_ _04747_ _04748_ vssd1 vssd1 vccd1 vccd1 _04749_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _05279_ _05355_ _03607_ _00217_ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__nand4_2
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18294_ _03107_ _07390_ vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17245_ _07603_ _07615_ vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__nor2_1
X_14457_ _04529_ _04531_ _04672_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_114_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11669_ _01217_ _01219_ _01227_ vssd1 vssd1 vccd1 vccd1 _01762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13408_ _03349_ _03365_ _03525_ _03526_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17176_ _07627_ _07628_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__or2_1
X_14388_ _04445_ net335 _04596_ _04597_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_40_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ _03152_ _06485_ _06486_ _06487_ vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13339_ _03279_ _03285_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16058_ _03011_ _03155_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ _05263_ _05171_ _05275_ vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09501_ cla_inst.in2\[16\] vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09432_ _03313_ vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_10 _00516_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_21 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 _01266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 _02200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 _03618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_65 _04537_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_76 _06799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_87 _08820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_98 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _05562_ _05584_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel vssd1
+ vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__and3_1
X_12710_ _02794_ _02802_ vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13690_ _03832_ _03833_ _03649_ _03751_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_57_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12641_ _02691_ _02711_ _02726_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15360_ _05656_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__xnor2_1
X_12572_ _02658_ _02663_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14311_ _01356_ _01962_ _04364_ _04363_ vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11523_ _01541_ _01543_ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15291_ _05581_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17030_ _08615_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__a21o_1
X_14242_ _04436_ _04437_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11454_ _01543_ _01545_ _01544_ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10405_ cla_inst.in1\[28\] vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__buf_2
XFILLER_0_123_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14173_ _04361_ _04363_ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__nor2_1
X_11385_ _01477_ _00879_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ _03218_ _03219_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__xor2_2
X_10336_ _00424_ _00426_ _09348_ _00273_ vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__o211a_1
X_18981_ clknet_4_1_0_clk _09366_ vssd1 vssd1 vccd1 vccd1 salida\[34\] sky130_fd_sc_hd__dfxtp_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _07504_ _00127_ _07559_ _00358_ vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__a22o_1
X_13055_ _03141_ _03146_ _03049_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__mux2_1
X_17932_ _07218_ _07486_ vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__nor2_1
X_12006_ _00563_ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__inv_4
X_17863_ _08366_ _08377_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__xor2_1
X_10198_ _00288_ _00289_ _00290_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__and3_2
XFILLER_0_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814_ _07233_ _07234_ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__xor2_1
X_17794_ _07630_ _07741_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__nor2_1
X_16745_ _07158_ _07159_ vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__nor2_1
X_13957_ _03974_ _03975_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__a21o_1
X_12908_ _02997_ _02998_ _03000_ _00591_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__or4_1
X_16676_ _06343_ _06342_ _06997_ _07084_ vssd1 vssd1 vccd1 vccd1 _07085_ sky130_fd_sc_hd__a31o_1
X_13888_ _03834_ net321 _04050_ _04051_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15627_ _05948_ _05875_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__nor2_1
X_18415_ _08971_ _08976_ vssd1 vssd1 vccd1 vccd1 _08977_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12839_ _02930_ _02931_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__xnor2_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18346_ _04537_ _07743_ _08900_ vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_139_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15558_ _05870_ _05871_ _05872_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__o21ai_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14509_ _04576_ _04577_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__o21ai_4
X_18277_ _07269_ _08141_ _08827_ _06721_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15489_ _02973_ _03564_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17228_ _06639_ _06627_ _02981_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__mux2_1
Xinput30 i_wb_addr[6] vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 i_wb_data[15] vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput52 i_wb_data[25] vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__buf_1
XFILLER_0_71_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput63 i_wb_data[6] vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_2
XFILLER_0_52_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17159_ _06764_ _07018_ _07194_ _07608_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09981_ _09226_ _09232_ vssd1 vssd1 vccd1 vccd1 _09240_ sky130_fd_sc_hd__or2_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11170_ _01261_ _01262_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ _00213_ vssd1 vssd1 vccd1 vccd1 _00214_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ ApproximateM_inst.lob_16.lob1.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00145_ sky130_fd_sc_hd__clkbuf_4
X_14860_ _05109_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__xnor2_1
X_13811_ _03774_ net171 _03966_ vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_98_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14791_ _02996_ _01139_ _01223_ _02993_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16530_ _06338_ _06348_ _06349_ vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13742_ net119 _03889_ _03891_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__nor3_1
XFILLER_0_98_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10954_ _06460_ _04067_ _01045_ _01046_ vssd1 vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _03166_ _03083_ _06430_ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__and3_1
X_13673_ cla_inst.in2\[31\] _00172_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__nand2_1
X_10885_ _00967_ _00976_ _00977_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18200_ _08582_ _08614_ _08667_ vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_39_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15412_ _03548_ _05623_ _05625_ _03125_ _05714_ vssd1 vssd1 vccd1 vccd1 _09364_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12624_ _02675_ _02680_ _02679_ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__a21oi_1
X_16392_ _06659_ _06668_ _06774_ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18131_ _08614_ _08590_ _08668_ vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__o21ai_1
X_15343_ _05636_ _05637_ _05632_ vssd1 vssd1 vccd1 vccd1 _05640_ sky130_fd_sc_hd__a21oi_1
X_12555_ _02608_ _02647_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11506_ _01595_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__xor2_2
X_18062_ _01997_ _08593_ _03930_ vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15274_ _05563_ _05564_ vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__nor2_1
X_12486_ _02515_ _02520_ _02519_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__o21a_1
XFILLER_0_123_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17013_ _07345_ _07349_ _07449_ vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__or3_1
X_14225_ _04390_ _04391_ _04392_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__or3_4
X_11437_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _03618_ _01527_
+ _01528_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14156_ _04175_ _04179_ _04177_ vssd1 vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__o21ba_1
X_11368_ _01458_ _01459_ _01455_ _01456_ vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__o211a_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13107_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _00401_ _00402_ _00411_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__o21a_1
X_14087_ _03662_ _05704_ _08757_ _03629_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__a22o_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ clknet_4_7_0_clk _09394_ vssd1 vssd1 vccd1 vccd1 salida\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _01382_ _01389_ _01390_ _01391_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__nand4_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _03041_ _06443_ _04336_ vssd1 vssd1 vccd1 vccd1 _08435_ sky130_fd_sc_hd__a21oi_1
X_13038_ _03127_ _03129_ _03048_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__mux2_1
X_18895_ clknet_4_11_0_clk _00049_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17846_ _07143_ _08262_ vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14989_ _05248_ _05253_ vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__xnor2_1
X_17777_ _07109_ _07649_ vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16728_ _07040_ _07043_ _07037_ vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ _07063_ _07065_ vssd1 vssd1 vccd1 vccd1 _07066_ sky130_fd_sc_hd__and2b_1
XFILLER_0_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18329_ _06403_ _06546_ _08883_ _03143_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_115_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09964_ _07080_ _07374_ _07406_ _07047_ vssd1 vssd1 vccd1 vccd1 _09112_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09895_ _08333_ _08344_ _08354_ vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__nand3_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ _04296_ _04285_ _04187_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12340_ _02418_ _02432_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ _02362_ _02363_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__xnor2_1
X_14010_ _04183_ _04184_ vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__nand2_1
X_11222_ _00862_ _01107_ vssd1 vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11153_ _01243_ _01245_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__nor2_2
X_10104_ _00196_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__buf_4
X_11084_ _01149_ _01150_ _01165_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__a21oi_2
X_15961_ _06306_ _06307_ vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__and2_1
X_17700_ _08198_ _08199_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__nor2_1
X_14912_ _02999_ _03055_ _05169_ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__nand3_1
X_10035_ _00125_ _00127_ _09188_ _00109_ vssd1 vssd1 vccd1 vccd1 _00128_ sky130_fd_sc_hd__a22o_1
X_18680_ net40 _09189_ _09217_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__o21a_1
X_15892_ _06190_ _06225_ _06231_ _06184_ _06233_ vssd1 vssd1 vccd1 vccd1 _06235_ sky130_fd_sc_hd__o221a_1
X_14843_ _03912_ _04082_ _05094_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__o21ai_1
X_17631_ _02846_ _02847_ _02465_ vssd1 vssd1 vccd1 vccd1 _08125_ sky130_fd_sc_hd__a21bo_1
X_17562_ _08045_ _08046_ _08048_ vssd1 vssd1 vccd1 vccd1 _08050_ sky130_fd_sc_hd__a21o_1
X_14774_ _09350_ _05486_ _05878_ _00112_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__a22o_1
X_11986_ _02073_ _02077_ _01984_ _02054_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__o211a_1
X_16513_ _03086_ _06509_ _08865_ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__and3b_1
X_13725_ _03861_ _03873_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10937_ _00936_ _00935_ _00934_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17493_ _07843_ _07847_ vssd1 vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16444_ _06775_ _06779_ _06832_ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__and3_1
X_13656_ _08713_ _09303_ _03795_ _03796_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__nand4_2
XFILLER_0_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ _00958_ _00960_ vssd1 vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12607_ _02693_ _02696_ _02699_ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__nor3b_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _06531_ _06533_ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _03674_ _03675_ _03720_ _03721_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ _00270_ _00271_ _00272_ _09348_ vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__a22o_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18114_ _08548_ _08562_ _08546_ vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__a21o_1
X_15326_ _03165_ _05307_ _05621_ _03039_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__o22a_1
X_12538_ _02628_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045_ _08482_ _08531_ _08575_ vssd1 vssd1 vccd1 vccd1 _08576_ sky130_fd_sc_hd__a21oi_1
X_15257_ _05537_ _05544_ vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__nand2_1
X_12469_ _02561_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__inv_2
XFILLER_0_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14208_ _03741_ _03902_ _04068_ _04236_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__nor4_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15188_ _05465_ _05470_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__xnor2_1
X_14139_ _04322_ _04324_ _04319_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18947_ clknet_4_3_0_clk _09386_ vssd1 vssd1 vccd1 vccd1 salida\[0\] sky130_fd_sc_hd__dfxtp_2
X_09680_ _06019_ vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__clkbuf_4
X_18878_ clknet_4_15_0_clk net248 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__dfxtp_1
X_17829_ _06734_ _08243_ _08340_ _06461_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09947_ _08692_ _08702_ _08919_ vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__a21o_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _07799_ _08169_ vssd1 vssd1 vccd1 vccd1 _08180_ sky130_fd_sc_hd__and2_2
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _01905_ _01907_ vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__or2_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11771_ _01106_ _01862_ _01863_ vssd1 vssd1 vccd1 vccd1 _01864_ sky130_fd_sc_hd__or3b_4
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13510_ _03635_ _03636_ _03631_ _03419_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__a211o_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _08082_ _00814_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__nor2_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14490_ _02986_ _07156_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__nand4_2
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13441_ _03560_ _03561_ _03098_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ _00696_ _00697_ _00743_ _00744_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16160_ _03003_ _03004_ _03018_ _06523_ vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__or4_4
XFILLER_0_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13372_ _03484_ _03486_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _00663_ _00664_ _00675_ vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15111_ _05260_ _05283_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12323_ _02414_ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__or2_1
X_16091_ _03068_ _06448_ vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15042_ _05216_ _05217_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__nand2_1
X_12254_ _02188_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11205_ _08713_ _08452_ _01002_ _01001_ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12185_ _02275_ _02276_ _02224_ vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__a21oi_1
X_18801_ _09298_ _09309_ vssd1 vssd1 vccd1 vccd1 _09310_ sky130_fd_sc_hd__and2_1
X_11136_ _01187_ _01192_ _01196_ _01197_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__a211oi_2
X_16993_ _07407_ _07427_ _07429_ vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__and3_1
X_18732_ _09255_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__clkbuf_1
X_11067_ _03345_ net242 _01031_ _07581_ vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__and4_1
X_15944_ _02976_ _04241_ _03918_ _03036_ vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__a31o_1
X_10018_ _00110_ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__inv_2
X_15875_ _06203_ _06215_ vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__nor2_1
X_18663_ net65 _03094_ _09193_ vssd1 vssd1 vccd1 vccd1 _09206_ sky130_fd_sc_hd__mux2_1
X_17614_ _06750_ _07859_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14826_ _05074_ _05076_ vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__nand2_2
X_18594_ net289 _09140_ _09153_ _09144_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14757_ _03006_ _02124_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__nand2_1
X_17545_ _03693_ _06441_ _06426_ vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__a21oi_1
X_11969_ _01913_ _01916_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13708_ _00163_ _01866_ _03853_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17476_ _06891_ _07390_ _07836_ _07834_ vssd1 vssd1 vccd1 vccd1 _07956_ sky130_fd_sc_hd__a31o_1
X_14688_ _04794_ _04796_ _04924_ _04925_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13639_ _04690_ _07406_ _03776_ _03777_ vssd1 vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__o2bb2a_1
X_16427_ _06813_ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16358_ _06736_ _06738_ _03098_ vssd1 vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15309_ _05499_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16289_ _06660_ _06663_ _00494_ vssd1 vssd1 vccd1 vccd1 _06664_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18028_ _08455_ _08549_ _08555_ vssd1 vssd1 vccd1 vccd1 _08557_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09801_ _05627_ _05725_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__or2_1
X_09732_ ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _06591_ sky130_fd_sc_hd__buf_4
X_09663_ _05322_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__clkbuf_8
X_09594_ _05072_ _05083_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__and2b_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13990_ _04161_ _04162_ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12941_ _02981_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15660_ _05890_ _05983_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__xnor2_1
X_12872_ op_code\[2\] op_code\[3\] vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__nand2b_2
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 _09374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_111 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _04835_ _04836_ _04839_ _04840_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__o211ai_2
XANTENNA_122 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 _04191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _01815_ _01915_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _05811_ _05821_ _05819_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__a21oi_1
XANTENNA_144 _08615_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_155 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 net172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _02589_ _02844_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__or2_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _04764_ _04765_ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__xor2_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11754_ _01082_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _01847_ sky130_fd_sc_hd__and4_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04722_ _00780_ _00782_ vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__a21o_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _06880_ _07194_ _07290_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__or3_2
X_14473_ _04551_ _04401_ net215 vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__and3b_1
XFILLER_0_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11685_ _01776_ _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nor2_1
X_16212_ _06579_ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19000_ clknet_4_4_0_clk _09367_ vssd1 vssd1 vccd1 vccd1 salida\[53\] sky130_fd_sc_hd__dfxtp_1
X_13424_ _03065_ _03075_ _02983_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__mux2_1
X_10636_ _00106_ _00212_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17192_ _07643_ _07644_ vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16143_ _02976_ _06505_ vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_141_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13355_ net131 _03373_ _03467_ _03468_ vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__o211ai_4
X_10567_ _00634_ _00635_ _00657_ _00658_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__nand4_4
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12306_ _02392_ _02394_ _02393_ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__o21a_1
X_16074_ _01248_ _06430_ vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__and2_1
X_13286_ _03390_ _03391_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__and3_2
X_10498_ _00164_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__buf_4
X_15025_ _05059_ _05186_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a21o_1
X_12237_ _02326_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__or2_1
X_12168_ _02258_ _02260_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__and2_1
X_11119_ _05573_ _05595_ _04395_ _03739_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__and4_1
X_12099_ _02191_ _02085_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__xnor2_1
X_16976_ _06951_ _07035_ _07410_ net237 vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__o22a_1
X_18715_ _09242_ vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__clkbuf_1
Xinput6 i_wb_addr[13] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ _06270_ _06271_ vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__nand2_1
X_18646_ net57 _09189_ _09192_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__o21a_1
X_15858_ _06196_ _06197_ vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14809_ _04920_ _04922_ vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18577_ _09113_ vssd1 vssd1 vccd1 vccd1 _09141_ sky130_fd_sc_hd__clkbuf_4
X_15789_ _06097_ _06123_ vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17528_ _08011_ _08012_ vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17459_ _06657_ _07708_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09715_ _04340_ _04362_ _05028_ cla_inst.in1\[16\] vssd1 vssd1 vccd1 vccd1 _06406_
+ sky130_fd_sc_hd__and4_1
X_09646_ _05649_ _05606_ _05617_ _05573_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__a22o_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _04875_ _04897_ vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__nor2_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11470_ _01550_ _01561_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ ApproximateM_inst.lob_16.lob2.mux.sel vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_61_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13140_ _03224_ _03225_ _03236_ vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10352_ _00442_ _00444_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13071_ _03161_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__nand2_1
X_10283_ _00333_ _00335_ _08681_ _09005_ vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__o211a_1
X_12022_ _02112_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__nor2_1
X_16830_ _07158_ _07159_ _07251_ vssd1 vssd1 vccd1 vccd1 _07252_ sky130_fd_sc_hd__a21oi_2
X_13973_ _04123_ _04124_ _04142_ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__nor3_4
XFILLER_0_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16761_ _06355_ _06790_ _07176_ _03094_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__a22o_1
X_18500_ _03916_ _06999_ _08141_ _09066_ _09067_ vssd1 vssd1 vccd1 vccd1 _09068_ sky130_fd_sc_hd__o311a_1
X_15712_ _01359_ _04125_ _06038_ _06039_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__and4_1
X_12924_ _03007_ _03011_ _03013_ _03016_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__or4_2
X_16692_ _07072_ _07075_ _07101_ _06723_ _02214_ vssd1 vssd1 vccd1 vccd1 _09415_ sky130_fd_sc_hd__o32a_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18431_ _03119_ _06266_ _07579_ _08141_ _08993_ vssd1 vssd1 vccd1 vccd1 _08994_ sky130_fd_sc_hd__o221a_1
X_15643_ _05958_ _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__or2_1
X_12855_ _02942_ _02947_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__xnor2_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11806_ _01876_ _01897_ _01898_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__and3_1
X_15574_ _05882_ _05889_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__nand2_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _08868_ _08918_ vssd1 vssd1 vccd1 vccd1 _08920_ sky130_fd_sc_hd__nor2_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _02863_ _02872_ _02878_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__and3_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _07537_ _01962_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17313_ _07776_ _07778_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__and2b_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _06591_ _03607_ _00774_ _00806_ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18293_ _04668_ _04679_ _07743_ vssd1 vssd1 vccd1 vccd1 _08845_ sky130_fd_sc_hd__nor3_1
X_14456_ _04670_ _04671_ _04484_ vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__o21ai_1
X_17244_ _07589_ _07601_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11668_ _01201_ _01759_ _01757_ _01758_ vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_142_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13407_ _03523_ _03524_ _03367_ _03369_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10619_ _00700_ _00701_ _00711_ vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17175_ _07622_ _07625_ _07626_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__a21oi_1
X_14387_ _04584_ _04585_ _04595_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__or3_4
XFILLER_0_4_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ _05246_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__inv_6
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16126_ _02728_ _03002_ _03021_ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__or3_2
X_13338_ _03280_ _03284_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__nand2_1
X_16057_ _06024_ _06410_ _06411_ _06328_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13269_ _00620_ net136 _03237_ _03238_ vssd1 vssd1 vccd1 vccd1 _03374_ sky130_fd_sc_hd__o211a_2
XFILLER_0_121_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15008_ _05273_ _05274_ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16959_ _07388_ _07391_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__nand2_1
X_09500_ _04056_ vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__buf_6
XFILLER_0_79_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09431_ sel_op\[0\] vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__clkbuf_4
X_18629_ salida\[31\] _09113_ _09117_ salida\[63\] _09127_ vssd1 vssd1 vccd1 vccd1
+ _09177_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_11 _00644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 _01266_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 _02533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_55 _03760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_66 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_88 _08820_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_99 _08934_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ _05671_ _05039_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__nand2_1
X_09629_ _05453_ _05464_ _05388_ _05050_ vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__nand4_2
X_12640_ _02700_ _02731_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__or3_4
XFILLER_0_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12571_ _02622_ _02659_ _02662_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__or3b_1
XFILLER_0_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14310_ _04359_ _04367_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__and2_1
XFILLER_0_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _01613_ _01614_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__and2b_1
X_15290_ _05481_ _05484_ _05482_ vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ _03859_ _04132_ _07015_ _07112_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__and4_1
X_11453_ _01543_ _01544_ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ _05736_ _07025_ _00317_ _00319_ _00318_ vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a32o_1
X_14172_ _00148_ _00149_ _08409_ _03750_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and4_1
X_11384_ _00204_ _00878_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13123_ _04001_ _05257_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__nand2_1
X_10335_ _00268_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__inv_2
X_18980_ clknet_4_0_0_clk _09355_ vssd1 vssd1 vccd1 vccd1 salida\[33\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _03145_ vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__inv_2
X_17931_ _08358_ _08359_ _08360_ _08356_ vssd1 vssd1 vccd1 vccd1 _08451_ sky130_fd_sc_hd__nor4b_1
X_10266_ _00358_ _07504_ _00127_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__and3_1
X_12005_ _02092_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__xnor2_1
X_17862_ _08367_ _08375_ vssd1 vssd1 vccd1 vccd1 _08377_ sky130_fd_sc_hd__xnor2_1
X_10197_ _08474_ _08485_ _08398_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__a21bo_1
X_16813_ _07127_ _07131_ _07128_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__o21ai_2
X_17793_ _08299_ _08301_ vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16744_ _07067_ _07070_ _07066_ vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__a21o_1
X_13956_ _03790_ _04125_ _03976_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12907_ _02999_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__clkbuf_4
X_13887_ _04004_ _04005_ _04048_ _04049_ vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__o22ai_2
X_16675_ _06598_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18414_ _08749_ _08810_ _08972_ _08975_ vssd1 vssd1 vccd1 vccd1 _08976_ sky130_fd_sc_hd__o31a_1
X_12838_ _02909_ _02911_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__or2b_2
X_15626_ _05786_ _05788_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__xnor2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18345_ _04537_ _07743_ _08900_ vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__or3_1
X_15557_ _05870_ _05871_ _05872_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nor3_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12769_ _01802_ _01804_ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__nand2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14508_ _04727_ _04728_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__xor2_2
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15488_ _05789_ _05796_ vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__nand2_1
X_18276_ _06401_ _06546_ _08826_ _03056_ vssd1 vssd1 vccd1 vccd1 _08827_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput20 i_wb_addr[26] vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__clkbuf_1
X_17227_ _06508_ _07683_ _07684_ vssd1 vssd1 vccd1 vccd1 _07685_ sky130_fd_sc_hd__and3_1
Xinput31 i_wb_addr[7] vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_1
X_14439_ _04475_ _04477_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 i_wb_data[16] vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput53 i_wb_data[26] vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_1
Xinput64 i_wb_data[7] vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__buf_2
XFILLER_0_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17158_ _07018_ _07195_ _07608_ _06766_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16109_ _03089_ _02125_ _03179_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__or3_1
X_09980_ _07537_ _09219_ _09197_ _09205_ vssd1 vssd1 vccd1 vccd1 _09232_ sky130_fd_sc_hd__o2bb2a_1
X_17089_ _07531_ _07532_ _07507_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10120_ _00212_ vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__buf_4
X_10051_ _00126_ _00133_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__or2_1
XFILLER_0_100_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13810_ _03775_ _03780_ vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__and2_1
X_14790_ _02999_ _01112_ _04893_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__nand3_1
XFILLER_0_98_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13741_ _03718_ _03890_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__nor2_1
X_10953_ _04493_ _04416_ _00949_ _03421_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__and4_1
XFILLER_0_39_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13672_ _03625_ _03628_ _03626_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16460_ _02974_ _06847_ _06849_ _06645_ vssd1 vssd1 vccd1 vccd1 _06850_ sky130_fd_sc_hd__a211o_1
X_10884_ _00966_ _00918_ net191 vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__nor3_1
X_15411_ _05711_ _05712_ _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__o21a_1
X_12623_ _02713_ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__nand2_1
X_16391_ _06669_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15342_ _05632_ _05636_ _05637_ vssd1 vssd1 vccd1 vccd1 _05639_ sky130_fd_sc_hd__and3_1
X_18130_ _08582_ _08667_ vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__xnor2_1
X_12554_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel _00177_ _02646_
+ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__nand3_1
XFILLER_0_65_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11505_ _04045_ _01596_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15273_ _05446_ _05448_ _05561_ vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__nor3_1
X_18061_ _02175_ _08423_ _02170_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12485_ _02576_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17012_ _07345_ _07349_ _07449_ vssd1 vssd1 vccd1 vccd1 _07451_ sky130_fd_sc_hd__o21a_1
X_14224_ _03539_ _04241_ _04415_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__a31o_1
X_11436_ _04548_ _03618_ _01527_ _01528_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__nand4_2
XFILLER_0_21_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14155_ _04342_ _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__xnor2_1
X_11367_ _01455_ _01456_ _01458_ _01459_ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _02965_ _02966_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__nor2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _00403_ _00410_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__xnor2_1
X_14086_ _04100_ _04105_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__nor2_1
X_18963_ clknet_4_6_0_clk _09393_ vssd1 vssd1 vccd1 vccd1 salida\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _00794_ _01381_ _01279_ _01380_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__a211o_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _06847_ _08036_ _03197_ _05800_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__a2bb2o_1
X_13037_ _03023_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__nand2_1
X_10249_ _07363_ _09248_ vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__nand2_1
X_18894_ clknet_4_11_0_clk _00048_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17845_ _08262_ _08357_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _08281_ _08282_ vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__nand2_1
X_14988_ _05251_ _05252_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16727_ _07021_ _07045_ vssd1 vssd1 vccd1 vccd1 _07140_ sky130_fd_sc_hd__nor2_1
X_13939_ _04092_ _03945_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__o21a_2
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16658_ _06936_ _06979_ _07064_ vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15609_ _05828_ _05893_ _05927_ _05928_ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_151_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16589_ _02728_ _06988_ _06989_ vssd1 vssd1 vccd1 vccd1 _06990_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18328_ _01417_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18259_ _08804_ _08806_ vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09963_ _07232_ _07080_ _07374_ _07406_ vssd1 vssd1 vccd1 vccd1 _09101_ sky130_fd_sc_hd__and4_1
X_09894_ _03377_ _04886_ _03837_ _03356_ vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__a22o_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _02242_ _02241_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _01104_ _01116_ vssd1 vssd1 vccd1 vccd1 _01314_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11152_ cla_inst.in2\[21\] _00108_ _01241_ _01244_ vssd1 vssd1 vccd1 vccd1 _01245_
+ sky130_fd_sc_hd__o2bb2a_1
X_10103_ ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00196_ sky130_fd_sc_hd__buf_6
XFILLER_0_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11083_ _01171_ _01175_ vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__xor2_2
X_15960_ _06304_ _06305_ vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__nand2_1
X_14911_ _05167_ _05168_ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__xnor2_1
X_10034_ _09212_ vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__clkbuf_8
X_15891_ _06221_ _06222_ vssd1 vssd1 vccd1 vccd1 _06233_ sky130_fd_sc_hd__nand2_1
X_17630_ _06559_ _08123_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__or2_1
X_14842_ _03912_ _04075_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nand2_1
X_17561_ _06653_ _06756_ _08047_ vssd1 vssd1 vccd1 vccd1 _08048_ sky130_fd_sc_hd__nor3_1
X_14773_ _03014_ _05921_ _04871_ _04870_ vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__a31o_1
X_11985_ _01984_ _02054_ _02073_ _02077_ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16512_ _02828_ _02968_ _06905_ vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__or3_1
X_13724_ _03862_ _03872_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__xor2_1
X_10936_ _00936_ _00934_ _00935_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__nand3_1
X_17492_ _07971_ _07972_ vssd1 vssd1 vccd1 vccd1 _07974_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16443_ _06828_ _06831_ vssd1 vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__xor2_1
X_13655_ _08724_ _09248_ _03795_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__a22o_1
X_10867_ _03717_ _03410_ _00956_ _00959_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12606_ _02697_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__xnor2_1
X_13586_ _03674_ _03675_ _03720_ _03721_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__and4_1
X_16374_ _06563_ _06756_ vssd1 vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__nor2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _00856_ _00889_ _00890_ vssd1 vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__nor3_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _08634_ _08649_ vssd1 vssd1 vccd1 vccd1 _08650_ sky130_fd_sc_hd__xor2_1
X_15325_ _03132_ _03193_ _03536_ vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__mux2_1
X_12537_ _02616_ _02629_ vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18044_ _08573_ _08574_ vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__nand2_1
X_15256_ _05537_ _05544_ vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__or2_1
X_12468_ _02502_ _02559_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__nand2_1
X_14207_ _04399_ _04400_ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__xor2_2
X_11419_ _04984_ _00131_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__nand2_1
X_15187_ _05468_ _05469_ vssd1 vssd1 vccd1 vccd1 _05470_ sky130_fd_sc_hd__or2_1
X_12399_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _00774_ vssd1
+ vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__and2_1
X_14138_ _04319_ _04322_ _04324_ vssd1 vssd1 vccd1 vccd1 _04325_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18946_ clknet_4_2_0_clk _00100_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__dfxtp_2
X_14069_ _02975_ _03547_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18877_ clknet_4_15_0_clk net313 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__dfxtp_1
X_17828_ _06387_ _06545_ _08339_ _03041_ vssd1 vssd1 vccd1 vccd1 _08340_ sky130_fd_sc_hd__a22o_1
X_17759_ _08153_ _08154_ _08152_ vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap150 _06804_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09946_ _08822_ _08908_ vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ cla_inst.in1\[27\] vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__buf_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _00120_ _06471_ vssd1 vssd1 vccd1 vccd1 _01863_ sky130_fd_sc_hd__and2_4
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _00812_ _08071_ _06765_ _00813_ vssd1 vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ _03129_ _03168_ _03048_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__mux2_1
X_10652_ _00696_ _00697_ _00743_ _00744_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__or4_4
XFILLER_0_137_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13371_ _03485_ _03305_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10583_ _00663_ _00664_ _00675_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15110_ _05384_ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__nand2_1
X_12322_ _02346_ _02349_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__xor2_1
X_16090_ _03143_ _03056_ _06447_ vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15041_ _05285_ _05286_ vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12253_ _02344_ _02345_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or2_1
X_11204_ _01295_ _01296_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12184_ _02275_ _02224_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__and3_1
X_18800_ _02997_ net50 _09301_ vssd1 vssd1 vccd1 vccd1 _09309_ sky130_fd_sc_hd__mux2_1
X_11135_ _01217_ _01219_ _01227_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16992_ _07408_ _07323_ _07425_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__nand3_1
X_18731_ _09245_ _09254_ vssd1 vssd1 vccd1 vccd1 _09255_ sky130_fd_sc_hd__and2_1
X_11066_ _03454_ _07548_ vssd1 vssd1 vccd1 vccd1 _01159_ sky130_fd_sc_hd__and2_1
X_15943_ _06265_ _06269_ _06287_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__o21ai_1
X_10017_ _00109_ _09349_ _09188_ _07591_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__and4_1
X_18662_ _09204_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__clkbuf_1
X_15874_ _06203_ _06215_ vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17613_ _07978_ _08105_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__xnor2_1
X_14825_ _05075_ vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__inv_2
X_18593_ salida\[16\] _09141_ _09142_ salida\[48\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09153_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17544_ _06379_ _06378_ _06377_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__a21o_1
X_14756_ _04997_ _04998_ _04862_ _04969_ vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11968_ _01905_ _02058_ _02060_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13707_ _00163_ _01866_ _03853_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__and3_1
X_10919_ _01008_ _01011_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17475_ _07143_ _07721_ _07844_ _07846_ vssd1 vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__o22ai_2
X_14687_ _04922_ _04923_ _04884_ vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__a21o_1
X_11899_ _01899_ _01904_ _01991_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__or3_4
X_16426_ _06812_ net150 vssd1 vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__and2_1
X_13638_ _03776_ _03777_ _04548_ _07406_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16357_ _03089_ _02272_ _03104_ _06626_ _06737_ vssd1 vssd1 vccd1 vccd1 _06738_ sky130_fd_sc_hd__o311a_1
X_13569_ _09350_ _04154_ _00165_ _00112_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15308_ _05600_ _05601_ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16288_ _06661_ _06662_ _03324_ vssd1 vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_140_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18027_ _08455_ _08549_ _08555_ vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15239_ _05441_ _05432_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09800_ _07145_ _07178_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__nand2_1
X_09731_ _05224_ _06062_ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__nand2_1
X_18929_ clknet_4_12_0_clk _00083_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel
+ sky130_fd_sc_hd__dfxtp_1
X_09662_ _05235_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__buf_4
X_09593_ _04427_ _04569_ _04384_ _04635_ vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09929_ _08724_ _05975_ vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__nand2_1
X_12940_ _02983_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__or2_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _00908_ _02963_ _00906_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__a21o_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_101 _09395_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_112 net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _01521_ _07015_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__a22o_1
XANTENNA_123 _02783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_134 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ _04001_ _09219_ _01813_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _05855_ _05907_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__xnor2_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 _08674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ _01504_ _00461_ _04634_ _04633_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__a31o_1
X_11753_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ _01082_ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_178 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _00779_ _00794_ _00795_ _00796_ vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__a211oi_4
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _06657_ net145 _07598_ _07597_ vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__a31o_1
X_14472_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__xnor2_2
X_11684_ _01733_ _01772_ _01775_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__nor3_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ _06578_ vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__buf_2
X_10635_ _00726_ _00727_ vssd1 vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13423_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17191_ _07643_ _07644_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13354_ _03434_ _03435_ _03466_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__o21ai_2
X_16142_ _06494_ _06503_ _03080_ vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__mux2_1
X_10566_ _00634_ _00635_ _00657_ _00658_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12305_ _02397_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__inv_2
X_13285_ _03214_ _03220_ _03213_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__a21bo_1
X_16073_ _06427_ _06429_ vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__nor2_1
X_10497_ _00589_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15024_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__and2b_1
X_12236_ _02327_ _02328_ vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12167_ _01106_ _01113_ _02259_ _00398_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__or4b_4
X_11118_ _05595_ _04395_ _04886_ _05573_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__a22o_1
X_12098_ _02086_ _02084_ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__or2_1
X_16975_ _00398_ _07311_ vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__nand2_4
X_18714_ _09209_ _09241_ vssd1 vssd1 vccd1 vccd1 _09242_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11049_ _01138_ _01140_ _01141_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__and3_1
X_15926_ _06200_ _03011_ _06246_ _03154_ vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__nand4_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 i_wb_addr[14] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
X_18645_ _06427_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09192_ sky130_fd_sc_hd__a21oi_1
X_15857_ _03016_ _05652_ vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__and2_1
X_14808_ _05034_ _05035_ _05055_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__o21ai_1
X_18576_ _09097_ vssd1 vssd1 vccd1 vccd1 _09140_ sky130_fd_sc_hd__buf_2
X_15788_ _06121_ _06122_ vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17527_ _07887_ _07889_ _07885_ vssd1 vssd1 vccd1 vccd1 _08012_ sky130_fd_sc_hd__o21ba_1
X_14739_ _04979_ _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17458_ _06800_ _07934_ _07935_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__a21o_1
X_16409_ _02974_ _03119_ _03534_ _06788_ _06794_ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__o311a_1
XFILLER_0_55_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17389_ _03107_ _07592_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__nand2_4
XFILLER_0_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09714_ _04690_ _05388_ vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__nand2_1
X_09645_ _05638_ vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09576_ _04088_ _03892_ _04886_ _03903_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__and4_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10420_ _09256_ vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__buf_4
XFILLER_0_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ _03728_ _00443_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ _00517_ _03024_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__and2_1
X_10282_ _00336_ _00372_ _00373_ _00374_ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__and4b_2
X_12021_ _02112_ _02113_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03432_ vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__and4bb_1
X_16760_ _02533_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__a21o_1
X_13972_ _04123_ _04124_ _04142_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o21a_1
X_15711_ _02991_ _03071_ _06037_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__nand3_1
X_12923_ _03015_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__clkbuf_4
X_16691_ _07081_ _07082_ _07100_ vssd1 vssd1 vccd1 vccd1 _07101_ sky130_fd_sc_hd__nand3_1
X_18430_ _06409_ _07274_ _08992_ _06720_ vssd1 vssd1 vccd1 vccd1 _08993_ sky130_fd_sc_hd__o211a_1
X_15642_ _05961_ _05963_ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__or2_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _02945_ _02946_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__and2_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _01756_ _01896_ _01892_ _01895_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a211o_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _08802_ _08870_ vssd1 vssd1 vccd1 vccd1 _08918_ sky130_fd_sc_hd__nor2_1
X_15573_ _05882_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _02873_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__xnor2_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _07772_ _07774_ _07775_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__or3_1
X_14524_ _04745_ _04746_ vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__nand2_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel _00210_ vssd1
+ vssd1 vccd1 vccd1 _01829_ sky130_fd_sc_hd__and2_2
X_18292_ _00786_ _00787_ _07743_ _08774_ vssd1 vssd1 vccd1 vccd1 _08844_ sky130_fd_sc_hd__o31a_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17243_ _07666_ _07663_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ _04484_ _04670_ _04671_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__or3_2
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _01757_ _01758_ _01201_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13406_ _03367_ _03369_ _03523_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_141_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10618_ _00709_ _00710_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__xnor2_1
X_17174_ _07622_ _07625_ _07626_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__and3_1
X_14386_ _04584_ _04585_ _04595_ vssd1 vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__o21ai_2
X_11598_ _01687_ _01688_ _01689_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _03152_ _07766_ _03150_ vssd1 vssd1 vccd1 vccd1 _06486_ sky130_fd_sc_hd__nor3_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ _06711_ _07733_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__nand2_1
X_13337_ _03447_ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16056_ _03013_ _03073_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__or2_1
X_13268_ net131 _03266_ _03291_ vssd1 vssd1 vccd1 vccd1 _03373_ sky130_fd_sc_hd__nor3_2
X_15007_ _01745_ _03142_ vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ _02308_ _02311_ vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__and2b_1
X_13199_ _03298_ _03299_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16958_ _06937_ _07332_ _07390_ _06542_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_154_11 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15909_ _06251_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__nand2_1
X_16889_ _07124_ _07042_ _07313_ _06561_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__o22a_1
X_09430_ _03281_ _03206_ _03260_ _03292_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18628_ net314 _09097_ _09175_ _09176_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18559_ net301 _09098_ _09129_ _09126_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_12 _00644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_45 _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_56 _03760_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_67 _04649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 _07123_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_89 _08880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _05355_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09559_ _04690_ _04700_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ _02622_ _02659_ _02662_ vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11521_ _01174_ _01612_ _01611_ vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14240_ _04132_ _07015_ _07123_ _04099_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__a22oi_1
X_11452_ _04548_ _00211_ _01541_ _01542_ vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10403_ _00494_ _00495_ _00344_ _00343_ vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a31o_1
X_14171_ _09350_ _08409_ _00715_ _00112_ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_1_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11383_ _00877_ _00223_ _01428_ vssd1 vssd1 vccd1 vccd1 _01476_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _05845_ _03215_ _03216_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__a21bo_1
X_10334_ _09348_ _00273_ _00424_ _00426_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a211oi_4
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ _00861_ _03144_ _03023_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o21ai_1
X_17930_ _08366_ _08377_ vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__or2_1
X_10265_ cla_inst.in2\[30\] vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__buf_2
X_12004_ _02093_ _02096_ _02094_ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__o21ai_1
X_17861_ _08373_ _08374_ vssd1 vssd1 vccd1 vccd1 _08375_ sky130_fd_sc_hd__nor2_1
X_10196_ _00281_ _00287_ _00286_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__a21o_1
X_16812_ _07133_ _07136_ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__and2b_1
X_17792_ _07207_ _07780_ _07623_ _06947_ vssd1 vssd1 vccd1 vccd1 _08301_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16743_ _07154_ _07157_ vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__xnor2_2
X_13955_ _03456_ vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ _01745_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__clkbuf_4
X_16674_ _06343_ _06997_ _06342_ vssd1 vssd1 vccd1 vccd1 _07083_ sky130_fd_sc_hd__a21oi_1
X_13886_ _04004_ _04005_ _04048_ _04049_ vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__or4_4
X_18413_ _08840_ _08972_ _08974_ vssd1 vssd1 vccd1 vccd1 _08975_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ _05945_ _05946_ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__nand2_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12837_ _02928_ _02929_ vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18344_ _08848_ _08899_ vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15556_ _05781_ _05782_ _05784_ vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__o21a_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _02858_ _02859_ _01795_ _02854_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14507_ _02188_ cla_inst.in1\[31\] vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18275_ _01359_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__a21o_1
X_11719_ _01783_ _01786_ _01751_ _01785_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15487_ _05789_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ _02758_ _02791_ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17226_ _07680_ _07681_ _07682_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__nand3_1
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput10 i_wb_addr[17] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_1
X_14438_ _00115_ _05921_ _04519_ _04518_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput21 i_wb_addr[27] vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput32 i_wb_addr[8] vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput43 i_wb_data[17] vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput54 i_wb_data[27] vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__buf_1
X_17157_ _07290_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput65 i_wb_data[8] vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__buf_2
X_14369_ _04575_ _04576_ _04984_ _00498_ vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__and4bb_2
X_16108_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17088_ _07507_ _07531_ _07532_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16039_ _03000_ _03044_ vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10050_ _08202_ _08148_ _08213_ _08235_ vssd1 vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__nor4_1
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13740_ _03507_ _03510_ _03718_ _03719_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10952_ _04416_ _00949_ _03421_ _04340_ vssd1 vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__a22o_1
X_13671_ _03660_ _03665_ _03813_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__a21bo_1
X_10883_ _00974_ _00975_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15410_ _05711_ _05712_ _04238_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__a21oi_1
X_12622_ _02677_ _02714_ vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__xnor2_1
X_16390_ _06771_ _06773_ vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15341_ _01356_ _00322_ _05633_ _05634_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12553_ ApproximateM_inst.lob_16.lob2.mux.sel _00774_ vssd1 vssd1 vccd1 vccd1 _02646_
+ sky130_fd_sc_hd__and2_2
X_11504_ _05595_ _03903_ _03914_ _06019_ vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18060_ _08586_ _08589_ _08591_ vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__a21oi_2
X_15272_ _05446_ _05448_ _05561_ vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__o21a_1
X_12484_ _02568_ _02569_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17011_ _07447_ _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__and2b_1
X_14223_ _03539_ _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__nor2_1
X_11435_ _04362_ _00774_ _00909_ _04340_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ net142 _01457_ _01389_ _01387_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__o211a_1
X_14154_ _01504_ _05888_ vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__nand2_1
X_10317_ _00408_ _00409_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__xor2_1
X_13105_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__clkbuf_4
X_14085_ _04097_ _04098_ vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__and2b_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _01387_ _01388_ _01383_ _01384_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__a211o_1
X_18962_ clknet_4_6_0_clk _09392_ vssd1 vssd1 vccd1 vccd1 salida\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _08832_ _08854_ vssd1 vssd1 vccd1 vccd1 _00341_ sky130_fd_sc_hd__or2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _08427_ _08429_ _08430_ vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__nand3_1
X_13036_ _03026_ _01503_ _02805_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__a21o_1
X_18893_ clknet_4_11_0_clk _00047_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17844_ _06961_ _06957_ _07706_ _08260_ vssd1 vssd1 vccd1 vccd1 _08357_ sky130_fd_sc_hd__or4_1
X_10179_ _09344_ _09347_ _06938_ _08311_ vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__o211ai_4
X_17775_ _07194_ _07318_ _07290_ _07313_ vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__or4_2
X_14987_ _09352_ _05986_ _05249_ _05250_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__o2bb2a_1
X_16726_ _07103_ _07138_ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__xnor2_1
X_13938_ _04100_ _04105_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16657_ _06976_ _06978_ vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__and2_1
X_13869_ _09349_ _03815_ _03837_ cla_inst.in2\[27\] vssd1 vssd1 vccd1 vccd1 _04031_
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_29_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15608_ _05914_ _05926_ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16588_ _02728_ _06509_ _03169_ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18327_ _03198_ _06152_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__nand2_1
X_15539_ _05449_ _00119_ _05852_ _05849_ vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18258_ _08804_ _08806_ vssd1 vssd1 vccd1 vccd1 _08807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17209_ _07664_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18189_ _08654_ _08657_ _08652_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09962_ _07363_ _07733_ vssd1 vssd1 vccd1 vccd1 _09091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09893_ _03465_ _03815_ vssd1 vssd1 vccd1 vccd1 _08344_ sky130_fd_sc_hd__and2_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _01093_ _01103_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11151_ _01242_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10102_ _00184_ vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__clkbuf_4
X_11082_ _01172_ _01174_ vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__and2_1
X_14910_ _05038_ _05042_ _05040_ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__o21ba_1
X_10033_ _00109_ _00125_ _09212_ _09188_ vssd1 vssd1 vccd1 vccd1 _00126_ sky130_fd_sc_hd__and4_1
X_15890_ _06076_ _06079_ _06185_ _06231_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__a211o_1
X_14841_ _05080_ _05081_ _05086_ _03125_ _05092_ vssd1 vssd1 vccd1 vccd1 _09358_ sky130_fd_sc_hd__a221o_1
X_17560_ _02124_ _07825_ vssd1 vssd1 vccd1 vccd1 _08047_ sky130_fd_sc_hd__nand2_1
X_14772_ _04910_ _04911_ vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11984_ _02073_ _02075_ _02076_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nor3_1
X_16511_ _02826_ _02827_ vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__nor2_1
X_13723_ _03863_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _01026_ _01027_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__xnor2_2
X_17491_ _07866_ _07873_ vssd1 vssd1 vccd1 vccd1 _07972_ sky130_fd_sc_hd__or2b_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16442_ _06654_ _06665_ _06829_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _05508_ _05464_ _07722_ _08169_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__nand4_2
X_10866_ _00957_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12605_ _02547_ _02546_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__and2b_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _06755_ vssd1 vssd1 vccd1 vccd1 _06756_ sky130_fd_sc_hd__clkbuf_4
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _03718_ _03719_ _03507_ _03510_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__o211ai_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _08311_ _00855_ _00823_ _00854_ vssd1 vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18112_ _08646_ _08647_ vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__or2_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _05614_ _05618_ _04823_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__o21a_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12536_ _02593_ _02627_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _08565_ _08571_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__or2_1
X_15255_ _05541_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__or2_1
X_12467_ _02502_ _02559_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14206_ _04228_ _04230_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__nor2_2
XFILLER_0_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ _09188_ _01509_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__a21bo_1
X_15186_ _09352_ _00318_ _05466_ _05467_ vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12398_ _02421_ _02488_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__nor3_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14137_ _03014_ _00557_ _04321_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__a22oi_1
X_11349_ _01337_ _01377_ _01440_ _01441_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18945_ clknet_4_2_0_clk _00099_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[31\] sky130_fd_sc_hd__dfxtp_2
X_14068_ _03541_ _03545_ _03099_ vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__mux2_1
X_13019_ _03026_ _03111_ _01963_ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a21o_1
X_18876_ clknet_4_14_0_clk net315 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17827_ _02985_ _06547_ _06550_ vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17758_ _08261_ _08262_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16709_ _07028_ _07029_ vssd1 vssd1 vccd1 vccd1 _07120_ sky130_fd_sc_hd__and2b_1
X_17689_ _07038_ _07745_ vssd1 vssd1 vccd1 vccd1 _08188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap140 _01380_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_1
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09945_ _08854_ _08897_ vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _07015_ vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__clkbuf_8
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _05617_ vssd1 vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__inv_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10651_ _00741_ _00742_ _00555_ _00698_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10582_ _00666_ _00674_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__xnor2_1
X_13370_ _03302_ _03303_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12321_ _02401_ _02413_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ _05304_ _05305_ _05309_ vssd1 vssd1 vccd1 vccd1 _09360_ sky130_fd_sc_hd__o21ai_1
X_12252_ _02343_ _02336_ _02342_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ _00808_ _00807_ vssd1 vssd1 vccd1 vccd1 _01296_ sky130_fd_sc_hd__and2b_1
X_12183_ _02271_ _02273_ _02274_ _02270_ vssd1 vssd1 vccd1 vccd1 _02276_ sky130_fd_sc_hd__o31ai_1
X_11134_ _01222_ _01225_ _01226_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__or3_1
X_16991_ _07426_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11065_ _01034_ _01033_ _01032_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__a21o_1
X_18730_ _03161_ net46 _09251_ vssd1 vssd1 vccd1 vccd1 _09254_ sky130_fd_sc_hd__mux2_1
X_15942_ _06265_ _06269_ _06287_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__or3_1
X_10016_ cla_inst.in2\[27\] vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__buf_2
X_18661_ _09176_ _09203_ vssd1 vssd1 vccd1 vccd1 _09204_ sky130_fd_sc_hd__and2_1
X_15873_ _06171_ _06214_ vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__xor2_1
X_17612_ _07974_ _07992_ _07991_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__a21oi_1
X_14824_ _05071_ _05073_ _04961_ _04939_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_99_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18592_ net291 _09140_ _09151_ _09144_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__o211a_1
X_17543_ _06379_ _06377_ _06378_ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__nand3_1
X_14755_ _04862_ _04969_ _04997_ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__o211ai_1
X_11967_ _02059_ _00357_ _07613_ _04034_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _03850_ _03852_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17474_ _07950_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__xor2_1
X_10918_ _05497_ _01009_ _01010_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__a21bo_1
X_14686_ _04884_ _04922_ _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nand3_2
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ _01987_ _01990_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__and2b_1
X_16425_ sel_op\[0\] vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__inv_4
XFILLER_0_117_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13637_ _04635_ _04427_ cla_inst.in1\[25\] cla_inst.in1\[24\] vssd1 vssd1 vccd1 vccd1
+ _03777_ sky130_fd_sc_hd__and4_1
Xsplit70 _05311_ vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__clkbuf_2
X_10849_ _03990_ _00211_ _00928_ _00927_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16356_ _03027_ _00593_ _02373_ _02982_ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__a211o_1
X_13568_ _03440_ _03442_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15307_ _05459_ _05501_ _05457_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12519_ _02609_ _02610_ _02611_ vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__nand3_1
X_16287_ _00644_ net213 _06517_ vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__or3_1
X_13499_ _06029_ _05649_ cla_inst.in1\[30\] _07755_ vssd1 vssd1 vccd1 vccd1 _03626_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _08553_ _08554_ vssd1 vssd1 vccd1 vccd1 _08555_ sky130_fd_sc_hd__xor2_2
X_15238_ _05510_ _05511_ _05514_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__or3b_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15169_ _05449_ _03044_ _05447_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ _05126_ _05115_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__or2b_1
X_18928_ clknet_4_8_0_clk _00082_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_09661_ _05192_ _05203_ _05802_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__and3_1
X_18859_ clknet_4_4_0_clk net258 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__dfxtp_1
X_09592_ _04635_ _04427_ _04569_ _04449_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__and4_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09928_ _08713_ vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__clkbuf_8
X_09859_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07973_ sky130_fd_sc_hd__buf_6
X_12870_ _02959_ _02962_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__nand2_2
XFILLER_0_99_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_102 _09398_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 net49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11821_ _01814_ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 _08674_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _04762_ _04763_ vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__xnor2_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _01658_ _01666_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__xnor2_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 _05410_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 _02646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _04318_ _04755_ _04744_ vssd1 vssd1 vccd1 vccd1 _00796_ sky130_fd_sc_hd__a21oi_2
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _04544_ _04546_ vssd1 vssd1 vccd1 vccd1 _04689_ sky130_fd_sc_hd__nor2_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _01733_ _01772_ _01775_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__o21a_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _06573_ _06577_ _01106_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13422_ _03540_ _03541_ _03061_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__mux2_1
X_10634_ _00109_ _09349_ _03618_ _00171_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__and4_1
X_17190_ _07484_ _07506_ _07533_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16141_ _03099_ _06498_ _06502_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__a21oi_1
X_13353_ _03434_ _03435_ _03466_ vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__or3_4
X_10565_ _00655_ _00656_ _00636_ _00637_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12304_ _02392_ _02395_ _02311_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ _07646_ _09354_ vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _03382_ _03383_ _03389_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__a21o_1
X_10496_ _00427_ _00430_ _00587_ _00588_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15023_ _05180_ _05291_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__xnor2_2
X_12235_ _02163_ _02161_ vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12166_ _04864_ vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__clkinv_4
X_11117_ _07352_ _05322_ _01127_ _01128_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__a22o_1
X_12097_ _02189_ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__inv_2
X_16974_ _07196_ _07197_ _07294_ vssd1 vssd1 vccd1 vccd1 _07409_ sky130_fd_sc_hd__and3_1
X_18713_ net55 _06408_ _09182_ vssd1 vssd1 vccd1 vccd1 _09241_ sky130_fd_sc_hd__mux2_1
X_11048_ _01109_ _01137_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__or2_1
X_15925_ _03011_ _06246_ _03154_ _06200_ vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__a22o_1
Xinput8 i_wb_addr[15] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
X_18644_ net69 vssd1 vssd1 vccd1 vccd1 _09191_ sky130_fd_sc_hd__buf_2
X_15856_ _06194_ _06195_ vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14807_ _05034_ _05035_ _05055_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__or3_2
XFILLER_0_99_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15787_ _06053_ _06055_ _06120_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__or3_1
X_18575_ net277 _09098_ _09139_ _09126_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__o211a_1
X_12999_ _03025_ _00881_ _02646_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a21o_1
X_17526_ _08009_ _08010_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__or2_1
X_14738_ _02059_ _03455_ vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17457_ _06755_ _07621_ _07933_ net331 vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__o22a_1
X_14669_ _04780_ _04787_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16408_ _03083_ _06789_ _06793_ vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17388_ _07038_ _07649_ _07859_ _06527_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__a22o_1
X_16339_ _03539_ _06705_ _06712_ _06718_ _06484_ vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18009_ _07390_ _07650_ vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09713_ _04853_ _04875_ _04897_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__o21ba_1
X_09644_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05638_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _03739_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__clkbuf_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _05333_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _00333_ _00335_ _08681_ _09005_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ _05638_ _04220_ _00217_ _00992_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__a22oi_1
X_13971_ _04127_ _04141_ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__xnor2_2
X_15710_ _02991_ _00495_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__a21o_1
X_12922_ _03014_ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__buf_2
X_16690_ _07083_ _07085_ _07093_ _07099_ vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__o211a_1
X_15641_ _03015_ _03067_ _05962_ _05959_ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__o2bb2a_1
X_12853_ _02943_ _02944_ _02926_ _02928_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__o211ai_2
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _01892_ _01895_ _01756_ _01896_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__o211ai_2
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _08915_ _08916_ vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__and2_1
X_15572_ _05885_ _05887_ vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__or2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12784_ _02875_ _02876_ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17311_ _07772_ _07774_ _07775_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__o21a_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ _00679_ _00678_ _01575_ _00715_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__nand4_1
XFILLER_0_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _01820_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__a21o_2
XFILLER_0_127_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18291_ _08797_ _08796_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17242_ _07662_ _07661_ vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__or2b_1
X_14454_ _04667_ _04669_ _04649_ vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11666_ _01198_ _01199_ _01200_ _01181_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13405_ _03521_ _03522_ _03370_ _03347_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o211a_1
X_10617_ _00204_ _00557_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__nand2_1
X_17173_ _06581_ _07511_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__nor2_1
X_14385_ _04586_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11597_ _01687_ _01688_ _01689_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__nand3_1
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16124_ _00517_ _03156_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__nor2_1
X_13336_ _03439_ _03446_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__nand2_1
X_10548_ _00639_ _00640_ vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16055_ _06330_ _06407_ _06409_ _06024_ vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__a211oi_2
X_13267_ _03341_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__inv_2
X_10479_ _00560_ _00561_ _00571_ vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__o21ai_1
X_15006_ _05271_ _05272_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__nand2_1
X_12218_ _02309_ _02308_ _02310_ vssd1 vssd1 vccd1 vccd1 _02311_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13198_ _00189_ _00191_ _04045_ _04067_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12149_ _07036_ _07069_ _00210_ _03607_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__and4_1
XFILLER_0_138_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16957_ _07389_ vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__clkbuf_4
X_15908_ _03007_ _03072_ _06249_ _06250_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__a211o_1
XFILLER_0_154_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16888_ _06561_ _07124_ _07042_ _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__nor4_1
X_18627_ _09124_ vssd1 vssd1 vccd1 vccd1 _09176_ sky130_fd_sc_hd__buf_4
X_15839_ _06121_ _06124_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18558_ salida\[1\] _09114_ _09118_ salida\[33\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09129_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ _07975_ _07976_ _07990_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18489_ _09018_ _09021_ _09052_ _09053_ _09019_ vssd1 vssd1 vccd1 vccd1 _09056_ sky130_fd_sc_hd__o2111a_1
XANTENNA_13 _00813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_24 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_35 _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_46 _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_57 _04074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_68 _04679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _07591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09627_ _05279_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09558_ _04384_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09489_ _03760_ _03935_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ _01174_ _01611_ _01612_ vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__and3_1
XFILLER_0_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11451_ _03990_ _00146_ _01515_ _01509_ _00197_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _09311_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__buf_4
X_14170_ net219 _04155_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11382_ _01426_ _01427_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__and2b_1
XFILLER_0_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ _04121_ _05322_ _05333_ _04088_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10333_ _00421_ _00422_ _00425_ _00378_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__o2bb2a_1
X_13052_ _03025_ _03143_ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__and2_1
X_10264_ _07570_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__buf_6
X_12003_ _02094_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__nand2_1
X_10195_ _00281_ _00286_ _00287_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__nand3_1
X_17860_ _08269_ _08271_ _08372_ vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16811_ _07229_ _07230_ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17791_ _07302_ _07303_ _07511_ _07621_ vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__or4_1
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13954_ _04120_ _04122_ _03949_ _04091_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__a211oi_4
X_16742_ _06973_ net205 _07155_ vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__a21oi_2
X_12905_ _01505_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__clkbuf_4
X_16673_ _02975_ _03916_ _03120_ _04243_ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__or4_1
X_13885_ _04046_ _04047_ _04006_ _03877_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18412_ _08917_ _08918_ _08921_ _08893_ vssd1 vssd1 vccd1 vccd1 _08974_ sky130_fd_sc_hd__a22o_1
X_12836_ _02926_ _02927_ _02901_ _02922_ vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a211o_1
X_15624_ _05866_ _05870_ _05944_ vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__or3_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15555_ _05868_ _05869_ _05752_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__a21oi_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _07592_ _08896_ _08898_ vssd1 vssd1 vccd1 vccd1 _08899_ sky130_fd_sc_hd__nand3_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _01795_ _02854_ _02858_ _02859_ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _04515_ cla_inst.in1\[30\] vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__nand2_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _01751_ _01785_ _01783_ _01786_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__o211ai_2
X_18274_ _03056_ _06447_ vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15486_ _05416_ _05793_ _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _02759_ _02789_ _02790_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14437_ _04514_ _04522_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__and2_1
X_17225_ _07680_ _07681_ _07682_ vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__a21o_1
Xinput11 i_wb_addr[18] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
X_11649_ _00164_ _01357_ _01680_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__and3_1
Xinput22 i_wb_addr[28] vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput33 i_wb_addr[9] vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput44 i_wb_data[18] vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
X_17156_ _06969_ _07109_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__nand2_1
X_14368_ _03881_ _03892_ cla_inst.in1\[27\] _07004_ vssd1 vssd1 vccd1 vccd1 _04576_
+ sky130_fd_sc_hd__and4_4
Xinput55 i_wb_data[28] vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__buf_1
Xinput66 i_wb_data[9] vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__buf_2
XFILLER_0_141_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _02728_ _03022_ vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__and2b_1
X_13319_ _03428_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17087_ _07508_ _07509_ _07530_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__or3_1
XFILLER_0_150_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14299_ _04499_ _04500_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__or2b_1
X_16038_ _06389_ _06390_ _04421_ vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__a21o_1
XFILLER_0_58_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17989_ _08512_ _08513_ _08514_ vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__nand3_1
XFILLER_0_74_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10951_ _01040_ _01043_ vssd1 vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13670_ _03661_ _03664_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10882_ _08615_ _00557_ _00945_ _00944_ vssd1 vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__a31o_2
X_12621_ _07602_ _02676_ _02678_ vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__a21bo_1
X_15340_ _05635_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12552_ _02635_ _02642_ _02641_ vssd1 vssd1 vccd1 vccd1 _02645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11503_ _05573_ _05595_ _03903_ vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and3_1
X_15271_ _05557_ _05560_ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__xor2_1
X_12483_ _02574_ _02575_ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17010_ _07445_ _07446_ _07379_ _07380_ vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14222_ _03063_ _03115_ _03916_ vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11434_ _04504_ _04427_ _00217_ _00909_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__nand4_2
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14153_ _04339_ _04341_ vssd1 vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__nor2_1
X_11365_ _01387_ _01389_ _01457_ net142 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_779 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13104_ _03197_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__clkbuf_4
X_10316_ _00253_ _00213_ _00256_ _00255_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a31o_1
X_14084_ _04107_ _04108_ _04119_ vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__nor3_1
X_18961_ clknet_4_6_0_clk _09391_ vssd1 vssd1 vccd1 vccd1 salida\[14\] sky130_fd_sc_hd__dfxtp_1
X_11296_ _01383_ _01384_ _01387_ _01388_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__o211ai_4
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _08427_ _08429_ _08430_ vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__a21o_1
X_13035_ _03023_ _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__nand2_1
X_10247_ _06993_ _00339_ _09112_ _09101_ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a31o_1
X_18892_ clknet_4_11_0_clk _00046_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[10\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17843_ _08353_ _08355_ vssd1 vssd1 vccd1 vccd1 _08356_ sky130_fd_sc_hd__xor2_1
X_10178_ _00268_ _00269_ _00161_ _00231_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17774_ net146 _07604_ _07664_ _07394_ vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__a22o_1
X_14986_ _05249_ _05250_ _09352_ _05975_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__and4bb_1
X_16725_ _07111_ _07137_ vssd1 vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__xor2_1
X_13937_ _04103_ _04104_ vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__xnor2_1
X_13868_ _03818_ _03820_ vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__nor2_1
X_16656_ _06973_ _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12819_ _02909_ _02910_ _02896_ _02897_ vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__o211ai_2
X_15607_ _05914_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ _04340_ _04416_ cla_inst.in1\[26\] cla_inst.in1\[25\] vssd1 vssd1 vccd1 vccd1
+ _03954_ sky130_fd_sc_hd__and4_2
X_16587_ _03169_ _06673_ vssd1 vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18326_ _03056_ _06447_ _03143_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15538_ _05850_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__inv_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15469_ _05774_ _05775_ _05716_ _05695_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__o211a_1
X_18257_ _08655_ _08733_ _08805_ vssd1 vssd1 vccd1 vccd1 _08806_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17208_ _00247_ _07311_ _07312_ vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18188_ _08729_ _08730_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17139_ _07496_ _07505_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _06678_ _06743_ vssd1 vssd1 vccd1 vccd1 _09080_ sky130_fd_sc_hd__or2_2
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _03629_ _03596_ _04657_ _03837_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__nand4_2
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11150_ _01241_ _01242_ cla_inst.in2\[21\] _09219_ vssd1 vssd1 vccd1 vccd1 _01243_
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_101_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10101_ _00178_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__buf_6
X_11081_ _05017_ _00165_ _01172_ _01173_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__nand4_1
X_10032_ cla_inst.in2\[26\] vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__clkbuf_4
X_14840_ _05090_ _05091_ _03199_ vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__o21a_1
X_14771_ _04750_ _04915_ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__nor2_1
X_11983_ _02071_ _02072_ _02067_ _02070_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__o211a_1
X_13722_ _03864_ _03869_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16510_ _06834_ _06901_ _06903_ _06559_ vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__a211o_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _03990_ _03618_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17490_ _07872_ _07871_ vssd1 vssd1 vccd1 vccd1 _07971_ sky130_fd_sc_hd__or2b_1
X_13653_ _05366_ cla_inst.in1\[28\] _07374_ _05410_ vssd1 vssd1 vccd1 vccd1 _03795_
+ sky130_fd_sc_hd__a22o_1
X_16441_ _06771_ _06773_ vssd1 vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__or2b_1
X_10865_ _00956_ _00957_ _03717_ _03410_ vssd1 vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__and4b_1
XFILLER_0_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12604_ _08865_ _01503_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__nand2_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16372_ _02977_ _06753_ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13584_ _03507_ _03510_ _03718_ _03719_ vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__a211o_1
X_10796_ _00859_ _00888_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__xnor2_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _05614_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18111_ _08635_ _08645_ vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__nor2_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ _02593_ _02627_ vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__or2b_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ _05449_ _01139_ _05542_ _05538_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__o2bb2a_1
X_18042_ _08565_ _08571_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__nand2_1
X_12466_ _07700_ _07799_ _00212_ _00206_ vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__and4_2
XFILLER_0_81_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14205_ _04397_ _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__nand2_2
XFILLER_0_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ _01151_ _01031_ _09179_ _04078_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a22o_1
X_15185_ _05466_ _05467_ _09352_ _07134_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__and4bb_1
X_12397_ _02489_ _02214_ _02419_ _02420_ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__o22a_1
X_14136_ _04320_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11348_ _01415_ _01439_ _01438_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__o21ai_2
X_18944_ clknet_4_2_0_clk _00098_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[30\] sky130_fd_sc_hd__dfxtp_1
X_14067_ _04245_ _04246_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__mux2_1
X_11279_ _01251_ _01270_ vssd1 vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__nand2_1
X_13018_ _01866_ vssd1 vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__clkbuf_4
X_18875_ clknet_4_14_0_clk net316 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__dfxtp_1
X_17826_ _03041_ _06443_ _08337_ vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _02200_ _06891_ _06969_ _08150_ vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__and4_1
X_14969_ _03008_ _00678_ _05878_ _06471_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__and4_1
X_16708_ _07117_ _07118_ vssd1 vssd1 vccd1 vccd1 _07119_ sky130_fd_sc_hd__nor2_1
X_17688_ _07038_ _07623_ _08095_ _08186_ vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__a31o_1
XFILLER_0_147_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16639_ _07041_ _07043_ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18309_ _08785_ _08791_ _08861_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap130 _02071_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_1
XFILLER_0_130_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap141 net325 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_1
XFILLER_0_111_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09944_ _08865_ _08876_ _08887_ _08843_ vssd1 vssd1 vccd1 vccd1 _08897_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _07635_ _07657_ vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__nand2_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10650_ _00555_ _00698_ _00741_ _00742_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10581_ _00672_ _00673_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12320_ _02411_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12251_ _02336_ _02342_ _02343_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__a21oi_1
X_11202_ _05224_ _05050_ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__nand2_1
X_12182_ _02270_ _02271_ _02273_ _02274_ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__or4_4
X_11133_ _01137_ _01221_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__and2_1
X_16990_ _07408_ _07323_ _07425_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__a21oi_2
X_11064_ _01034_ _01032_ _01033_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__nand3_1
X_15941_ _06284_ _06286_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__xnor2_2
X_10015_ _09219_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__clkbuf_4
X_18660_ net64 _00881_ _09193_ vssd1 vssd1 vccd1 vccd1 _09203_ sky130_fd_sc_hd__mux2_1
X_15872_ _06211_ _06212_ vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__nor2_1
X_17611_ _08101_ _08102_ vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__nand2_1
X_14823_ _04961_ _04939_ _05071_ _05073_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__o211ai_2
X_18591_ salida\[15\] _09141_ _09142_ salida\[47\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09151_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17542_ _08025_ _08026_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__or2_1
X_14754_ _04992_ _04993_ _04996_ vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__nand3_2
X_11966_ _03728_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__buf_8
XFILLER_0_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10917_ _05638_ _05377_ _05028_ _00992_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__a22o_1
X_13705_ _03851_ _03687_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__nand2_1
X_14685_ _04920_ _04921_ _04902_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__a21o_1
X_17473_ _07833_ _07838_ _07952_ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__o21ai_2
X_11897_ _01988_ _01987_ _01989_ vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__or3_4
X_13636_ _00294_ _07102_ cla_inst.in1\[24\] _04351_ vssd1 vssd1 vccd1 vccd1 _03776_
+ sky130_fd_sc_hd__a22oi_1
X_16424_ _00210_ _06528_ _06530_ _06810_ sel_op\[0\] vssd1 vssd1 vccd1 vccd1 _06811_
+ sky130_fd_sc_hd__o32a_1
X_10848_ _00925_ _00926_ _00940_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13567_ _00115_ _00247_ _03500_ _03499_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__a31o_1
XFILLER_0_109_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16355_ _03049_ _06622_ _06735_ _06626_ vssd1 vssd1 vccd1 vccd1 _06736_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10779_ cla_inst.in2\[24\] _00174_ _00196_ _00871_ vssd1 vssd1 vccd1 vccd1 _00872_
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_125_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15306_ _05598_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__nand2_1
X_12518_ _02559_ _02608_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16286_ _03281_ _03003_ _06520_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13498_ _05649_ _09256_ _09303_ _06029_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18025_ _07108_ _07745_ vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__nand2_1
X_15237_ _05428_ _05396_ _05509_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__a21o_1
X_12449_ _02540_ _02541_ vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15168_ _07635_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14119_ _00644_ _02476_ _03455_ _00513_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__and4_1
X_15099_ _05265_ _05269_ _05266_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18927_ clknet_4_13_0_clk _00081_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ _05192_ _05203_ _05802_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__a21oi_4
X_18858_ clknet_4_7_0_clk net280 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__dfxtp_1
X_17809_ _08208_ _08210_ _08206_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__a21o_1
X_09591_ _05017_ _05050_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__nand2_1
X_18789_ _09300_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09927_ _05213_ vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__buf_4
X_09858_ cla_inst.in1\[24\] vssd1 vssd1 vccd1 vccd1 _07962_ sky130_fd_sc_hd__clkbuf_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _07178_ _07189_ _07199_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__nand3_4
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _01908_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__xor2_1
XANTENNA_103 _09399_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_114 net69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 _02987_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ _01828_ _01841_ _01842_ net138 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a211oi_2
XANTENNA_169 _06555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _04318_ _04744_ _04755_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__and3_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _04686_ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__or2b_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11682_ _01729_ _01774_ vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__xnor2_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13421_ _03058_ _03070_ _03049_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__mux2_1
X_10633_ _00149_ _00206_ _00172_ _00151_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _00494_ _06470_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__and3_1
X_13352_ _03437_ _03464_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _00636_ _00637_ _00655_ _00656_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_107_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _02308_ _02310_ _02309_ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16071_ _00127_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__clkinv_4
X_13283_ _03382_ _03383_ _03389_ vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__nand3_1
X_10495_ _00585_ _00586_ _00418_ _00421_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_106_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ _05288_ _05289_ vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ _02324_ _02323_ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12165_ _07853_ _00557_ _02257_ vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__and3_2
X_11116_ _01206_ _01208_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__nand2_1
X_12096_ _02188_ _05017_ _07559_ _07602_ vssd1 vssd1 vccd1 vccd1 _02189_ sky130_fd_sc_hd__and4_1
X_16973_ _07307_ _07309_ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__nand2_1
X_18712_ _09239_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__clkbuf_1
X_11047_ _00845_ _01139_ _01108_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__a21o_2
X_15924_ _06260_ _06261_ vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__nor2_1
Xinput9 i_wb_addr[16] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_1
X_18643_ _09183_ vssd1 vssd1 vccd1 vccd1 _09190_ sky130_fd_sc_hd__buf_2
X_15855_ _03010_ _03013_ _03154_ _03072_ vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14806_ _05053_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__xnor2_2
X_18574_ salida\[9\] _09114_ _09118_ salida\[41\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09139_ sky130_fd_sc_hd__a221o_1
X_15786_ _06053_ _06055_ _06120_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12998_ _03085_ _03088_ _03090_ vssd1 vssd1 vccd1 vccd1 _03091_ sky130_fd_sc_hd__mux2_1
X_17525_ _07881_ _07891_ _08008_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14737_ _04977_ _04978_ vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__nor2_1
X_11949_ _02028_ _02041_ vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17456_ _02127_ _07933_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14668_ _04781_ _04786_ vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16407_ _06336_ _06790_ _06792_ _06543_ _06461_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__a221o_1
X_13619_ _03454_ _05311_ vssd1 vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__and2_1
XFILLER_0_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17387_ _02044_ _07743_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__nor2_4
X_14599_ _04827_ _04828_ _03538_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16338_ _03547_ _06717_ _03117_ vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a21o_1
X_16269_ _03547_ _06642_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _08533_ _08534_ vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09712_ _06340_ _06351_ _06362_ vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__nand3_4
X_09643_ _05573_ _05595_ _05606_ _05617_ vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _04121_ _04657_ _04864_ _04088_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10280_ _09152_ _09338_ _00370_ _00371_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_131_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13970_ _04139_ _04140_ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__nor2_1
X_12921_ _00362_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15640_ _05960_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__inv_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _02926_ _02928_ _02943_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a211o_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _01741_ _01755_ _01754_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a21o_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15571_ _03015_ _03142_ _05886_ _05883_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _02858_ _02860_ vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__nor2_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _07625_ _07626_ _07622_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__a21bo_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14522_ _00678_ _08409_ _00715_ _00679_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__a22o_1
X_11734_ _01594_ _01599_ vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__xnor2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _08736_ _08809_ _08749_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_139_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17241_ _02127_ _06723_ _07675_ _07699_ vssd1 vssd1 vccd1 vccd1 _09390_ sky130_fd_sc_hd__o22a_1
X_14453_ _04649_ _04667_ _04669_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor3_1
X_11665_ _01710_ _01716_ _01717_ _01718_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__and4_1
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13404_ _03370_ _03347_ _03521_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__a211oi_4
X_10616_ _00707_ _00708_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__xor2_2
X_14384_ _04587_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17172_ _07038_ net146 _07623_ _06527_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__a22o_1
X_11596_ _01646_ _01653_ _01652_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13335_ _03439_ _03446_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16123_ _06483_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__clkbuf_4
X_10547_ _06029_ _06051_ _07384_ _07015_ vssd1 vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__and4_1
XFILLER_0_134_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ _00661_ net327 _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__o211a_1
X_16054_ _03016_ _06408_ vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__nor2_1
X_10478_ _00562_ _00570_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__xnor2_1
X_15005_ _05270_ _05264_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or2b_1
X_12217_ _02306_ _02307_ _02295_ _02299_ vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__a211oi_1
X_13197_ _00191_ _00398_ _00247_ _00189_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a22oi_1
X_12148_ _07069_ _00210_ _03607_ _07036_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12079_ _01810_ _01903_ _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__a21o_1
X_16956_ _04034_ _03324_ _06814_ _07386_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__a211oi_2
X_15907_ _06249_ _06250_ _06200_ _03072_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__o211ai_1
X_16887_ _07313_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ salida\[30\] _09113_ _09117_ salida\[62\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09175_ sky130_fd_sc_hd__a221o_2
XFILLER_0_154_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15838_ _06175_ _06176_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18557_ _09127_ vssd1 vssd1 vccd1 vccd1 _09128_ sky130_fd_sc_hd__buf_2
X_15769_ _01417_ _04125_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17508_ _07975_ _07976_ _07990_ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18488_ _09052_ _09053_ _09054_ vssd1 vssd1 vccd1 vccd1 _09055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_14 _01108_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _03108_ _06440_ vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__nor2_1
XANTENNA_25 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_36 _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_47 _02969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_58 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_69 _05625_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput110 net110 vssd1 vssd1 vccd1 vccd1 o_wb_data[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ _05268_ _05431_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__xnor2_2
X_09557_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04690_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09488_ _03870_ _03925_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11450_ _04690_ _00211_ _01541_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__nand4_2
XFILLER_0_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _06993_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11381_ _00163_ _00881_ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _04088_ _04121_ _05333_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__and3_1
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ net338 _00377_ _09346_ _00274_ vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13051_ _03142_ vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__clkbuf_4
X_10263_ _00353_ _00354_ _09271_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__o21ai_1
X_12002_ _05301_ _00180_ _00130_ _05279_ vssd1 vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__a22o_1
X_10194_ _00278_ _00279_ _00280_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16810_ _07193_ _07228_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__nand2_1
X_17790_ _08173_ _08178_ _08297_ vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__a21oi_1
X_16741_ _07059_ _07061_ vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__and2b_1
X_13953_ _03949_ _04091_ _04120_ _04122_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__o211a_4
X_12904_ _02996_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__buf_2
X_16672_ _06426_ _06435_ _07076_ _07079_ vssd1 vssd1 vccd1 vccd1 _07081_ sky130_fd_sc_hd__o31a_1
X_13884_ _04006_ _03877_ _04046_ _04047_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__a211oi_2
X_18411_ _08872_ _08921_ vssd1 vssd1 vccd1 vccd1 _08972_ sky130_fd_sc_hd__or2b_1
X_15623_ _05866_ _05870_ _05944_ vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _02901_ _02922_ _02926_ _02927_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__o211ai_4
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _06374_ _00558_ _04995_ vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__a21o_1
X_15554_ _05752_ _05868_ _05869_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__and3_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _02856_ _02857_ _01790_ _02855_ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__a211oi_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14505_ _08615_ _03456_ _04589_ _04588_ _04725_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__a32o_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _07084_ _08821_ _08823_ vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11717_ _01808_ _01809_ vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__nor2_4
X_15485_ _05612_ _05708_ _05709_ _05794_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__o211a_1
X_12697_ _02756_ _02757_ _02758_ _02754_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ _07566_ _07567_ _07565_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_582 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14436_ _04516_ _04521_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__and2b_1
X_11648_ _01642_ net125 _01739_ _01740_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__o211ai_4
Xinput12 i_wb_addr[19] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput23 i_wb_addr[29] vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 i_wb_cyc vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_2
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput45 i_wb_data[19] vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_2
X_17155_ _06891_ _07109_ _07499_ _07605_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__a31o_1
XFILLER_0_142_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14367_ _03793_ _07374_ _07406_ _03859_ vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__a22oi_1
X_11579_ _07799_ _05845_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__and2_2
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput56 i_wb_data[29] vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_1
Xinput67 i_wb_stb vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_4
X_16106_ _03121_ _06454_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__nor2_1
X_13318_ _03254_ _03256_ _03426_ _03427_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__a211oi_4
X_14298_ _04339_ _04343_ _04341_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__o21ba_1
X_17086_ _07508_ _07509_ _07530_ vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_110_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16037_ _00592_ _04336_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__or2_2
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ _03351_ _03352_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17988_ _08429_ _08430_ _08427_ vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__a21bo_1
X_16939_ _03079_ _06698_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18609_ net257 _09157_ _09164_ _09162_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _01041_ _01042_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__xnor2_2
X_09609_ _05246_ vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__buf_4
X_10881_ _00968_ _00973_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12620_ _07091_ _07363_ _07570_ _07602_ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__and4_1
X_12551_ _02635_ _02641_ _02642_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__nand3_1
XFILLER_0_108_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11502_ _06711_ _00715_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15270_ _01317_ _05558_ _05559_ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_108_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12482_ _02504_ _02571_ _02573_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__nand3_1
XFILLER_0_62_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11433_ _01514_ _01524_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__xor2_1
X_14221_ _03078_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14152_ _00190_ _00192_ _06482_ _04591_ vssd1 vssd1 vccd1 vccd1 _04341_ sky130_fd_sc_hd__and4_1
X_11364_ _00123_ _00848_ _00849_ vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ _00404_ _00407_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__xnor2_1
X_13103_ _03036_ _03123_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__nor2_2
XFILLER_0_132_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14083_ _04261_ _04264_ _03539_ vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__mux2_1
X_18960_ clknet_4_6_0_clk _09390_ vssd1 vssd1 vccd1 vccd1 salida\[13\] sky130_fd_sc_hd__dfxtp_1
X_11295_ _01385_ _01284_ _01386_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__nand3_2
XFILLER_0_131_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _08330_ _08331_ _08329_ vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__o21bai_2
X_13034_ _03028_ _02779_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__nor2_1
X_10246_ _07744_ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__buf_4
XFILLER_0_28_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18891_ clknet_4_11_0_clk _00045_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_17842_ net146 net145 vssd1 vssd1 vccd1 vccd1 _08355_ sky130_fd_sc_hd__nand2_1
X_10177_ _00161_ _00231_ _00268_ _00269_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__a211o_2
X_17773_ _08162_ _08163_ _08161_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__o21ai_2
X_14985_ _00148_ _00149_ _06062_ _05257_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__and4_1
X_16724_ _07133_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__xor2_1
X_13936_ _04001_ _07123_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16655_ _07059_ _07061_ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__xnor2_1
X_13867_ _00107_ _04012_ _03867_ _03866_ vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__a31o_1
X_15606_ _05924_ _05925_ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12818_ _02896_ _02897_ _02909_ _02910_ vssd1 vssd1 vccd1 vccd1 _02911_ sky130_fd_sc_hd__a211o_1
X_16586_ _03206_ _06986_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__nor2_1
X_13798_ _00294_ _07004_ _07102_ _04504_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__a22oi_1
X_18325_ _03201_ _08878_ _08879_ vssd1 vssd1 vccd1 vccd1 _08880_ sky130_fd_sc_hd__and3_2
X_15537_ _05849_ _00119_ _05449_ _05850_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__and4b_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _02751_ _02836_ _02839_ _02841_ vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__o31a_1
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18256_ _08732_ _08731_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__or2b_1
X_15468_ _05716_ _05695_ _05774_ _05775_ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17207_ _07661_ _07662_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__xnor2_1
X_14419_ _00702_ _05486_ _05878_ _00195_ vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_53_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18187_ _08636_ _08644_ _08646_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__a21oi_1
X_15399_ _05499_ _05602_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17138_ _07552_ _07553_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09960_ _06993_ _09059_ _07428_ _07417_ vssd1 vssd1 vccd1 vccd1 _09070_ sky130_fd_sc_hd__a31o_1
X_17069_ _07124_ _07126_ _07511_ _06561_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _06373_ _06504_ _06515_ vssd1 vssd1 vccd1 vccd1 _08322_ sky130_fd_sc_hd__nand3_2
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ _00147_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__buf_4
X_11080_ _00294_ _00210_ _00205_ _04504_ vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__a22o_1
X_10031_ _00110_ _00114_ vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _05012_ _05013_ _04867_ _04968_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__o211ai_2
X_11982_ _02053_ _02074_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__nand2_1
X_13721_ _03867_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__xnor2_1
X_10933_ _01024_ _01025_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16440_ _06824_ _06827_ vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__xnor2_1
X_13652_ _03791_ _03792_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__nor2_1
X_10864_ ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel cla_inst.in2\[16\] vssd1
+ vssd1 vccd1 vccd1 _00957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ _02672_ _02673_ _02692_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a21oi_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _03324_ _06752_ net343 vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o21ai_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _03715_ _03716_ _03676_ _03677_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__a211oi_2
X_10795_ _00860_ _00865_ _00867_ _00887_ vssd1 vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ _08635_ _08645_ vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__and2_1
X_15322_ _05416_ _05615_ _05616_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__a21oi_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _02618_ _02625_ _02626_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__o21ai_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18041_ _08490_ _08570_ vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__xnor2_1
X_15253_ _05539_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__inv_2
X_12465_ _02544_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__xnor2_1
X_14204_ _04393_ _04394_ _04396_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11416_ _04078_ _01151_ _00871_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__and3_1
X_15184_ _00148_ _00149_ _00308_ _05964_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__and4_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12396_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _02489_ sky130_fd_sc_hd__inv_4
XFILLER_0_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14135_ _04320_ _04012_ _00362_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__and4b_1
XFILLER_0_10_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11347_ _01415_ _01438_ _01439_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__or3_4
XFILLER_0_39_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18943_ clknet_4_2_0_clk _00097_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[29\] sky130_fd_sc_hd__dfxtp_2
X_11278_ _01252_ _01269_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__or2b_1
X_14066_ _03079_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__clkbuf_4
X_10229_ _07025_ vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__buf_4
X_13017_ _03040_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__nand2_1
X_18874_ clknet_4_15_0_clk net249 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__dfxtp_1
X_17825_ _03041_ _06443_ _06424_ vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__a21oi_1
X_17756_ _06961_ _07706_ _08260_ _07018_ vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__o22a_1
X_14968_ _05230_ vssd1 vssd1 vccd1 vccd1 _05231_ sky130_fd_sc_hd__inv_2
X_16707_ _06766_ _06875_ _07114_ _07116_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__o22a_1
X_13919_ _03538_ _03124_ _04076_ _04085_ _03199_ vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__a32o_1
X_17687_ _08094_ _08092_ vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__and2b_1
X_14899_ _05018_ _05027_ _05025_ vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16638_ _06579_ _07042_ vssd1 vssd1 vccd1 vccd1 _07043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16569_ _06878_ _06879_ _00194_ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18308_ _08859_ _08860_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18239_ _08784_ _08785_ vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap120 net319 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_1
XFILLER_0_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09943_ _08832_ vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _07319_ _07940_ _08115_ vssd1 vssd1 vccd1 vccd1 _08137_ sky130_fd_sc_hd__a21o_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10580_ _00670_ _00671_ _00667_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _02218_ _02220_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ _00974_ _00975_ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12181_ _02128_ _02258_ vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__and2_1
X_11132_ _07853_ _01223_ _01224_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__a21oi_4
X_11063_ _01154_ _01155_ vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__xnor2_1
X_15940_ _06258_ _06285_ vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__nand2_1
X_10014_ _00106_ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__clkbuf_4
X_15871_ _06209_ _06210_ vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__and2_1
X_17610_ _08099_ _08100_ vssd1 vssd1 vccd1 vccd1 _08102_ sky130_fd_sc_hd__nand2_1
X_14822_ _05069_ _05070_ _04896_ _04963_ vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__a211o_1
X_18590_ net285 _09140_ _09150_ _09144_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17541_ _08025_ _08026_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__nand2_1
X_14753_ _04992_ _04993_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11965_ _02007_ _02057_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13704_ _03682_ _03683_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__or2b_1
X_10916_ _00992_ _05638_ net235 vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__and3_1
X_17472_ _07707_ _07832_ vssd1 vssd1 vccd1 vccd1 _07952_ sky130_fd_sc_hd__or2_1
X_14684_ _04902_ _04920_ _04921_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__nand3_1
X_11896_ _01986_ _01980_ _01984_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__and3_1
X_16423_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ _03184_ vssd1 vssd1 vccd1 vccd1 _06810_ sky130_fd_sc_hd__o41a_1
X_13635_ _03600_ _03601_ _03599_ vssd1 vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ _00931_ _00938_ _00939_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16354_ _01677_ _06637_ vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__or2_1
X_13566_ _03495_ _03503_ _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10778_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00871_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15305_ _05596_ _05597_ _05552_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12517_ _00120_ _00213_ _00207_ _07711_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16285_ _02728_ net344 vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__nor2_1
X_13497_ _03395_ _03403_ _03402_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18024_ _08551_ _08552_ vssd1 vssd1 vccd1 vccd1 _08553_ sky130_fd_sc_hd__nand2_2
X_15236_ _03082_ _05307_ _05425_ _03039_ _05523_ vssd1 vssd1 vccd1 vccd1 _09362_ sky130_fd_sc_hd__o221ai_2
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _02501_ _02507_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15167_ _03014_ _01223_ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _02458_ _02459_ _02452_ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14118_ _02476_ _03456_ _00665_ _00644_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15098_ _05371_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14049_ _04225_ _04226_ _04227_ vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__and3_2
X_18926_ clknet_4_13_0_clk _00080_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_18857_ clknet_4_4_0_clk net266 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__dfxtp_1
X_17808_ _08316_ _08317_ vssd1 vssd1 vccd1 vccd1 _08318_ sky130_fd_sc_hd__xor2_1
X_09590_ _05039_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__clkbuf_8
X_18788_ _09298_ _09299_ vssd1 vssd1 vccd1 vccd1 _09300_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17739_ _02973_ _06645_ vssd1 vssd1 vccd1 vccd1 _08243_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09926_ _06493_ _06450_ vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__or2b_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _07036_ _07069_ _05693_ cla_inst.in1\[22\] vssd1 vssd1 vccd1 vccd1 _07951_
+ sky130_fd_sc_hd__nand4_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _06993_ _07025_ _07145_ _07167_ vssd1 vssd1 vccd1 vccd1 _07199_ sky130_fd_sc_hd__a22o_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 _09402_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_115 net82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _03201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_137 _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _01670_ _01676_ _01679_ _01680_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nor4_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10701_ _00779_ _00792_ _00793_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__nand3_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _01507_ _01773_ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__or2b_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13420_ _03046_ _03054_ _03049_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__mux2_1
X_10632_ _07537_ _00147_ _00520_ _00359_ _00132_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__a32o_1
XFILLER_0_64_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10563_ _00653_ _00654_ _00638_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__a21bo_1
X_13351_ _03438_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12302_ _02393_ _02392_ _02394_ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__nor3_1
X_16070_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _03386_ _03387_ vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__xor2_2
X_10494_ _00418_ _00421_ _00585_ _00586_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _05139_ _05183_ _05136_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__a21oi_2
X_12233_ _02321_ _02325_ vssd1 vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12164_ _00515_ _02127_ vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11115_ _06982_ _00443_ _01206_ _01207_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__nand4_2
X_12095_ _04373_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__clkbuf_8
X_16972_ _07385_ _07405_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__xnor2_1
X_11046_ _05986_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__clkbuf_4
X_18711_ _09209_ _09238_ vssd1 vssd1 vccd1 vccd1 _09239_ sky130_fd_sc_hd__and2_1
X_15923_ _02969_ _06264_ _06265_ _06268_ vssd1 vssd1 vccd1 vccd1 _09374_ sky130_fd_sc_hd__o31ai_4
X_18642_ _09183_ vssd1 vssd1 vccd1 vccd1 _09189_ sky130_fd_sc_hd__buf_2
X_15854_ _03012_ _03154_ _03072_ _03010_ vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__a22o_1
X_14805_ _01873_ _03055_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18573_ net271 _09098_ _09138_ _09126_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__o211a_1
X_15785_ _06118_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__and2_1
X_12997_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__clkbuf_4
X_17524_ _07881_ _07891_ _08008_ vssd1 vssd1 vccd1 vccd1 _08009_ sky130_fd_sc_hd__a21oi_2
X_14736_ _04099_ _04034_ _00502_ _09248_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11948_ _02031_ _02039_ _02040_ vssd1 vssd1 vccd1 vccd1 _02041_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17455_ _04034_ _06889_ vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__nand2_1
X_14667_ _04619_ _04789_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11879_ _01869_ _01970_ _01938_ _01969_ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16406_ _06431_ _06791_ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__nor2_1
X_13618_ _03531_ _03509_ _06613_ net223 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17386_ _07856_ _07857_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _03916_ _03546_ vssd1 vssd1 vccd1 vccd1 _04828_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16337_ _03164_ _06470_ _06713_ _06716_ vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__a31o_1
X_13549_ _00169_ _08409_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16268_ _06639_ _06641_ _03061_ vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18007_ _07665_ _07596_ _08453_ vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__and3_1
X_15219_ _05503_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16199_ _03410_ _03673_ _06529_ _06565_ vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__or4_4
XFILLER_0_77_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09711_ _04919_ _04930_ _04842_ vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__a21bo_1
X_18909_ clknet_4_10_0_clk _00063_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[27\] sky130_fd_sc_hd__dfxtp_4
X_09642_ cla_inst.in1\[21\] vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09573_ _03804_ vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__buf_6
XFILLER_0_96_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _06319_ _06329_ _06267_ vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__a21bo_1
X_12920_ _03012_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__clkbuf_4
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _00893_ _00897_ _00895_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a21oi_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _01892_ _01893_ _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__nor3_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _05884_ vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__inv_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _01374_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer90 _00925_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14521_ _03005_ _00557_ vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__nand2_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _01824_ _01825_ vssd1 vssd1 vccd1 vccd1 _01826_ sky130_fd_sc_hd__or2b_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _07678_ _07685_ _07696_ _07698_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__or4b_1
X_14452_ _04650_ _04525_ _04666_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__and3_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _01610_ _01619_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13403_ _03518_ _03519_ _03337_ _03339_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10615_ _00564_ _00567_ _00565_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_107_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17171_ _02127_ _06814_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__nor2_4
XFILLER_0_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14383_ _04590_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__xor2_1
X_11595_ _01684_ _01686_ _01685_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16122_ _08865_ _02965_ _06422_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nor3_1
X_13334_ _03442_ _03445_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__or2_1
X_10546_ _06084_ _07384_ _08158_ _06040_ vssd1 vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16053_ _03149_ vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13265_ _00696_ net320 _03341_ _03342_ vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10477_ _00568_ _00569_ vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15004_ _05264_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12216_ _02277_ _02279_ _02274_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ _00737_ _00739_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12147_ _02234_ _02239_ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__xnor2_1
X_12078_ _01995_ _01996_ _01999_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__o22ai_1
X_16955_ _06563_ _06756_ _07332_ _07387_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__or4_1
X_11029_ _08039_ _04449_ _04471_ _00992_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__a22o_1
X_15906_ _03013_ _06246_ _06248_ vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16886_ _00247_ _07311_ _07312_ vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__nand3_4
X_15837_ _06161_ _06174_ vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__nor2_1
X_18625_ net303 _09157_ _09174_ _09162_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__o211a_1
X_15768_ _02991_ _03153_ vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__nand2_1
X_18556_ net68 _09096_ vssd1 vssd1 vccd1 vccd1 _09127_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14719_ _03121_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__nor2_1
X_17507_ _07979_ _07989_ vssd1 vssd1 vccd1 vccd1 _07990_ sky130_fd_sc_hd__xnor2_1
X_18487_ _09018_ _09021_ _09019_ vssd1 vssd1 vccd1 vccd1 _09054_ sky130_fd_sc_hd__o21a_1
X_15699_ _03009_ _03012_ _09059_ _00322_ vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__and4_1
X_17438_ _07910_ _07914_ _07912_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 _02989_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17369_ _07833_ _07838_ vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__xnor2_2
XANTENNA_59 _04406_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput100 net100 vssd1 vssd1 vccd1 vccd1 o_wb_data[25] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput111 net111 vssd1 vssd1 vccd1 vccd1 o_wb_data[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09625_ _05344_ _05421_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__and2b_1
X_09556_ _04438_ _04482_ _04657_ _04646_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09487_ _03881_ _03892_ _03903_ _03914_ vssd1 vssd1 vccd1 vccd1 _03925_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10400_ _00340_ _00347_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ _01470_ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__xor2_1
XFILLER_0_150_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10331_ _00378_ _00421_ _00422_ _00423_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__and4b_2
XFILLER_0_103_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10262_ _00353_ _09271_ _00354_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__or3_1
X_13050_ _00322_ vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__buf_2
X_12001_ _05410_ _05301_ _00146_ _00197_ vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__nand4_1
X_10193_ _00284_ _00285_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16740_ _07152_ _07153_ vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__xnor2_2
X_13952_ _04107_ _04108_ _04119_ vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__or3_4
X_12903_ _00191_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__clkbuf_4
X_16671_ _06462_ _07078_ vssd1 vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__nor2_1
X_13883_ _04043_ _04044_ _03828_ _04007_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__o211a_1
X_15622_ _05941_ _05942_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and2_1
X_18410_ _08969_ _08970_ vssd1 vssd1 vccd1 vccd1 _08971_ sky130_fd_sc_hd__or2_1
X_12834_ _02924_ _02925_ _02923_ _02907_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__a211o_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _08895_ _04023_ _07743_ vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__or3_1
X_15553_ _05864_ _05865_ _05776_ _05778_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__a211o_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _01790_ _02855_ _02856_ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__o211a_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14504_ _04515_ vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__buf_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _05557_ _06401_ _06400_ vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__a21oi_1
X_11716_ _01806_ _01807_ _01507_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a21oi_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _05616_ _05790_ vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__nand2_1
X_12696_ _02782_ _02786_ _02787_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__and4_1
XFILLER_0_126_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17223_ _06368_ _07355_ _04725_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__or3b_1
X_14435_ _04325_ _04523_ vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11647_ _01721_ _01738_ _01737_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__a21o_1
Xinput13 i_wb_addr[1] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput24 i_wb_addr[2] vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_2
XFILLER_0_25_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17154_ _06657_ _07604_ _07498_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__and3_1
Xinput35 i_wb_data[0] vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14366_ _04571_ _04572_ _04567_ net333 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__a211o_1
Xinput46 i_wb_data[1] vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
X_11578_ _05878_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput57 i_wb_data[2] vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_4
Xinput68 i_wb_we vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_4
XFILLER_0_40_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__clkbuf_4
X_13317_ _03424_ _03425_ _03411_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a21oi_2
X_10529_ _00451_ _00453_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__nand2_1
X_17085_ _07510_ _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__xor2_1
X_14297_ _04497_ _04498_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__xnor2_1
X_16036_ _06386_ _06387_ _06388_ vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__a21bo_1
X_13248_ _00713_ _00717_ _00712_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _03276_ _03277_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__and2_1
X_17987_ _03044_ _08428_ _03000_ vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__or3b_2
X_16938_ _06704_ _06710_ _03079_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16869_ _07292_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__xnor2_2
X_18608_ salida\[21\] _09159_ _09160_ salida\[53\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18539_ net148 vssd1 vssd1 vccd1 vccd1 _09109_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09608_ cla_inst.in1\[20\] vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__clkbuf_8
X_10880_ _00969_ _00972_ vssd1 vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ ApproximateM_inst.lob_16.lob2.genblk1\[13\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04493_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _02635_ _02641_ _02642_ vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11501_ _01589_ _01592_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12481_ _02571_ _02573_ _02504_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14220_ _02975_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__nor2_2
X_11432_ _01514_ _01524_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14151_ _00192_ _06482_ _05921_ _00190_ vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a22oi_1
X_11363_ _01396_ _01404_ _01397_ _01398_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__or4_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _03194_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__inv_2
X_10314_ _00405_ _00406_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__and2b_1
X_14082_ _03547_ _04262_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nor2_1
X_11294_ _01385_ _01284_ _01386_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__a21o_2
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17910_ _04336_ _08428_ _03368_ vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__or3b_1
X_13033_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__clkbuf_4
X_10245_ _09070_ _09137_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18890_ clknet_4_13_0_clk _00044_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10176_ _00267_ _00266_ _08289_ _07919_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__a211oi_2
X_17841_ _08351_ _08352_ vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__nand2_1
X_14984_ _03321_ _06094_ _00460_ _03322_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__a22oi_1
X_17772_ _08176_ _08177_ _08175_ vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__o21ai_1
X_13935_ _04101_ _04102_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__nand2_1
X_16723_ _07031_ _07044_ _07135_ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16654_ _06967_ _06975_ _07060_ vssd1 vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__o21ai_1
X_13866_ _03863_ _03871_ _04027_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__a21bo_1
X_15605_ _05915_ _05923_ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__and2_1
X_12817_ _02907_ _02908_ _01468_ _01490_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16585_ _06984_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__xor2_1
X_13797_ _05975_ _03763_ _03765_ _03766_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15536_ _07668_ _00318_ _05758_ _03009_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__a22o_1
X_18324_ _02887_ _08877_ vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _02838_ _02840_ _02837_ vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__a21o_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18255_ _08802_ _08803_ vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__and2_1
X_15467_ _05773_ _05757_ _05759_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ _02769_ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__and2_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17206_ _07538_ _07545_ _07536_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__o21ba_1
X_14418_ _01504_ _05856_ _04497_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__and3_1
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18186_ _08727_ _08728_ vssd1 vssd1 vccd1 vccd1 _08729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_396 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15398_ _05596_ _05699_ vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17137_ _07549_ _07551_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__and2b_1
X_14349_ _04552_ _04554_ _04555_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17068_ _04012_ _06889_ vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__nand2_4
XFILLER_0_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16019_ _06367_ _06369_ _00786_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__a21bo_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _06949_ _08278_ _08289_ _08300_ vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__or4b_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10030_ _08191_ _00122_ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11981_ _01967_ _02027_ _02052_ vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__or3_1
X_13720_ cla_inst.in2\[25\] _04012_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2_1
X_10932_ _03771_ _04242_ _00176_ _04078_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13651_ _06040_ _06084_ _00509_ _00513_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10863_ _04078_ _03771_ _00949_ _03421_ vssd1 vssd1 vccd1 vccd1 _00956_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12602_ _02654_ _02660_ _02661_ vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__a21oi_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ net212 _06517_ _06520_ _06751_ vssd1 vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _03676_ _03677_ _03715_ _03716_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__o211a_1
X_10794_ _00868_ _00886_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15321_ _05520_ _05516_ _05517_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12533_ _02622_ _02624_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__nand2_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18040_ _08568_ _08569_ vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__nand2_1
X_15252_ _05538_ _01139_ _05449_ _05539_ vssd1 vssd1 vccd1 vccd1 _05541_ sky130_fd_sc_hd__and4b_1
XFILLER_0_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12464_ _02550_ _02556_ vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ _04393_ _04394_ _04396_ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__or3_4
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _03662_ _07591_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__nand2_2
XFILLER_0_124_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15183_ _09350_ _05715_ _05975_ _00112_ vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__a22oi_1
X_12395_ _05671_ _00197_ _02486_ _02487_ _09188_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ _00678_ _04045_ _04067_ _00679_ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__a22o_1
X_11346_ _01413_ _01414_ _01312_ _01378_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18942_ clknet_4_2_0_clk _00096_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[28\] sky130_fd_sc_hd__dfxtp_1
X_14065_ _03540_ _03554_ _02980_ vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__mux2_1
X_11277_ _01238_ _01273_ _01368_ _01369_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__o211a_1
X_13016_ _03025_ _03108_ _02272_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a21o_1
X_10228_ _05747_ _07025_ _00317_ _00320_ vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__and4_1
X_18873_ clknet_4_14_0_clk net246 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__dfxtp_1
X_17824_ _06388_ _06387_ _06386_ vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__a21o_1
X_10159_ _00203_ _00166_ vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14967_ _00678_ _00443_ _06471_ _00679_ vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__a22o_1
X_17755_ _07933_ vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__buf_2
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16706_ _06766_ _06875_ _07114_ _07116_ vssd1 vssd1 vccd1 vccd1 _07117_ sky130_fd_sc_hd__nor4_1
X_13918_ _04080_ _04084_ _03921_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__mux2_1
X_17686_ _08183_ _08184_ vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__or2b_1
X_14898_ _05009_ _05154_ vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _00173_ _00175_ _04460_ _04482_ vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__and4_2
X_16637_ _06957_ vssd1 vssd1 vccd1 vccd1 _07042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16568_ _06939_ _06966_ vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18307_ _08858_ _08844_ vssd1 vssd1 vccd1 vccd1 _08860_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15519_ _05746_ _05745_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__or2b_1
X_16499_ _06801_ _06818_ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18238_ _08707_ _08710_ _08783_ vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18169_ _08704_ _08708_ vssd1 vssd1 vccd1 vccd1 _08710_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap121 _03884_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_1
XFILLER_0_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap143 _00603_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_1
X_09942_ _07123_ vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _07319_ _07940_ _08115_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__nand3_4
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _00968_ _00973_ vssd1 vssd1 vccd1 vccd1 _01293_ sky130_fd_sc_hd__nand2_1
X_12180_ _00846_ _00716_ _02272_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _00515_ _01136_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__nor2_4
XFILLER_0_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ _04984_ _00218_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__nand2_1
X_10013_ cla_inst.in2\[25\] vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__clkbuf_4
X_15870_ _06209_ _06210_ vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14821_ _04896_ _04963_ _05069_ _05070_ vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14752_ _04725_ _04125_ _04994_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__and3_2
X_17540_ _07911_ _07912_ _07910_ vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__a21o_1
X_11964_ _02006_ _02001_ _02004_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13703_ _03847_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__nand2_1
X_10915_ _05671_ _05322_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17471_ _07942_ _07949_ vssd1 vssd1 vccd1 vccd1 _07950_ sky130_fd_sc_hd__xor2_1
X_14683_ _04917_ _04918_ _04903_ _04791_ vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__o211ai_1
X_11895_ _01675_ _01864_ _01981_ vssd1 vssd1 vccd1 vccd1 _01988_ sky130_fd_sc_hd__or3_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13634_ _03612_ _03613_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__nand2_2
X_16422_ _07657_ _06541_ _06807_ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__and3_1
X_10846_ _00932_ _00933_ _00937_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__nand3_1
XFILLER_0_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16353_ _06727_ _06733_ _03079_ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__mux2_2
X_13565_ _03496_ _03502_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__nand2_1
Xsplit84 _06571_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlymetal6s2s_1
X_10777_ _00200_ _00869_ vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15304_ _05552_ _05596_ _05597_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12516_ _02608_ _02559_ vssd1 vssd1 vccd1 vccd1 _02609_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16284_ _06654_ _06658_ vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__and2_1
X_13496_ _03620_ _03621_ _03393_ _03587_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a211o_4
XFILLER_0_136_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15235_ _05518_ _05521_ _05522_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__a21o_1
X_18023_ _07194_ _07290_ _07511_ _07621_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__or4_1
X_12447_ _02538_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15166_ _05445_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__nor2_1
X_12378_ _02400_ _02461_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__xor2_2
X_14117_ _04115_ _04109_ vssd1 vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__and2b_1
X_11329_ cla_inst.in2\[20\] _00878_ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15097_ _01505_ _00322_ vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14048_ _04052_ _04055_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__or2b_1
X_18925_ clknet_4_11_0_clk _00079_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_4
X_18856_ clknet_4_4_0_clk net256 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__dfxtp_1
X_17807_ _08187_ _08200_ _08198_ vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__a21o_1
X_18787_ _02985_ net45 _09276_ vssd1 vssd1 vccd1 vccd1 _09299_ sky130_fd_sc_hd__mux2_1
X_15999_ _07058_ _01264_ vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17738_ _06385_ _06546_ _08241_ _01678_ vssd1 vssd1 vccd1 vccd1 _08242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17669_ _08159_ _08164_ vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09925_ _06384_ _06439_ vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__or2b_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _07210_ _07308_ _07297_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__a21o_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _05736_ _05986_ _06105_ _06073_ vssd1 vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__a31o_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _09403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_116 _00131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _03790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _05888_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 _08762_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _00762_ _00763_ _00778_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__a21o_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ cla_inst.in2\[20\] _01503_ _01240_ _01506_ vssd1 vssd1 vccd1 vccd1 _01773_
+ sky130_fd_sc_hd__a22o_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10631_ _09353_ _00207_ _00548_ _00547_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__a31o_1
X_13350_ _03449_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__xnor2_1
X_10562_ _00638_ _00653_ _00654_ vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12301_ _02390_ _02391_ _02385_ net123 vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_133_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _03728_ _06062_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10493_ _00583_ _00584_ net339 _00424_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15020_ _05243_ _05287_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__xor2_2
XFILLER_0_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12232_ _02323_ _02324_ vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12163_ _02254_ _02255_ vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11114_ _07254_ _05039_ _00439_ _07232_ vssd1 vssd1 vccd1 vccd1 _01207_ sky130_fd_sc_hd__a22o_1
X_12094_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__nand2_1
X_16971_ _07392_ _07404_ vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__xnor2_1
X_18710_ net54 _03068_ _09182_ vssd1 vssd1 vccd1 vccd1 _09238_ sky130_fd_sc_hd__mux2_1
X_11045_ _01109_ _01137_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__nand2_1
X_15922_ _04958_ _05307_ _06266_ _03039_ vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__o22a_1
X_18641_ _09187_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__clkbuf_1
X_15853_ _06118_ _06173_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__and2b_1
X_14804_ _05051_ _05052_ vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nand2_1
X_18572_ salida\[8\] _09114_ _09118_ salida\[40\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09138_ sky130_fd_sc_hd__a221o_1
X_15784_ _06098_ _06099_ _06117_ vssd1 vssd1 vccd1 vccd1 _06119_ sky130_fd_sc_hd__or3_1
X_12996_ _03047_ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__clkbuf_4
X_17523_ _07999_ _08007_ vssd1 vssd1 vccd1 vccd1 _08008_ sky130_fd_sc_hd__xnor2_1
X_14735_ _04034_ _00502_ _09311_ _04099_ vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_52_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11947_ _02035_ _02038_ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17454_ _07896_ _07898_ vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__nor2_1
X_14666_ _04899_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11878_ _01969_ _01938_ _01970_ _01869_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13617_ _03366_ cla_inst.in1\[20\] _05377_ _03345_ vssd1 vssd1 vccd1 vccd1 _03755_
+ sky130_fd_sc_hd__a22o_1
X_16405_ _03083_ _06430_ vssd1 vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__nor2_1
X_10829_ _00920_ _00921_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__and2b_1
X_14597_ _03543_ _03555_ _02979_ vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__mux2_1
X_17385_ _07727_ _07719_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__and2b_1
X_13548_ _03678_ _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__nor2_1
X_16336_ _03077_ _06715_ vssd1 vssd1 vccd1 vccd1 _06716_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16267_ _06467_ _06640_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__and2_1
X_13479_ net330 _03597_ _03602_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__a21o_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15218_ _05429_ _05390_ _05502_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__or3_1
X_18006_ _07313_ _07487_ _07593_ _07318_ vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__o22a_1
XFILLER_0_140_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16198_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel _03826_ sel_op\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__or3b_1
X_15149_ _05390_ _05391_ _05394_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__or3_1
X_09710_ _06267_ _06329_ _06319_ vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__a21o_1
X_18908_ clknet_4_10_0_clk _00062_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[26\] sky130_fd_sc_hd__dfxtp_1
X_09641_ cla_inst.in1\[22\] vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__buf_4
X_18839_ clknet_4_0_0_clk net302 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__dfxtp_1
X_09572_ _03990_ _04482_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__nand2_8
XFILLER_0_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09908_ _08398_ _08485_ _08474_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__a21o_1
X_09839_ cla_inst.in1\[29\] vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__clkbuf_4
X_12850_ _00893_ _00895_ _00897_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__and3_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _01707_ _01891_ _01887_ _01890_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__o211a_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _01370_ _01373_ _01371_ _01372_ vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__o211a_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer80 _04683_ vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer91 _00375_ vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__clkbuf_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _04739_ _04740_ _04598_ _04701_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__o211ai_4
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _01816_ _01819_ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__xnor2_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _04650_ _04525_ _04666_ vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__a21oi_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11663_ _01741_ _01754_ _01755_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__nand3_2
XFILLER_0_37_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13402_ _03337_ _03339_ _03518_ _03519_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10614_ _00705_ _00706_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__xnor2_2
X_17170_ _06561_ _07124_ _07318_ _07621_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__or4_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14382_ _06460_ _03455_ vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__nand2_1
X_11594_ _01684_ _01685_ _01686_ vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__nand3_2
XFILLER_0_36_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16121_ _04241_ _06474_ _06480_ _03117_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ _00362_ _00207_ _03441_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_24_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ _00457_ _00462_ _00456_ vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _06404_ _06405_ vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13264_ _03368_ _03311_ _03310_ vssd1 vssd1 vccd1 vccd1 _03369_ sky130_fd_sc_hd__nand3_2
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10476_ _00253_ _00166_ _00406_ _00405_ vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15003_ _05267_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12215_ _02295_ _02299_ _02306_ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__o211a_1
X_13195_ _03293_ _03294_ _00661_ net327 vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__a211o_4
X_12146_ _02235_ _02238_ vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12077_ _02081_ _02167_ _02169_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__o21ai_1
X_16954_ _06374_ _03324_ _06814_ _07386_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__a211o_2
X_11028_ _01097_ _01101_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__xnor2_1
X_15905_ _03013_ _06246_ _06248_ vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__and3_1
X_16885_ _02124_ _06871_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ salida\[29\] _09159_ _09160_ salida\[61\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09174_ sky130_fd_sc_hd__a221o_1
X_15836_ _06161_ _06174_ vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18555_ net295 _09098_ _09122_ _09126_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__o211a_1
X_12979_ _03071_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__clkbuf_4
X_15767_ _02992_ _03071_ _06037_ _06041_ vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17506_ _07987_ _07988_ vssd1 vssd1 vccd1 vccd1 _07989_ sky130_fd_sc_hd__nor2_1
X_14718_ _04957_ _04958_ _03538_ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18486_ _03155_ _08428_ _03011_ vssd1 vssd1 vccd1 vccd1 _09053_ sky130_fd_sc_hd__or3b_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15698_ _03012_ _09059_ _00322_ _03010_ vssd1 vssd1 vccd1 vccd1 _06025_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17437_ _07911_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__inv_2
X_14649_ _04880_ _04881_ net196 _04756_ vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_27 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_49 _03265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17368_ _07836_ _07837_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16319_ _02489_ _03152_ _06487_ _06485_ vssd1 vssd1 vccd1 vccd1 _06697_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17299_ _07739_ _07740_ _07761_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput101 net101 vssd1 vssd1 vccd1 vccd1 o_wb_data[26] sky130_fd_sc_hd__clkbuf_4
Xoutput112 net112 vssd1 vssd1 vccd1 vccd1 o_wb_data[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09624_ _05366_ _05322_ _05388_ _05410_ vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09555_ _04646_ _04373_ _04395_ _04657_ vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__and4_4
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ _03826_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__buf_6
XFILLER_0_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10330_ net338 _00377_ _09346_ _00274_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10261_ cla_inst.in2\[31\] _07613_ _00351_ _00352_ vssd1 vssd1 vccd1 vccd1 _00354_
+ sky130_fd_sc_hd__a22oi_1
X_12000_ _05224_ _00178_ vssd1 vssd1 vccd1 vccd1 _02093_ sky130_fd_sc_hd__nand2_2
X_10192_ _03990_ _05497_ vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _04107_ _04108_ _04119_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__o21ai_2
X_12902_ _02992_ _01417_ _01359_ _02994_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__or4_1
X_13882_ _03828_ _04007_ _04043_ _04044_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__a211oi_2
X_16670_ _06341_ _06546_ _07077_ _00881_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__a22o_1
X_12833_ _02923_ _02907_ _02924_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__o211ai_4
X_15621_ _05841_ _05940_ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__or2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _06374_ _06368_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15552_ _05866_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__inv_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _01238_ _01272_ _01271_ vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__o21ai_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _04719_ _04720_ _04721_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11715_ _01507_ _01806_ _01807_ vssd1 vssd1 vccd1 vccd1 _01808_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15483_ _05792_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__inv_2
X_18271_ _05557_ _06400_ _06401_ vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__and3_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12695_ _02755_ _02785_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__or2_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17222_ _04725_ _06510_ _02127_ vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14434_ _04645_ _04648_ vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__xor2_4
X_11646_ _01721_ _01737_ _01738_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__nand3_4
XFILLER_0_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 i_wb_addr[20] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 i_wb_addr[30] vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14365_ _04567_ net181 _04571_ _04572_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__o211ai_4
X_17153_ _07396_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 i_wb_data[10] vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_2
X_11577_ _01655_ _01668_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput47 i_wb_data[20] vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__clkbuf_2
X_13316_ _03411_ _03424_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and3_2
Xinput58 i_wb_data[30] vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_1
XFILLER_0_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16104_ _06462_ vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__buf_4
Xinput69 reset vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__buf_4
X_10528_ _00617_ _00618_ _00619_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__a21oi_2
X_17084_ _07518_ _07528_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__xnor2_1
X_14296_ _01504_ _05856_ vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ _03349_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16035_ _02985_ _01695_ vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__nand2_1
X_10459_ _00544_ _00551_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13178_ _03269_ _03275_ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__nand2_1
X_12129_ _02185_ _02186_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__or2_1
X_17986_ _03000_ _06511_ _00813_ vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16937_ _06360_ _06545_ _07368_ _03101_ vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__a22o_1
X_16868_ _06657_ _07108_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__nand2_1
X_18607_ _09127_ vssd1 vssd1 vccd1 vccd1 _09163_ sky130_fd_sc_hd__clkbuf_4
X_15819_ _06155_ vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__inv_2
X_16799_ _03324_ _06529_ _06814_ _02099_ vssd1 vssd1 vccd1 vccd1 _07218_ sky130_fd_sc_hd__a211o_2
XFILLER_0_90_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18538_ _09099_ _09100_ _09102_ _09107_ vssd1 vssd1 vccd1 vccd1 _09108_ sky130_fd_sc_hd__nor4_2
XFILLER_0_74_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18469_ _07256_ _09022_ _09025_ _09034_ vssd1 vssd1 vccd1 vccd1 _09035_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _05224_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__buf_4
X_09538_ _04471_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__buf_12
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ _03717_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _01589_ _01592_ vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ _02572_ vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11431_ _01518_ _01523_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14150_ _04181_ _04180_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__or2b_1
X_11362_ _01401_ _01403_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__or2b_1
X_13101_ _03165_ _03193_ _02975_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10313_ _00183_ _03432_ _03618_ _00184_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14081_ _03568_ _03571_ _03099_ vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11293_ _00811_ _00815_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__xnor2_1
X_13032_ _06765_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__nor2_2
X_10244_ _09080_ _09131_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17840_ _07035_ _07125_ _07487_ _07593_ vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__or4_2
X_10175_ _07919_ _08289_ _00266_ _00267_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__o211a_2
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17771_ _08275_ _08276_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__nor2_1
X_14983_ _07635_ _05888_ _05127_ _05125_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__a31o_1
X_16722_ _06945_ _07030_ vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or2b_1
X_13934_ _04099_ _04132_ _07962_ _05715_ vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__nand4_1
XFILLER_0_88_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16653_ _06939_ _06966_ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__nand2_1
X_13865_ _03864_ _03869_ vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__nand2_1
X_15604_ _05915_ _05923_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__nor2_1
X_12816_ _01468_ _01490_ _02907_ _02908_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a211oi_2
X_16584_ _06866_ _06900_ _06902_ vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__a21bo_1
X_13796_ _03777_ _03778_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18323_ _02887_ _08877_ vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__or2_1
XFILLER_0_139_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15535_ _03009_ _07668_ _01317_ _05758_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__and4_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12747_ _02746_ _02750_ vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__or2b_1
XFILLER_0_45_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18254_ _08798_ _08801_ vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15466_ _05757_ _05759_ _05773_ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__a21oi_1
X_12678_ _02762_ _02770_ vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17205_ _07648_ _07660_ vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__xnor2_1
X_11629_ _01215_ _01209_ _01214_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__nand3_2
X_14417_ _00877_ _03044_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18185_ _08632_ _08649_ _08633_ vssd1 vssd1 vccd1 vccd1 _08728_ sky130_fd_sc_hd__o21ba_1
X_15397_ _05697_ _05698_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17136_ _07561_ _07564_ _07585_ _06723_ _02259_ vssd1 vssd1 vccd1 vccd1 _09389_ sky130_fd_sc_hd__o32a_2
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14348_ _04552_ _04554_ _03202_ vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14279_ _03014_ _00716_ _04476_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a22oi_1
X_17067_ _07401_ _07403_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16018_ _04725_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__or2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _08486_ _08492_ vssd1 vssd1 vccd1 vccd1 _08493_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11980_ _02067_ _02070_ net130 _02072_ vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__a211oi_4
X_10931_ _04078_ _03771_ _04242_ _00772_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13650_ _06084_ _03455_ _00513_ _03790_ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a22oi_1
X_10862_ net194 _00953_ _00954_ vssd1 vssd1 vccd1 vccd1 _00955_ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12601_ _02650_ net203 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__or2b_1
X_13581_ _03713_ _03714_ _03696_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__o21ai_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _00884_ _00885_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__nor2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15320_ _05516_ _05517_ _05407_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__and3b_1
X_12532_ _02622_ _02624_ vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__xnor2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15251_ _07668_ _01223_ _00461_ _03009_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a22o_1
X_12463_ _02550_ _02554_ _02555_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14202_ _04188_ _04190_ _04186_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_50_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11414_ cla_inst.in2\[20\] _01503_ _01240_ _01506_ vssd1 vssd1 vccd1 vccd1 _01507_
+ sky130_fd_sc_hd__and4_2
X_15182_ _07635_ _00461_ _05334_ _05332_ vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12394_ _06019_ _08039_ _09212_ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14133_ _00679_ _00678_ _04045_ _04154_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__and4_1
X_11345_ _01362_ _01437_ vssd1 vssd1 vccd1 vccd1 _01438_ sky130_fd_sc_hd__xnor2_1
X_18941_ clknet_4_2_0_clk _00095_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[27\] sky130_fd_sc_hd__dfxtp_2
X_14064_ _03550_ _03552_ _03099_ vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__mux2_1
X_11276_ _01337_ _01367_ _01366_ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__o21ai_1
X_13015_ _03107_ vssd1 vssd1 vccd1 vccd1 _03108_ sky130_fd_sc_hd__buf_4
X_10227_ _00318_ _00319_ vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__nand2_1
X_18872_ clknet_4_14_0_clk net305 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__dfxtp_1
X_17823_ _06388_ _06386_ _06387_ vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__nand3_1
X_10158_ _00204_ _00214_ _00225_ vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17754_ _08155_ _08157_ vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__and2b_1
X_14966_ _03005_ _05921_ vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10089_ _00173_ _00175_ _00178_ _00181_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__nand4_1
X_16705_ _06653_ _06944_ _07115_ _06571_ vssd1 vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13917_ _04082_ _04083_ _02780_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__mux2_1
X_17685_ _08063_ _08149_ _08182_ vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14897_ _05143_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__xor2_1
X_16636_ _07037_ _07040_ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__nand2_1
X_13848_ _00702_ _04700_ _08409_ _00195_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16567_ _06940_ _06965_ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__xor2_1
X_13779_ _03509_ _08746_ _08049_ _03531_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18306_ _08844_ _08858_ vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__and2b_1
X_15518_ _05828_ _05829_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16498_ _06890_ vssd1 vssd1 vccd1 vccd1 _06891_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18237_ _08707_ _08710_ _08783_ vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__nand3_1
X_15449_ _05739_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18168_ _08704_ _08708_ vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17119_ _07462_ _07463_ _07460_ vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__o21bai_2
Xmax_cap122 _02521_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap144 _01178_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_1
X_18099_ _08632_ _08633_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _05736_ vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09872_ _08017_ _08093_ _08104_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__a21o_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _06094_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__buf_4
XFILLER_0_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11061_ _01152_ _01153_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__and2b_1
X_10012_ _09351_ _09353_ _07646_ _09354_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__and4_1
X_14820_ _05067_ _05068_ _04932_ _04964_ vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__a211o_2
XFILLER_0_99_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14751_ _04856_ _04855_ vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__nand2_1
X_11963_ _01941_ _02055_ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__nand2_1
X_13702_ _03845_ _03846_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__nand2_1
X_10914_ _01004_ _01006_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17470_ _07947_ _07948_ vssd1 vssd1 vccd1 vccd1 _07949_ sky130_fd_sc_hd__or2_1
X_14682_ _04903_ _04791_ _04917_ _04918_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11894_ _01980_ _01984_ _01986_ vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16421_ _06802_ _06806_ _03535_ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__a21oi_2
X_13633_ _03768_ _03769_ _03770_ vssd1 vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__a21oi_2
X_10845_ _00932_ _00933_ _00937_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xsplit74 _06560_ vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlymetal6s2s_1
X_16352_ _06729_ _06731_ _03098_ vssd1 vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__mux2_1
X_13564_ _03494_ _03505_ vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__nand2_1
X_10776_ _00253_ _00194_ _00198_ _00199_ vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15303_ _05593_ _05594_ _05478_ _05553_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12515_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel _00218_ _02607_
+ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__and3_1
X_13495_ _03393_ net134 _03620_ _03621_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__o211ai_4
X_16283_ _06572_ _06581_ _06657_ _06527_ vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_136_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18022_ _07396_ _07780_ _07623_ _07394_ vssd1 vssd1 vccd1 vccd1 _08551_ sky130_fd_sc_hd__a22o_1
X_15234_ _05518_ _05521_ _03930_ vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__o21ai_1
X_12446_ _02475_ _02478_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15165_ _03008_ _07515_ _00460_ _05856_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__and4_1
XFILLER_0_23_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12377_ _02176_ _02469_ vssd1 vssd1 vccd1 vccd1 _02470_ sky130_fd_sc_hd__and2_4
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14116_ _04137_ _04136_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__and2b_1
X_11328_ _01358_ _01420_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__xor2_1
X_15096_ _05369_ _05370_ vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18924_ clknet_4_11_0_clk _00078_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_14047_ _04222_ _04223_ _04224_ vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__o21ai_1
X_11259_ _01350_ _01339_ _01340_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__nor3_1
X_18855_ clknet_4_7_0_clk net276 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__dfxtp_1
X_17806_ _08314_ _08315_ vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__and2_1
X_18786_ _09125_ vssd1 vssd1 vccd1 vccd1 _09298_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15998_ _06343_ _06344_ _06345_ _06346_ vssd1 vssd1 vccd1 vccd1 _06347_ sky130_fd_sc_hd__and4_1
X_17737_ _02987_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__a21o_1
X_14949_ _02989_ _03456_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ _08159_ _08164_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16619_ _06567_ _06570_ _06946_ _00357_ vssd1 vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__o211a_1
X_17599_ _08088_ _08089_ vssd1 vssd1 vccd1 vccd1 _08090_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09924_ _06373_ _08322_ _08659_ _08670_ vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__a211o_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _07908_ _07897_ _06960_ _05812_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__a211oi_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _06993_ _07025_ _07145_ _07167_ vssd1 vssd1 vccd1 vccd1 _07178_ sky130_fd_sc_hd__nand4_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 op_code\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_117 _00166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_128 _04034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_139 _06765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ _00512_ _00518_ vssd1 vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10561_ _00651_ _00652_ _00643_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12300_ _02258_ _02260_ _02386_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13280_ _00459_ _03384_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10492_ net339 _00424_ _00583_ _00584_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__o211a_4
XFILLER_0_134_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12231_ _02313_ _02318_ _02317_ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12162_ _02240_ _02253_ vssd1 vssd1 vccd1 vccd1 _02255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11113_ _07047_ _07254_ _05497_ _04580_ vssd1 vssd1 vccd1 vccd1 _01206_ sky130_fd_sc_hd__nand4_2
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12093_ _02177_ _02182_ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__xor2_1
X_16970_ _07401_ _07403_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__xor2_1
X_11044_ _01105_ _00514_ _01136_ _00813_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__or4_4
X_15921_ _04955_ _04957_ _03536_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18640_ _09176_ _09186_ vssd1 vssd1 vccd1 vccd1 _09187_ sky130_fd_sc_hd__and2_1
X_15852_ _06183_ _06187_ _06190_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__o21ai_1
X_14803_ _05036_ _05037_ _05049_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__nand3_1
X_18571_ net273 _09098_ _09136_ _09126_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__o211a_1
X_15783_ _06098_ _06099_ _06117_ vssd1 vssd1 vccd1 vccd1 _06118_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12995_ _03023_ _03087_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__nand2_1
X_17522_ _08004_ _08005_ vssd1 vssd1 vccd1 vccd1 _08007_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14734_ _04972_ _04974_ _04838_ _04839_ vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__o211ai_2
X_11946_ _02035_ _02038_ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17453_ _07891_ _07892_ _07895_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__and3_1
X_14665_ _00164_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__nand2_2
X_11877_ _01865_ _01867_ _01868_ _01861_ vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__o31ai_2
X_16404_ _06544_ vssd1 vssd1 vccd1 vccd1 _06790_ sky130_fd_sc_hd__clkbuf_4
X_13616_ _03588_ _03589_ _03590_ vssd1 vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__nor3_2
X_17384_ _07726_ _07720_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__and2b_1
X_10828_ _03771_ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel _04220_
+ cla_inst.in2\[16\] vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__a22o_1
X_14596_ _02979_ _03551_ _04825_ vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16335_ _03050_ _02563_ _03173_ _06470_ _06714_ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__o311a_1
X_13547_ cla_inst.in2\[24\] _00174_ _04886_ _03903_ vssd1 vssd1 vccd1 vccd1 _03679_
+ sky130_fd_sc_hd__and4_1
X_10759_ _00829_ _00851_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16266_ _00167_ _03101_ _00593_ _00558_ _03028_ _02982_ vssd1 vssd1 vccd1 vccd1 _06640_
+ sky130_fd_sc_hd__mux4_1
X_13478_ _03595_ _03597_ _03602_ vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__nand3_1
XFILLER_0_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18005_ _07039_ _07708_ _08460_ _08357_ vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__a31o_1
X_15217_ _05429_ _05390_ _05502_ vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_140_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12429_ _02450_ _02455_ _02454_ vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__o21ai_1
X_16197_ _03281_ _06529_ _06520_ vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15148_ _05402_ _05403_ vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15079_ _09350_ _05964_ _06094_ _00112_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a22oi_1
X_18907_ clknet_4_10_0_clk _00061_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[25\] sky130_fd_sc_hd__dfxtp_1
X_09640_ _05584_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__clkbuf_4
X_18838_ clknet_4_0_0_clk net296 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09571_ _04810_ _04821_ _04831_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__nand3_1
X_18769_ _09273_ _09284_ vssd1 vssd1 vccd1 vccd1 _09285_ sky130_fd_sc_hd__and2_1
XFILLER_0_148_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09907_ _08398_ _08474_ _08485_ vssd1 vssd1 vccd1 vccd1 _08496_ sky130_fd_sc_hd__nand3_1
X_09838_ _07733_ vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__buf_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _06982_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__clkbuf_8
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _01872_ _01875_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__xnor2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _00591_ _01264_ _01263_ _01261_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__a31o_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer70 _00694_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlymetal6s4s_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer81 net243 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer92 _00378_ vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _01821_ _01822_ _01823_ vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__o21ba_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14450_ _04664_ _04665_ vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nand2_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _01739_ _01740_ _01642_ net125 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13401_ _03516_ _03517_ _03371_ _03372_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__a211oi_2
X_10613_ _00253_ _00398_ vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14381_ _04515_ _04588_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a21bo_1
X_11593_ _01208_ _01683_ _01682_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a21o_1
X_16120_ _03164_ _06476_ _06479_ _03547_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13332_ _03440_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ _00476_ _00480_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16051_ _02992_ _03068_ vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__or2_1
X_10475_ _00566_ _00567_ vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__xnor2_1
X_13263_ _00592_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__buf_4
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15002_ _01504_ _08876_ vssd1 vssd1 vccd1 vccd1 _05269_ sky130_fd_sc_hd__nand2_1
X_12214_ _02302_ _02305_ _02304_ vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__o21ai_1
X_13194_ _00661_ net327 _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _02236_ _02237_ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12076_ _02168_ _01991_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__xnor2_1
X_16953_ _06460_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__inv_2
X_11027_ _01118_ _01119_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__nor2_1
X_15904_ _06247_ vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__buf_2
X_16884_ _01962_ _06812_ _06871_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__o21ai_4
X_18623_ net308 _09157_ _09173_ _09162_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835_ _06118_ _06173_ vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18554_ _09125_ vssd1 vssd1 vccd1 vccd1 _09126_ sky130_fd_sc_hd__buf_2
X_15766_ _06047_ _06046_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2b_1
X_12978_ _00495_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__clkbuf_4
X_17505_ _07985_ _07986_ vssd1 vssd1 vccd1 vccd1 _07988_ sky130_fd_sc_hd__nor2_1
X_14717_ _03547_ _03572_ vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18485_ _03011_ _06512_ _03155_ vssd1 vssd1 vccd1 vccd1 _09052_ sky130_fd_sc_hd__a21bo_1
X_11929_ _02007_ _02008_ vssd1 vssd1 vccd1 vccd1 _02022_ sky130_fd_sc_hd__xor2_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15697_ _03015_ _00339_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__and2_2
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17436_ _07910_ _07911_ _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__and3b_1
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14648_ _04741_ _04756_ _04880_ _04881_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 _01697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ _07018_ _07387_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__nor2_1
X_14579_ _04805_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__nor2_2
XFILLER_0_28_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16318_ _02982_ _06490_ _06695_ _06626_ vssd1 vssd1 vccd1 vccd1 _06696_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17298_ _07739_ _07740_ _07761_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16249_ _06470_ _06620_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__nand2_1
Xoutput102 net102 vssd1 vssd1 vccd1 vccd1 o_wb_data[27] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput113 net113 vssd1 vssd1 vccd1 vccd1 o_wb_data[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _05399_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__buf_4
X_09554_ _03739_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09485_ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03903_ sky130_fd_sc_hd__buf_4
XFILLER_0_66_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ cla_inst.in2\[31\] _07613_ _00351_ _00352_ vssd1 vssd1 vccd1 vccd1 _00353_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10191_ _00282_ _00283_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__nor2_1
X_13950_ _04117_ _04118_ vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__or2_1
X_12901_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__buf_2
X_13881_ _04041_ _04042_ _04024_ vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _05841_ _05940_ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__nand2_1
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _00856_ _00890_ _00889_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__o21ai_2
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _05776_ _05778_ _05864_ _05865_ vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__o211a_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _01238_ _01271_ _01272_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _04719_ _04720_ _04721_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__and3_2
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11714_ _01804_ _01805_ _01784_ _01787_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__a211o_1
X_18270_ _02881_ _08819_ vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__xnor2_4
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _05615_ _05790_ vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _02505_ _00134_ _00108_ _00845_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a22o_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17221_ _02633_ _07676_ _07677_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__a21oi_2
X_14433_ _01873_ _04647_ vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__nand2_2
XFILLER_0_126_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11645_ _01719_ _01720_ _01621_ _01640_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17152_ _07589_ _07601_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__xnor2_1
Xinput15 i_wb_addr[21] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
X_14364_ _02986_ _06732_ _04568_ _04570_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput26 i_wb_addr[31] vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11576_ _01655_ _01668_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__or2_1
Xinput37 i_wb_data[11] vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_2
XFILLER_0_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput48 i_wb_data[21] vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_2
X_16103_ _06461_ vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__clkbuf_4
X_13315_ _03422_ _03423_ _03416_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a21o_1
Xinput59 i_wb_data[31] vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_2
X_10527_ _00617_ _00618_ _00619_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__and3_4
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17083_ _07525_ _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ _04495_ _04496_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nor2_1
X_16034_ _02985_ _01695_ vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__or2_2
X_13246_ _03347_ _03348_ _00747_ _03203_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__a211o_1
X_10458_ _00545_ _00550_ vssd1 vssd1 vccd1 vccd1 _00551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10389_ _00468_ _00469_ _00481_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a21o_2
X_13177_ _03269_ _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12128_ _02218_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__nand2_1
X_17985_ _02167_ _02174_ _08424_ _08510_ _03202_ vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__o311a_2
X_16936_ _00644_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _07368_ sky130_fd_sc_hd__a21o_1
X_12059_ _02151_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__inv_2
X_16867_ _07288_ _07291_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__xor2_2
X_15818_ _03010_ _03012_ _03071_ _03149_ vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and4_1
X_18606_ net279 _09157_ _09161_ _09162_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _07038_ _06969_ _07216_ _06527_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__a22o_1
X_18537_ _09103_ _09104_ _09105_ _09106_ vssd1 vssd1 vccd1 vccd1 _09107_ sky130_fd_sc_hd__or4_2
X_15749_ _06074_ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18468_ _06412_ _06421_ _09026_ _09033_ vssd1 vssd1 vccd1 vccd1 _09034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17419_ _07767_ _07768_ _07770_ vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__or3_1
X_18399_ _04406_ _07592_ _08957_ vssd1 vssd1 vccd1 vccd1 _08959_ sky130_fd_sc_hd__a21o_1
XFILLER_0_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _05213_ vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09537_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04471_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09468_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03717_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11430_ _01519_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _01415_ _01438_ _01439_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__nor3_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10312_ _00184_ _00183_ _03432_ _00205_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__and4_1
X_13100_ _03178_ _03192_ _02780_ vssd1 vssd1 vccd1 vccd1 _03193_ sky130_fd_sc_hd__mux2_1
X_11292_ _01281_ _01282_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__or2b_1
X_14080_ _04247_ _04258_ _04260_ vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__o21ai_1
X_10243_ _08681_ _09005_ _00333_ _00335_ vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_30_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ _02728_ _02965_ _03239_ _03217_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__or4b_4
X_10174_ _00245_ _00246_ _00265_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__nand3_2
X_17770_ _08259_ _08166_ _08274_ vssd1 vssd1 vccd1 vccd1 _08276_ sky130_fd_sc_hd__nor3_1
X_14982_ _05146_ _05149_ vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nand2_1
X_16721_ _07122_ _07132_ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__xnor2_1
X_13933_ _04132_ _07962_ _00308_ _04099_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16652_ _07049_ _07057_ vssd1 vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__xnor2_1
X_13864_ _03861_ _03873_ vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__nand2_1
X_15603_ _05920_ _05922_ vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__or2_1
X_12815_ _02899_ _02906_ _02905_ vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__a21oi_1
X_16583_ _06981_ _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or2b_1
X_13795_ _03945_ _03947_ _03948_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18322_ _08875_ _08759_ _02893_ vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__o21a_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ _03006_ _04647_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__nand2_1
X_12746_ _02837_ _02838_ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _08798_ _08801_ vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__nand2_1
X_15465_ _05771_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12677_ _02753_ _02761_ vssd1 vssd1 vccd1 vccd1 _02770_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17204_ _07658_ _07659_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__nor2_1
X_14416_ _04626_ _04627_ _04470_ _04488_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _01621_ _01640_ _01719_ _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_108_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18184_ _08725_ _08726_ vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__nor2_1
X_15396_ _05549_ _05598_ _05696_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17135_ _07256_ _07568_ _07569_ _07584_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__a31o_1
X_14347_ _04401_ _04410_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ _01649_ _01650_ _01651_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__and3_1
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17066_ _07415_ _07423_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__nor2_1
X_14278_ _04475_ vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _00716_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__clkbuf_4
X_13229_ _03317_ _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__xnor2_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _08490_ _08491_ vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__nor2_1
X_16919_ _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__and2_4
X_17899_ _08120_ _08219_ _08414_ _08416_ _08325_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__o311a_1
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ _00939_ _00938_ _00931_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__a21o_1
X_10861_ _00925_ _00926_ _00940_ vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _02672_ _02673_ _02692_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__and3_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _03696_ _03713_ _03714_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__or3_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10792_ _00883_ _00876_ _00880_ vssd1 vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__nor3_1
XFILLER_0_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12531_ _02567_ _02623_ vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__xnor2_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _03009_ _07668_ _01223_ _00461_ vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and4_1
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12462_ _02545_ _02549_ _02548_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14201_ _04390_ _04391_ _04392_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11413_ _00877_ _07646_ _09354_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15181_ _05353_ _05354_ vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12393_ _08039_ _00871_ _07548_ _06019_ vssd1 vssd1 vccd1 vccd1 _02486_ sky130_fd_sc_hd__a22o_1
X_14132_ _03005_ _00166_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__nand2_1
X_11344_ _01416_ _01436_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18940_ clknet_4_2_0_clk _00094_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[26\] sky130_fd_sc_hd__dfxtp_2
X_14063_ _02976_ _04241_ _03038_ _04243_ vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__or4_1
X_11275_ _01337_ _01366_ _01367_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__or3_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13014_ _01962_ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__clkbuf_8
X_10226_ _06029_ _05649_ _07112_ vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__and3_1
X_18871_ clknet_4_14_0_clk net254 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__dfxtp_1
X_10157_ _00222_ _00224_ vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__and2b_1
X_17822_ _08329_ _08330_ _08331_ vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17753_ _08171_ _08181_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__nand2_1
X_14965_ _05226_ _05227_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__and2b_1
X_10088_ _00180_ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__buf_6
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16704_ net147 _07024_ _03790_ vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__o21ai_4
X_13916_ _03138_ _03190_ _00494_ vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__mux2_1
X_17684_ _08063_ _08149_ _08182_ vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__o21ba_1
X_14896_ _05151_ _05152_ vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__nor2_1
X_16635_ _06762_ _07038_ _07039_ _06527_ vssd1 vssd1 vccd1 vccd1 _07040_ sky130_fd_sc_hd__a22o_1
X_13847_ _03830_ _03814_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16566_ _06941_ _06964_ vssd1 vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _03772_ _03773_ _03783_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nor3_2
XFILLER_0_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15517_ _05809_ _05810_ _05827_ vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__nor3_1
X_18305_ _08856_ _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12729_ _02813_ _02821_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16497_ _06811_ _06889_ _00193_ vssd1 vssd1 vccd1 vccd1 _06890_ sky130_fd_sc_hd__and3b_1
X_18236_ _08781_ _08782_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15448_ _05752_ _05753_ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _08705_ _08706_ _08707_ vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__and3_1
X_15379_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17118_ _00558_ _07355_ _02347_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap123 _02389_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_1
X_18098_ _08617_ _08618_ _08631_ vssd1 vssd1 vccd1 vccd1 _08633_ sky130_fd_sc_hd__a21oi_1
Xmax_cap134 _03587_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__buf_1
XFILLER_0_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09940_ _08832_ _08843_ _05682_ _07156_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__and4b_1
X_17049_ _07113_ net145 _07489_ _06542_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _08060_ _08082_ _08028_ _07286_ vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__o211a_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11060_ _01151_ _00176_ _00145_ _04078_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__a22o_1
X_10011_ _07657_ vssd1 vssd1 vccd1 vccd1 _09354_ sky130_fd_sc_hd__buf_4
X_14750_ _04989_ _04990_ _04991_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a21o_1
X_11962_ _01938_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__o21ai_1
X_13701_ _03845_ _03846_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__or2_1
X_10913_ _05235_ _01005_ _00983_ _00982_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__a31o_1
X_14681_ _04904_ _04905_ _04916_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__nor3_1
X_11893_ _01895_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16420_ _06803_ _06520_ net150 _06805_ sel_op\[0\] vssd1 vssd1 vccd1 vccd1 _06806_
+ sky130_fd_sc_hd__a2111o_1
X_13632_ _03768_ _03769_ _03770_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__and3_1
X_10844_ _00934_ _00935_ _00936_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _03049_ _06618_ _06730_ _06626_ vssd1 vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__o211a_1
X_13563_ _03276_ _03504_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ _00163_ _00214_ vssd1 vssd1 vccd1 vccd1 _00868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15302_ _05478_ _05553_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__a211oi_4
X_12514_ _00514_ _02214_ vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__nor2_2
X_16282_ _06655_ vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__buf_2
X_13494_ _03606_ _03608_ _03619_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__or3_4
XFILLER_0_42_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18021_ _08456_ _08457_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__nor2_1
X_15233_ _05407_ _05416_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__a21oi_1
X_12445_ _02534_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__or2b_1
XFILLER_0_112_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ _07515_ _00461_ _05856_ _03008_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__a22oi_1
X_12376_ _02330_ _02467_ _02468_ _02328_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14115_ _04297_ _04298_ _04107_ _04266_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a211oi_2
X_11327_ _01315_ _01419_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15095_ _00192_ _08876_ _05368_ vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14046_ _04222_ _04223_ _04224_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__or3_4
X_18923_ clknet_4_13_0_clk _00077_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_11258_ _01339_ _01340_ _01350_ vssd1 vssd1 vccd1 vccd1 _01351_ sky130_fd_sc_hd__o21a_1
X_10209_ _00288_ _00289_ _00290_ vssd1 vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__a21oi_1
X_18854_ clknet_4_6_0_clk net290 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__dfxtp_1
X_11189_ _00789_ _00790_ vssd1 vssd1 vccd1 vccd1 _01282_ sky130_fd_sc_hd__xor2_2
X_17805_ _08183_ _08255_ _08313_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__or3_1
X_18785_ _09297_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__dlymetal6s2s_1
X_15997_ _05736_ _00194_ vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__or2_2
X_14948_ _05116_ _05117_ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__or2_1
X_17736_ _01678_ _06442_ _08239_ vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14879_ _05132_ _05133_ vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__and2_1
X_17667_ _08162_ _08163_ vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__xnor2_1
X_16618_ _07020_ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17598_ _07207_ _07665_ _07650_ _06947_ vssd1 vssd1 vccd1 vccd1 _08089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16549_ _06942_ _06943_ _06084_ vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_128_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _08763_ _06398_ _06399_ _07084_ _08764_ vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__a311o_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09923_ _08529_ _08648_ _08637_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__o21a_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _05812_ _06960_ _07897_ _07908_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__o211a_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _07080_ _07156_ _07134_ _07058_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__a22o_1
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 _04125_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ _00643_ _00651_ _00652_ vssd1 vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__nand3_2
XFILLER_0_64_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ _00580_ _00581_ _00582_ _00537_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_106_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ _02135_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12161_ _02240_ _02253_ vssd1 vssd1 vccd1 vccd1 _02254_ sky130_fd_sc_hd__or2_4
XFILLER_0_31_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11112_ _01126_ _01131_ _01130_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a21o_1
X_12092_ _02114_ _02184_ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__nor2_1
X_11043_ _06689_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__inv_4
X_15920_ net192 _06235_ _06263_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__a21oi_2
X_15851_ _06131_ _06180_ vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_14802_ _05036_ _05037_ _05049_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__a21o_1
X_15782_ _06113_ _06115_ vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__xnor2_1
X_18570_ salida\[7\] _09114_ _09118_ salida\[39\] _09128_ vssd1 vssd1 vccd1 vccd1
+ _09136_ sky130_fd_sc_hd__a221o_1
X_12994_ _03026_ _03086_ _02720_ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__a21o_1
X_17521_ _06750_ _07745_ _08003_ vssd1 vssd1 vccd1 vccd1 _08005_ sky130_fd_sc_hd__a21oi_1
X_14733_ _04838_ _04839_ _04972_ _04974_ vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11945_ _02036_ _02037_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_143_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17452_ _07929_ vssd1 vssd1 vccd1 vccd1 _09392_ sky130_fd_sc_hd__inv_2
XFILLER_0_129_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14664_ _01317_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__clkbuf_4
X_11876_ _01933_ _01934_ _01935_ vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16403_ _03912_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__a21o_1
X_13615_ _03606_ _03608_ _03619_ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__nor3_1
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10827_ cla_inst.in2\[16\] ApproximateM_inst.lob_16.lob2.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _00920_ sky130_fd_sc_hd__and4_1
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17383_ _07747_ _07748_ _07760_ _07758_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__a31o_1
X_14595_ _03079_ _02980_ _03533_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ _03161_ _02607_ _03170_ vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or3_1
X_13546_ _00183_ _04657_ _04864_ _00184_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a22oi_1
X_10758_ _00831_ _00844_ _00850_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16265_ _03152_ _02272_ _03104_ _06467_ _06638_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__o311a_1
X_13477_ _03600_ _03601_ vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__xor2_1
X_10689_ _04001_ _04045_ _00765_ _00781_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15216_ _05459_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__xor2_1
X_18004_ _08484_ _08494_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__or2b_1
XFILLER_0_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _02515_ _02519_ _02520_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__nor3_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ _06562_ vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__buf_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15147_ _05398_ _05401_ vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__and2b_1
X_12359_ _02443_ _02445_ _02375_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15078_ _05231_ _05234_ _05232_ vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14029_ _03993_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__xor2_1
X_18906_ clknet_4_10_0_clk _00060_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[24\] sky130_fd_sc_hd__dfxtp_2
X_18837_ _09336_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__clkbuf_1
X_09570_ _03487_ _03542_ _03443_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21bo_1
X_18768_ _04725_ net39 _09276_ vssd1 vssd1 vccd1 vccd1 _09284_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17719_ _08016_ _08018_ _08121_ vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__nor3_1
X_18699_ net50 _03052_ _09182_ vssd1 vssd1 vccd1 vccd1 _09230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09906_ _08365_ _08376_ _08387_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _07722_ vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__buf_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _06971_ vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__buf_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _06202_ _06213_ _06224_ vssd1 vssd1 vccd1 vccd1 _06234_ sky130_fd_sc_hd__nand3_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer60 _05377_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__clkbuf_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer71 cla_inst.in1\[18\] vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_2
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer82 _03772_ vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _04493_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel _00179_
+ _00129_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__and4_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer93 _00333_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _01742_ _01753_ vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _03371_ _03372_ _03516_ _03517_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__o211a_2
X_10612_ _00703_ _00704_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14380_ _02188_ cla_inst.in1\[30\] _09303_ _04515_ vssd1 vssd1 vccd1 vccd1 _04589_
+ sky130_fd_sc_hd__a22o_1
X_11592_ _01647_ _01649_ vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _03440_ _00206_ _07526_ _03441_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__and4b_1
XFILLER_0_51_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10543_ _00474_ _00475_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__and2_1
X_16050_ _06402_ _06403_ _05721_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _03307_ _03309_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10474_ _00170_ _04067_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15001_ _05265_ _05266_ vssd1 vssd1 vccd1 vccd1 _05267_ sky130_fd_sc_hd__nor2_1
X_12213_ _02302_ _02304_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__or3_1
X_13193_ net131 _03266_ _03291_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12144_ _02110_ _02109_ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12075_ _01899_ _01904_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__nor2_1
X_16952_ _07285_ _07295_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__nand2_1
X_11026_ _01072_ _01074_ _01117_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__and3_1
X_15903_ _03011_ _03154_ vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__and2_1
X_16883_ _07307_ _07309_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__xor2_1
X_18622_ salida\[28\] _09159_ _09160_ salida\[60\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15834_ _06171_ _06172_ vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18553_ _09124_ vssd1 vssd1 vccd1 vccd1 _09125_ sky130_fd_sc_hd__buf_4
X_15765_ _05966_ _06045_ vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2b_1
X_12977_ _00121_ _03069_ _03024_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17504_ _07985_ _07986_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11928_ _02017_ _02020_ vssd1 vssd1 vccd1 vccd1 _02021_ sky130_fd_sc_hd__and2_1
X_14716_ _03569_ _03582_ _02978_ vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__mux2_1
X_15696_ _06004_ vssd1 vssd1 vccd1 vccd1 _06023_ sky130_fd_sc_hd__inv_2
X_18484_ _09047_ _06559_ _09050_ vssd1 vssd1 vccd1 vccd1 _09051_ sky130_fd_sc_hd__or3b_4
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _04867_ _04868_ _04879_ vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__and3_1
X_17435_ _07802_ _07803_ _07801_ vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__a21bo_1
X_11859_ _01950_ _01951_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03399_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__and4b_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14578_ _04803_ _04804_ _04628_ _04698_ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__a211oi_1
XANTENNA_29 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _07834_ _07835_ vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13529_ _03656_ _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__or2_2
X_16317_ _03047_ _07766_ _03150_ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17297_ _07749_ _07760_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16248_ _06618_ _06619_ _03152_ vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput103 net103 vssd1 vssd1 vccd1 vccd1 o_wb_data[28] sky130_fd_sc_hd__clkbuf_4
Xoutput114 net114 vssd1 vssd1 vccd1 vccd1 o_wb_data[9] sky130_fd_sc_hd__clkbuf_4
X_16179_ _06544_ vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09622_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05399_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09553_ _04635_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__buf_6
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09484_ _03771_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__buf_6
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10190_ _03848_ _03782_ _04569_ _04384_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__and4_1
X_12900_ _00189_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__clkbuf_4
X_13880_ _04024_ _04041_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__nor3_1
X_12831_ _00891_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__inv_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _05861_ _05862_ _05757_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__o21ai_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _01790_ _01798_ _01799_ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__nor3_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ net179 _04579_ _04573_ vssd1 vssd1 vccd1 vccd1 _04721_ sky130_fd_sc_hd__a21bo_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _01784_ _01787_ _01804_ _01805_ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__o211ai_2
X_15481_ _05614_ _05710_ vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__nor2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _02755_ _02785_ vssd1 vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__nand2_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _01139_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__clkbuf_4
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17220_ _02633_ _07676_ _03201_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ _01735_ _01736_ vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17151_ _07590_ _07600_ vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__xnor2_1
X_14363_ _02986_ _07134_ _04568_ _04570_ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__nand4_2
XFILLER_0_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput16 i_wb_addr[22] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
X_11575_ _01658_ _01666_ _01667_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__a21boi_1
Xinput27 i_wb_addr[3] vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__clkbuf_4
X_16102_ _02966_ _06459_ vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__nor2_1
Xinput38 i_wb_data[12] vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_2
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13314_ _03416_ _03422_ _03423_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__nand3_2
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ _00445_ _00446_ _00438_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__a21bo_1
Xinput49 i_wb_data[22] vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_2
X_17082_ _07523_ _07524_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__nand2_1
X_14294_ _00173_ _00175_ _05388_ _05050_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__and4_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16033_ _06383_ _06385_ _03588_ vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13245_ _00747_ _03203_ _03347_ _03348_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10457_ _00548_ _00549_ vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13176_ _03272_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__or2_1
X_10388_ _00476_ _00480_ vssd1 vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__xnor2_1
X_12127_ _02219_ _02209_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__xnor2_1
X_17984_ _02167_ _08424_ _02174_ vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__o21ai_1
X_12058_ _02148_ _02134_ _02149_ _02150_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__or4b_4
X_16935_ _03101_ _06436_ _07366_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11009_ _01098_ _01100_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__or2b_1
X_16866_ _06562_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nor2_1
X_18605_ _09125_ vssd1 vssd1 vccd1 vccd1 _09162_ sky130_fd_sc_hd__buf_2
X_15817_ _03012_ _03072_ _03149_ _03010_ vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16797_ _03324_ _06529_ _06814_ _02099_ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18536_ net9 net12 net11 net15 vssd1 vssd1 vccd1 vccd1 _09106_ sky130_fd_sc_hd__or4_1
X_15748_ net197 _06079_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18467_ _03036_ _06295_ _09029_ _09032_ vssd1 vssd1 vccd1 vccd1 _09033_ sky130_fd_sc_hd__o211ai_1
X_15679_ _06002_ _06003_ _05957_ _05931_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17418_ _07891_ _07892_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18398_ _04406_ _07592_ _08957_ vssd1 vssd1 vccd1 vccd1 _08958_ sky130_fd_sc_hd__nand3_1
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17349_ _06421_ _07806_ _07807_ _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09605_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05213_ sky130_fd_sc_hd__buf_4
X_09536_ _04449_ vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09467_ _03553_ _03563_ _03695_ vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nand3_1
XFILLER_0_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _01362_ _01437_ vssd1 vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _00170_ _00165_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__nand2_1
X_11291_ _01299_ _01302_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13030_ _02971_ _03122_ vssd1 vssd1 vccd1 vccd1 _09355_ sky130_fd_sc_hd__nand2_1
X_10242_ _00330_ _00331_ _00334_ _00305_ vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__o2bb2a_1
X_10173_ _00245_ _00246_ _00265_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14981_ _05156_ _05155_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__and2b_1
X_16720_ _07129_ _07131_ vssd1 vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__xnor2_2
X_13932_ _04097_ _04098_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__xor2_2
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13863_ _03862_ _03872_ vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__or2_1
X_16651_ _07055_ _07056_ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__xnor2_1
X_12814_ _02899_ _02905_ _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__and3_2
X_15602_ _05918_ _05919_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__nor2_1
X_13794_ _03945_ _03947_ _03948_ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__nor3b_4
X_16582_ _06934_ _06935_ _06980_ vssd1 vssd1 vccd1 vccd1 _06983_ sky130_fd_sc_hd__or3b_4
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18321_ _02871_ _02881_ vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__nand2_1
X_15533_ _05737_ _05755_ _05844_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__or3_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _02749_ _02748_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__or2b_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15464_ _05688_ _05770_ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__or2_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _08725_ _08726_ _08728_ _08799_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14415_ _04470_ _04488_ _04626_ _04627_ vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17203_ _06750_ _07650_ _07656_ vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__a21oi_1
X_11627_ _01716_ _01717_ _01718_ _01710_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__a22o_1
X_15395_ _05549_ _05598_ _05696_ vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a21oi_1
X_18183_ _08715_ _08723_ vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14346_ _04399_ _04400_ vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17134_ _03198_ _04956_ _07572_ _07583_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__a211o_1
X_11558_ _07352_ _05050_ _01647_ _01648_ vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _00467_ _00486_ _00487_ _00488_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17065_ _07421_ _07422_ vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__nor2_1
X_14277_ _04475_ _00715_ _07526_ _04476_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__and4b_1
XFILLER_0_111_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11489_ _01529_ _01530_ _01532_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16016_ _06331_ _06365_ _06366_ vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13228_ _03318_ _03330_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__xor2_2
XFILLER_0_21_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _03254_ _03255_ _03247_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__a21o_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17967_ _08487_ _08488_ _08489_ vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16918_ _07248_ _07252_ _07249_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__o21ai_2
X_17898_ _08252_ _08324_ vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16849_ _00167_ _07179_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18519_ _03913_ _07086_ _08141_ _09087_ vssd1 vssd1 vccd1 vccd1 _09088_ sky130_fd_sc_hd__o31a_1
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10860_ _00948_ _00952_ vssd1 vssd1 vccd1 vccd1 _00953_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _04231_ _04253_ _04263_ vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__a21bo_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10791_ _00876_ _00880_ _00883_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _02482_ _02532_ vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__or2_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12461_ _02551_ _02553_ vssd1 vssd1 vccd1 vccd1 _02554_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14200_ _04390_ _04391_ _04392_ vssd1 vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__nor3_2
XFILLER_0_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11412_ _01504_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__buf_4
X_15180_ _05362_ _05360_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and2b_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ _02422_ _02430_ vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14131_ _04127_ _04141_ _04139_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__a21o_1
X_11343_ _01434_ _01435_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14062_ _03533_ _03549_ _03099_ vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__mux2_2
X_11274_ _01335_ _01336_ _01079_ _01147_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__o211a_1
X_13013_ _03103_ _03105_ _03090_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__mux2_1
X_10225_ _06732_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__buf_4
X_18870_ clknet_4_13_0_clk net245 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__dfxtp_1
X_17821_ _08329_ _08330_ _08331_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__or3_1
X_10156_ _00164_ _00248_ vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__nand2_1
X_17752_ _08167_ _08170_ vssd1 vssd1 vccd1 vccd1 _08257_ sky130_fd_sc_hd__nand2_1
X_14964_ _05223_ _05225_ _05119_ vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__a21o_1
X_10087_ _00179_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__buf_4
X_16703_ _07113_ _06655_ _06946_ _07026_ vssd1 vssd1 vccd1 vccd1 _07114_ sky130_fd_sc_hd__and4_1
X_13915_ _04081_ _03185_ _03060_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__mux2_1
X_17683_ _08171_ _08181_ vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__xnor2_1
X_14895_ _05149_ _05150_ _05144_ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a21oi_1
X_16634_ _07033_ _07034_ _00207_ vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__o21a_4
X_13846_ _03857_ _03858_ _03874_ vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13777_ _03201_ vssd1 vssd1 vccd1 vccd1 _03930_ sky130_fd_sc_hd__clkbuf_8
X_16565_ _06950_ _06963_ vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__xor2_1
X_10989_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _01082_ sky130_fd_sc_hd__buf_4
X_18304_ _08853_ _08855_ vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__nor2_1
X_15516_ _05809_ _05810_ _05827_ vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12728_ _02810_ _02812_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16496_ _06812_ net150 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__nand2_8
XFILLER_0_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18235_ _08776_ _08780_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__and2_1
X_15447_ _05740_ _05662_ _05751_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__and3_1
X_12659_ _02742_ _02743_ _02735_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18166_ _07332_ _07665_ _08260_ _08625_ vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__or4b_2
X_15378_ _07668_ _01139_ _01223_ _03009_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ _02347_ _06510_ _02259_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14329_ _04531_ _04532_ _04492_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__o21ai_2
Xmax_cap124 _00600_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18097_ _08617_ _08618_ _08631_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap135 _03375_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_1
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17048_ _02188_ _06889_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__and2_2
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09870_ _07286_ _08028_ _08082_ _08060_ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__a211o_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18999_ clknet_4_7_0_clk _09365_ vssd1 vssd1 vccd1 vccd1 salida\[52\] sky130_fd_sc_hd__dfxtp_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10010_ _09352_ vssd1 vssd1 vccd1 vccd1 _09353_ sky130_fd_sc_hd__buf_4
X_09999_ _07482_ _07908_ _09339_ _09340_ vssd1 vssd1 vccd1 vccd1 _09342_ sky130_fd_sc_hd__a211o_2
X_11961_ _01979_ _01983_ _01982_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10912_ _04700_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__clkbuf_8
X_13700_ _00203_ _05921_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__nand2_1
X_14680_ _04904_ _04905_ _04916_ vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__o21a_1
X_11892_ _01892_ _01894_ _01893_ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ _03595_ _03602_ _03597_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10843_ _03345_ net170 _00145_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__nand4_2
XFILLER_0_67_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13562_ _03692_ _03694_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__xor2_2
X_16350_ _01677_ _06623_ vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__or2_1
X_10774_ _00860_ _00866_ vssd1 vssd1 vccd1 vccd1 _00867_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15301_ _05574_ _05592_ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__and2_1
X_12513_ _02556_ _02594_ _02603_ vssd1 vssd1 vccd1 vccd1 _02606_ sky130_fd_sc_hd__a21oi_1
X_16281_ _06427_ _06651_ vssd1 vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__nor2_2
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13493_ _03606_ _03608_ _03619_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18020_ _08546_ _08547_ vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15232_ _05404_ _05406_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__and2b_1
X_12444_ _02535_ _02536_ vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__xor2_2
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ _03006_ _01678_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12375_ _02321_ _02325_ _02327_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__a21o_1
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14114_ _04107_ _04266_ _04297_ _04298_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__o211a_2
XFILLER_0_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11326_ _00105_ _01418_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__nor2_2
X_15094_ _00192_ _08876_ _05368_ vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__a21oi_1
X_14045_ _04046_ _04048_ vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__nor2_1
X_18922_ clknet_4_9_0_clk _00076_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_11257_ _01341_ _01349_ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10208_ _00299_ _00300_ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18853_ clknet_4_6_0_clk net292 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__dfxtp_1
X_11188_ net214 _00958_ vssd1 vssd1 vccd1 vccd1 _01281_ sky130_fd_sc_hd__nor2_1
X_17804_ _08183_ _08255_ _08313_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__o21ai_2
X_10139_ _00142_ _00159_ vssd1 vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__nor2_1
X_18784_ _09273_ _09296_ vssd1 vssd1 vccd1 vccd1 _09297_ sky130_fd_sc_hd__and2_1
X_15996_ _06084_ _00878_ vssd1 vssd1 vccd1 vccd1 _06345_ sky130_fd_sc_hd__or2_2
X_17735_ _06425_ _06443_ vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__nor2_1
X_14947_ _05113_ _05114_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17666_ _07039_ net145 vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__nand2_1
X_14878_ _05124_ _05131_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ _06950_ _06963_ vssd1 vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__nor2_1
X_13829_ _09166_ cla_inst.in2\[29\] _03673_ _00211_ vssd1 vssd1 vccd1 vccd1 _03987_
+ sky130_fd_sc_hd__and4_1
X_17597_ _07302_ _07303_ _07314_ _07516_ vssd1 vssd1 vccd1 vccd1 _08088_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16548_ _06562_ _06571_ _06874_ _06944_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__or4_4
XFILLER_0_58_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16479_ sel_op\[0\] _06804_ vssd1 vssd1 vccd1 vccd1 _06870_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18218_ _08763_ _06399_ _06398_ vssd1 vssd1 vccd1 vccd1 _08764_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18149_ _06397_ _06790_ _08688_ _03052_ vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _08529_ _08637_ _08648_ vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__nor3_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _07886_ _07493_ _07482_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__nand3b_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _07102_ vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_119 _02099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10490_ _00537_ _00580_ _00581_ _00582_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__or4_4
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12160_ _02243_ _02251_ _02252_ vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11111_ _01181_ _01201_ _01077_ _01203_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12091_ _05747_ _00213_ _02112_ _02113_ vssd1 vssd1 vccd1 vccd1 _02184_ sky130_fd_sc_hd__o2bb2a_1
X_11042_ _01121_ _01133_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__nand2_1
X_15850_ _04562_ _05623_ _06152_ _03124_ _06189_ vssd1 vssd1 vccd1 vccd1 _09372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801_ _05047_ _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__xnor2_1
X_15781_ _06035_ _06044_ _06114_ vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12993_ _00223_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__clkbuf_4
X_17520_ _06750_ _07745_ _08003_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__and3_1
X_14732_ _02986_ _08224_ _04970_ _04971_ vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__a22oi_2
X_11944_ _01948_ _01947_ vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17451_ _07905_ _07909_ _07928_ _06463_ _03108_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__a32o_2
X_14663_ _04896_ _04898_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11875_ _01961_ _01965_ _01966_ _01967_ vssd1 vssd1 vccd1 vccd1 _01968_ sky130_fd_sc_hd__or4_4
XFILLER_0_129_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16402_ _06337_ _06335_ _06336_ _06598_ _06786_ vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__a311o_1
X_13614_ _03622_ _03623_ _03646_ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nand3_2
X_10826_ _00912_ _00913_ _00917_ vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__a21oi_1
X_17382_ _07851_ _07852_ vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14594_ _04818_ _04820_ _04823_ vssd1 vssd1 vccd1 vccd1 _04824_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16333_ _01503_ _03083_ _03166_ _03086_ _06477_ _03161_ vssd1 vssd1 vccd1 vccd1 _06713_
+ sky130_fd_sc_hd__mux4_1
X_13545_ _03464_ _03437_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__and2b_1
X_10757_ _00848_ _00123_ _00849_ vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_54_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _03990_ _05964_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__nand2_1
X_16264_ _03089_ _06637_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__or2_1
X_10688_ _03859_ _03793_ _04056_ _03673_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003_ _08499_ _08500_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15215_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__and2_1
X_12427_ _02448_ _02514_ _02513_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16195_ _07657_ _06541_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15146_ _03035_ _03116_ _03537_ vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__mux2_1
X_12358_ _02450_ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__inv_2
X_11309_ _01320_ _01322_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__or2b_1
X_15077_ _05250_ _05251_ vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or2_1
X_12289_ _02228_ _02351_ _02350_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14028_ _04196_ _04204_ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__xnor2_1
X_18905_ clknet_4_10_0_clk _00059_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18836_ net60 op_code\[3\] _09331_ vssd1 vssd1 vccd1 vccd1 _09336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18767_ _09283_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__buf_1
X_15979_ _00908_ _02963_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17718_ _08120_ _08219_ vssd1 vssd1 vccd1 vccd1 _08220_ sky130_fd_sc_hd__nor2_1
X_18698_ net49 _09190_ _09229_ vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17649_ _03120_ _05425_ _08140_ _08144_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09905_ _08442_ _08463_ vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09836_ cla_inst.in1\[28\] vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__clkbuf_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _06971_ sky130_fd_sc_hd__buf_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _03509_ _03804_ _03399_ _03531_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a22o_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer50 net212 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer61 _05377_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__clkbuf_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer72 net234 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer83 _03595_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer94 _01926_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _01751_ _01752_ vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__nor2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _00173_ _00175_ _04056_ _00563_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__and4_2
XFILLER_0_138_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11591_ _01208_ _01682_ _01683_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__nand3_2
XFILLER_0_106_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _09172_ _00218_ _00178_ _09166_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__a22o_1
X_10542_ _00632_ _00633_ _00450_ _00603_ vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__a211o_4
XFILLER_0_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13261_ _03352_ _03351_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or2b_1
X_10473_ _00564_ _00565_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15000_ _00189_ _00191_ _07134_ _00309_ vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__and4_1
X_12212_ _02151_ _02301_ _02290_ net322 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__a211oi_1
X_13192_ net131 _03266_ _03291_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__or3_4
XFILLER_0_103_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _06971_ _03837_ vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12074_ _02164_ _02166_ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__and2_1
X_16951_ _07331_ _07338_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__nand2_1
X_11025_ _01072_ _01074_ _01117_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__a21oi_1
X_15902_ _05652_ vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__buf_2
X_16882_ _07208_ _07211_ _07206_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__a21bo_1
X_18621_ net267 _09157_ _09171_ _09162_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__o211a_1
X_15833_ _06112_ _06162_ _06169_ vssd1 vssd1 vccd1 vccd1 _06172_ sky130_fd_sc_hd__nor3_1
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18552_ net69 vssd1 vssd1 vccd1 vccd1 _09124_ sky130_fd_sc_hd__inv_2
X_15764_ _06095_ _06096_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12976_ _03025_ _03068_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17503_ _07868_ _07870_ _07867_ vssd1 vssd1 vccd1 vccd1 _07986_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14715_ _02975_ _04955_ vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__nor2_1
X_11927_ _01952_ _02019_ vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__nor2_1
X_18483_ _08978_ _09013_ _09049_ _09012_ _09046_ vssd1 vssd1 vccd1 vccd1 _09050_ sky130_fd_sc_hd__a221o_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15695_ _06017_ _06018_ _06022_ vssd1 vssd1 vccd1 vccd1 _09369_ sky130_fd_sc_hd__o21ai_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17434_ _03107_ _07355_ _06374_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__or3b_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14646_ _04867_ _04868_ _04879_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__a21oi_1
X_11858_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel _06008_ vssd1 vssd1 vccd1
+ vccd1 _01951_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_19 _01115_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _00262_ _00901_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__and2_1
X_17365_ _06764_ _07487_ _07593_ _06653_ vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__o22a_1
X_14577_ _04628_ _04698_ _04803_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__o211a_1
X_11789_ _01828_ _01840_ _01836_ _01839_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16316_ _03199_ _03133_ _06693_ vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__a21o_1
X_13528_ _07537_ _00213_ _03655_ _03657_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17296_ _07758_ _07759_ vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16247_ _03026_ _03052_ _01114_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ _03579_ _03581_ _03098_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput104 net104 vssd1 vssd1 vccd1 vccd1 o_wb_data[29] sky130_fd_sc_hd__clkbuf_4
X_16178_ _06422_ _06459_ vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15129_ _05404_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _05377_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18819_ _09125_ _09323_ vssd1 vssd1 vccd1 vccd1 _09324_ sky130_fd_sc_hd__and2_1
X_09552_ _04493_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__buf_8
XFILLER_0_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09483_ cla_inst.in2\[16\] vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ _07526_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12830_ _02899_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__inv_2
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _01791_ _01797_ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__nand2_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _04712_ _04713_ _04718_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__a21o_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _01802_ _01803_ _01776_ _01788_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__a211o_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15480_ _05786_ _05788_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__xor2_2
X_12692_ _02783_ _02784_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__or2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _04643_ _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _01687_ _01688_ _01689_ _01701_ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17150_ _07598_ _07599_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__xnor2_2
X_14362_ _03651_ _03662_ _07102_ _05704_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__nand4_2
X_11574_ _01663_ _01665_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 i_wb_addr[23] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__clkbuf_1
Xinput28 i_wb_addr[4] vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16101_ op_code\[2\] op_code\[3\] vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__or2_2
Xinput39 i_wb_data[13] vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__buf_2
X_13313_ _03419_ _03420_ _03251_ _03252_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__o211ai_2
X_10525_ _00610_ _00611_ _00616_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__a21o_1
X_14293_ _00702_ _00443_ _06471_ _00195_ vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__a22oi_1
X_17081_ _07523_ _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__or2_1
X_13244_ _03343_ _03344_ _03346_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__o21ai_2
X_16032_ _02987_ _01678_ vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__or2_1
X_10456_ _00106_ _00206_ vssd1 vssd1 vccd1 vccd1 _00549_ sky130_fd_sc_hd__nand2_1
X_13175_ _00362_ _00878_ _03271_ _03273_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__a22oi_1
X_10387_ _00477_ _00479_ vssd1 vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12126_ _02181_ _02204_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__nor2_1
X_17983_ _08447_ _08419_ _08505_ _08508_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__o31a_1
X_12057_ _02065_ _02147_ _02143_ _02146_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__a211o_1
X_16934_ _03101_ _06436_ _06424_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__a21oi_1
X_11008_ _01098_ _01100_ vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__xnor2_1
X_16865_ _03324_ _03003_ _06814_ _07289_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__a211o_2
X_18604_ salida\[20\] _09159_ _09160_ salida\[52\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09161_ sky130_fd_sc_hd__a221o_1
X_15816_ _03007_ _03067_ vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__nand2_1
X_16796_ _07212_ _07214_ vssd1 vssd1 vccd1 vccd1 _07215_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18535_ net5 net8 net7 net10 vssd1 vssd1 vccd1 vccd1 _09105_ sky130_fd_sc_hd__or4_1
X_15747_ _05795_ _06075_ _06077_ _06078_ vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__o211a_1
X_12959_ _01112_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18466_ _03913_ _06913_ _08141_ _09031_ _06721_ vssd1 vssd1 vccd1 vccd1 _09032_ sky130_fd_sc_hd__o311a_1
XFILLER_0_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15678_ _05957_ _05931_ _06002_ _06003_ vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__o211a_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17417_ _07883_ _07890_ vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__or2_1
X_14629_ _04852_ _04854_ _04859_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18397_ _08955_ _08956_ vssd1 vssd1 vccd1 vccd1 _08957_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _03198_ _05096_ _06543_ _07809_ _07816_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17279_ _02124_ _07592_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__nand2_4
XFILLER_0_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19018_ clknet_4_9_0_clk _00003_ vssd1 vssd1 vccd1 vccd1 sel_op\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09604_ _04733_ _04624_ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__or2b_1
X_09535_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel vssd1 vssd1 vccd1 vccd1
+ _04449_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ _03585_ _03640_ _03684_ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10310_ _00203_ _00248_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_132_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11290_ _01297_ _01298_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10241_ _00303_ _00304_ _08529_ _08659_ vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__a211oi_1
X_10172_ _00249_ _00264_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14980_ _05009_ _05154_ vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and2b_1
X_13931_ _03933_ _03934_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__nand2_1
X_16650_ _06749_ _06969_ vssd1 vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__nand2_1
X_13862_ _04021_ _04022_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__xor2_2
XFILLER_0_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15601_ _05918_ _05919_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__and2_1
X_12813_ _00854_ _02898_ _01465_ _01466_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o211ai_1
X_16581_ _06934_ _06935_ _06980_ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__o21ba_1
X_13793_ _03762_ _03767_ _03761_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18320_ _08872_ _08840_ _08841_ vssd1 vssd1 vccd1 vccd1 _08874_ sky130_fd_sc_hd__and3_1
X_15532_ _05737_ _05755_ _05844_ vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__o21ai_2
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12744_ _02634_ _02668_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__xnor2_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _08730_ _08729_ vssd1 vssd1 vccd1 vccd1 _08799_ sky130_fd_sc_hd__or2b_1
X_15463_ _05688_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__nand2_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12675_ _02766_ _02767_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ _06750_ _07650_ _07656_ vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__and3_1
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14414_ _04608_ _04609_ _04625_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__a21oi_1
X_11626_ _01710_ _01716_ _01717_ _01718_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__nand4_2
X_18182_ _08715_ _08723_ vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__and2_1
X_15394_ _05694_ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17133_ _06462_ _07574_ _07576_ _07582_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__or4_1
X_14345_ _04550_ _04551_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11557_ _05682_ _03750_ _01597_ _01596_ _04143_ vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _00291_ _00431_ _00465_ _00466_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__o211a_1
X_17064_ _07484_ _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__xor2_1
X_14276_ _07504_ _04012_ _04045_ _00358_ vssd1 vssd1 vccd1 vccd1 _04476_ sky130_fd_sc_hd__a22o_1
X_11488_ _01573_ _01574_ _01580_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nand3_2
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16015_ _02347_ _00558_ vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__and2_1
X_10439_ _00529_ _00530_ _00349_ _00531_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__o211ai_4
X_13227_ _03319_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _03247_ _03254_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__nand3_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _02140_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__and2_1
X_13089_ _02505_ _02259_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__nor2_1
X_17966_ _08487_ _08488_ _08489_ vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__and3_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16917_ _07345_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__nor2_1
X_17897_ _08016_ _08121_ _08414_ vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__or3_1
XFILLER_0_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16848_ _06424_ _06436_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779_ _06563_ _07195_ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nor2_1
X_18518_ _06680_ _09086_ vssd1 vssd1 vccd1 vccd1 _09087_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18449_ _09011_ _09012_ vssd1 vssd1 vccd1 vccd1 _09013_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_384 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09518_ net227 net169 _03421_ _04242_ vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__nand4_2
X_10790_ _00882_ _00208_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__xnor2_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _03498_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__buf_6
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12460_ _06971_ _00177_ _02551_ _02552_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__nand4_2
XFILLER_0_47_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11411_ _00170_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12391_ _02482_ _02483_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14130_ _04313_ _04314_ _04123_ _04145_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__a211oi_4
X_11342_ _01421_ _01433_ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11273_ _01267_ _01365_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__xnor2_1
X_14061_ _03913_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10224_ _06051_ _07156_ _07134_ _06040_ vssd1 vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__a22o_1
X_13012_ _02373_ _03104_ _03040_ vssd1 vssd1 vccd1 vccd1 _03105_ sky130_fd_sc_hd__o21ai_2
X_17820_ _08231_ _08233_ _08230_ vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__a21boi_2
X_10155_ _00247_ vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__clkbuf_4
X_17751_ _08185_ _08201_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__nor2_1
X_14963_ _05119_ _05223_ _05225_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10086_ ApproximateM_inst.lob_16.lob1.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00179_ sky130_fd_sc_hd__buf_4
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16702_ _06567_ _06570_ _00357_ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__o21a_1
X_13914_ _03177_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__inv_2
X_17682_ _08172_ _08179_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__xnor2_1
X_14894_ _05144_ _05149_ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__and3_1
X_16633_ _06807_ vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__clkbuf_4
X_13845_ _04002_ _04003_ _03811_ _03833_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__o211a_1
X_16564_ _06959_ _06962_ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__xnor2_1
X_13776_ _03904_ _03905_ _03929_ vssd1 vssd1 vccd1 vccd1 _09380_ sky130_fd_sc_hd__o21ai_2
X_10988_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _01081_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18303_ _08853_ _08855_ vssd1 vssd1 vccd1 vccd1 _08856_ sky130_fd_sc_hd__and2_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15515_ _05825_ _05826_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__nor2_1
X_12727_ _02803_ _02819_ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__nor2_1
X_16495_ _06867_ _06887_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18234_ _08776_ _08780_ vssd1 vssd1 vccd1 vccd1 _08781_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15446_ _05740_ _05662_ _05751_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12658_ _02746_ _02750_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11609_ _01585_ _01602_ _01700_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__a211oi_2
X_18165_ _07665_ _07708_ _08150_ _07216_ vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__a22o_1
X_15377_ _03006_ _04336_ vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12589_ _02597_ _02640_ _02639_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17116_ _07562_ _03930_ _07563_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__and3_1
X_14328_ _04492_ _04531_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__or3_4
XFILLER_0_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18096_ _08629_ _08630_ vssd1 vssd1 vccd1 vccd1 _08631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap125 _01707_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__clkbuf_2
Xmax_cap147 _07023_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_1
X_17047_ _06563_ _06572_ _07387_ _07487_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__or4_2
X_14259_ _04445_ _04446_ _04456_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ clknet_4_7_0_clk _09364_ vssd1 vssd1 vccd1 vccd1 salida\[51\] sky130_fd_sc_hd__dfxtp_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _08353_ _08355_ vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09998_ _09339_ _09340_ _07482_ _07908_ vssd1 vssd1 vccd1 vccd1 _09341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11960_ _02027_ _02052_ _01967_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__o21ai_2
X_10911_ _01000_ _01003_ vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11891_ _01979_ _01982_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__or3_4
X_13630_ _03761_ _03762_ _03767_ vssd1 vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__a21o_1
X_10842_ net169 _00179_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ net227 vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__a22o_1
X_13561_ _00164_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10773_ _00118_ _00865_ vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15300_ _05574_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _02556_ _02594_ _02603_ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__and3_1
X_16280_ _06561_ _06572_ _06579_ _06653_ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__or4_1
X_13492_ _03609_ _03617_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15231_ _05516_ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__or2b_1
X_12443_ _00357_ _02487_ _02486_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15162_ _05432_ _05441_ vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12374_ _02398_ _02465_ _02466_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _04283_ net133 _04295_ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__or3_1
X_11325_ _01356_ _07646_ _09354_ _01417_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__a22oi_1
X_15093_ _00189_ _07134_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__and2_1
X_14044_ net319 _04219_ _04221_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__o21a_1
X_11256_ _01347_ _01348_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__nor2_1
X_18921_ clknet_4_13_0_clk _00075_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[7\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _08615_ _05856_ _08572_ _08561_ vssd1 vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a31o_1
X_11187_ _00969_ _00971_ _00970_ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__o21ba_1
X_18852_ clknet_4_6_0_clk net286 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__dfxtp_1
X_17803_ _08294_ _08312_ vssd1 vssd1 vccd1 vccd1 _08313_ sky130_fd_sc_hd__xor2_1
X_10138_ _00162_ _00230_ vssd1 vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__nand2_2
X_18783_ _02987_ net44 _09276_ vssd1 vssd1 vccd1 vccd1 _09296_ sky130_fd_sc_hd__mux2_1
X_15995_ _05747_ _00223_ vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__nand2_1
X_17734_ _03588_ _06385_ _06383_ vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__a21o_1
X_14946_ _05173_ _05174_ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__or2b_1
X_10069_ _00160_ _00141_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17665_ _08160_ _08161_ vssd1 vssd1 vccd1 vccd1 _08162_ sky130_fd_sc_hd__nand2_1
X_14877_ _05124_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or2_1
X_16616_ _06937_ _07018_ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__or2_1
X_13828_ cla_inst.in2\[31\] _00207_ vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__nand2_1
X_17596_ _07038_ _07623_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16547_ _06942_ _06943_ _06084_ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__a21bo_2
X_13759_ _03909_ _03910_ _02981_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16478_ _03003_ _03004_ _06523_ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__or3_1
XFILLER_0_143_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18217_ _02994_ _04900_ vssd1 vssd1 vccd1 vccd1 _08763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15429_ _05685_ _05732_ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18148_ _02997_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18079_ _06421_ _08597_ _08598_ _08606_ _08612_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__a311o_1
XFILLER_0_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _08496_ _08507_ _08518_ vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _07482_ _07493_ _07886_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__a21bo_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _07058_ _07091_ _07123_ _07134_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__nand4_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _01074_ _01075_ _01202_ _01053_ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__o2bb2a_1
X_12090_ _02177_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__nand2_1
X_11041_ _01121_ _01133_ vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__or2_1
X_14800_ _02999_ _04900_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__nand2_1
X_15780_ _06043_ _06036_ vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12992_ _03024_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14731_ _02986_ _07384_ _04970_ _04971_ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__and4_1
X_11943_ _00832_ _04886_ vssd1 vssd1 vccd1 vccd1 _02036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ _06836_ _07913_ _07915_ _07927_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__o31a_1
X_14662_ _04885_ _04768_ _04895_ vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__and3_1
X_11874_ _01864_ _01964_ vssd1 vssd1 vccd1 vccd1 _01967_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16401_ _06337_ _06336_ _06335_ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__a21oi_1
X_13613_ _03649_ _03650_ _03670_ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nor3_1
X_17381_ _07822_ _07729_ _07850_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__and3_1
X_10825_ _00912_ _00913_ _00917_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__and3_1
X_14593_ _03930_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16332_ _03916_ _06710_ vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__and2_1
X_13544_ _03438_ _03463_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10756_ _00831_ _00844_ vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16263_ _03026_ _03108_ _01963_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__a21o_1
X_13475_ _03598_ _03599_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10687_ _04668_ _04679_ _04711_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__o21ai_1
X_18002_ _08509_ _08511_ _08528_ _06723_ _00813_ vssd1 vssd1 vccd1 vccd1 _09399_ sky130_fd_sc_hd__o32a_1
X_15214_ _05460_ _05384_ _05498_ vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__nand3_1
XFILLER_0_124_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12426_ _02439_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__xnor2_1
X_16194_ net334 vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__buf_2
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15145_ _04823_ _05417_ _05418_ _05424_ vssd1 vssd1 vccd1 vccd1 _09361_ sky130_fd_sc_hd__a31o_1
X_12357_ _02416_ _02448_ net128 _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _01399_ _01400_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__or2_1
X_15076_ _05258_ _05256_ vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__and2b_1
X_12288_ _02378_ _02379_ _02368_ _02376_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__o211a_1
X_14027_ _04197_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__xnor2_1
X_18904_ clknet_4_10_0_clk _00058_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[22\] sky130_fd_sc_hd__dfxtp_4
X_11239_ _01313_ _01314_ _01330_ _01331_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__a211o_2
X_18835_ _09335_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__clkbuf_1
X_18766_ _09273_ _09282_ vssd1 vssd1 vccd1 vccd1 _09283_ sky130_fd_sc_hd__and2_1
X_15978_ _06323_ _06324_ _06325_ _03039_ vssd1 vssd1 vccd1 vccd1 _09378_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_117_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17717_ _08014_ _08119_ vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__nor2_1
X_14929_ _05065_ _05067_ _05187_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18697_ _01136_ _09183_ net69 vssd1 vssd1 vccd1 vccd1 _09229_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17648_ _06630_ _08141_ _08143_ _06720_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17579_ _07751_ _07394_ _07604_ _07039_ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ _03728_ _08452_ vssd1 vssd1 vccd1 vccd1 _08463_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _07700_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__clkbuf_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _05943_ _06138_ _05812_ _05823_ vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__a211oi_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _03465_ _03914_ vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__and2_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer40 _02693_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__buf_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer51 _00956_ vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer62 _03590_ vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_6
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer73 _03772_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer95 _04549_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__buf_6
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _00702_ _04154_ _00165_ _00195_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11590_ _06982_ _00443_ _01206_ _01207_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ _00450_ net143 _00632_ _00633_ vssd1 vssd1 vccd1 vccd1 _00634_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13260_ _03125_ _03133_ _03196_ _03199_ _03364_ vssd1 vssd1 vccd1 vccd1 _09366_ sky130_fd_sc_hd__a221o_1
X_10472_ _00173_ _00183_ _03673_ _00211_ vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__and4_1
X_12211_ _02131_ _02303_ vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _03267_ _03290_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12142_ _02211_ _02213_ vssd1 vssd1 vccd1 vccd1 _02235_ sky130_fd_sc_hd__nor2_1
X_12073_ _02165_ _02080_ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__xnor2_2
X_16950_ _07328_ _07329_ vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__or2b_1
X_11024_ _01104_ _01116_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__xnor2_1
X_15901_ _06242_ _06243_ vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__and2_1
X_16881_ _07305_ _07306_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__xnor2_1
X_15832_ _06112_ _06162_ _06169_ vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__o21a_1
X_18620_ salida\[27\] _09159_ _09160_ salida\[59\] _09163_ vssd1 vssd1 vccd1 vccd1
+ _09171_ sky130_fd_sc_hd__a221o_1
XFILLER_0_99_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15763_ _06088_ _06093_ vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nand2_1
X_18551_ salida\[0\] _09114_ _09118_ salida\[32\] _09121_ vssd1 vssd1 vccd1 vccd1
+ _09122_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12975_ _03067_ vssd1 vssd1 vccd1 vccd1 _03068_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14714_ _03562_ _03577_ _03079_ vssd1 vssd1 vccd1 vccd1 _04955_ sky130_fd_sc_hd__mux2_1
X_17502_ _07982_ _07983_ vssd1 vssd1 vccd1 vccd1 _07985_ sky130_fd_sc_hd__xnor2_1
X_11926_ _06711_ _04067_ _02018_ _01951_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_87_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18482_ _08969_ _09011_ vssd1 vssd1 vccd1 vccd1 _09049_ sky130_fd_sc_hd__or2_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15694_ _03547_ _04249_ _05307_ _06021_ _03039_ vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__o32a_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _06374_ _06511_ _02044_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__a21oi_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _04877_ _04878_ vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__and2_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11857_ _06008_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _01950_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10808_ _00249_ _00264_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__or2b_1
X_17364_ _06655_ _06762_ _07489_ _07596_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__and4_1
X_14576_ _04758_ _04759_ _04801_ _04802_ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11788_ _01540_ _01879_ _01880_ vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__nand3_2
XFILLER_0_103_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16315_ _06508_ _06676_ _06677_ _06692_ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13527_ _03654_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__inv_2
X_10739_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00832_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17295_ _07756_ _07757_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__and2_1
XFILLER_0_153_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16246_ _03027_ _03044_ _01224_ vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13458_ _03090_ _03189_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _01105_ _00514_ _02099_ _00212_ vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__or4b_4
XFILLER_0_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16177_ _06418_ _06422_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__nor2_4
X_13389_ _03494_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__xnor2_1
Xoutput105 net105 vssd1 vssd1 vccd1 vccd1 o_wb_data[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15128_ _05405_ _05296_ vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__or2_2
XFILLER_0_121_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15059_ _05223_ _05329_ vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__xor2_1
XFILLER_0_49_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09620_ cla_inst.in1\[18\] vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__buf_6
X_18818_ _03013_ net56 _09301_ vssd1 vssd1 vccd1 vccd1 _09323_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09551_ _04329_ _04613_ vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__xnor2_2
X_18749_ _09245_ _09268_ vssd1 vssd1 vccd1 vccd1 _09269_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09482_ _03793_ _03815_ _03837_ _03859_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09818_ cla_inst.in2\[28\] vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__buf_2
X_09749_ _06732_ vssd1 vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__inv_4
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _00591_ _01248_ _01247_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__a31o_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _01776_ _01788_ _01802_ net210 vssd1 vssd1 vccd1 vccd1 _01804_ sky130_fd_sc_hd__o211ai_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12691_ _07788_ _07570_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14430_ _04503_ _04505_ _04502_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__o21ai_4
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _01733_ _01734_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ _03377_ _07102_ _05693_ _03356_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11573_ _01663_ _01665_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput18 i_wb_addr[24] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_1
X_16100_ _06326_ _04823_ _06327_ _06458_ vssd1 vssd1 vccd1 vccd1 _09418_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13312_ _03251_ _03252_ _03419_ _03420_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a211o_2
Xinput29 i_wb_addr[5] vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__clkbuf_1
X_10524_ _00610_ _00611_ _00616_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__nand3_1
X_17080_ _07419_ _07420_ _07416_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__o21a_1
X_14292_ _04345_ _04344_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16031_ _06380_ _06381_ _06382_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__a21bo_1
X_13243_ _03343_ _03344_ _03346_ vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__or3_4
XFILLER_0_122_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ _00546_ _00547_ vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13174_ _03270_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__inv_2
X_10386_ _08158_ _00319_ _00478_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _02213_ _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__nor2_1
X_17982_ _06559_ _08506_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _02107_ _02133_ _02122_ _02132_ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__o211a_1
X_16933_ _06361_ _06359_ _06360_ _06598_ _07364_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__a311oi_1
X_11007_ _01084_ _01099_ vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__and2b_1
X_16864_ _05453_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__inv_2
X_18603_ _09117_ vssd1 vssd1 vccd1 vccd1 _09160_ sky130_fd_sc_hd__clkbuf_4
X_15815_ _03537_ _04560_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__a21o_1
X_16795_ _06766_ _06875_ _07116_ _07213_ vssd1 vssd1 vccd1 vccd1 _07214_ sky130_fd_sc_hd__o31a_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18534_ net29 net31 net30 net33 vssd1 vssd1 vccd1 vccd1 _09104_ sky130_fd_sc_hd__or4_2
X_15746_ _05945_ _06013_ _06014_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__o21ba_1
X_12958_ _03043_ _03046_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11909_ _04362_ _01031_ _09179_ _04340_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15677_ _06000_ _06001_ _05968_ vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__a21o_1
X_18465_ _06411_ _06546_ _09030_ _03073_ vssd1 vssd1 vccd1 vccd1 _09031_ sky130_fd_sc_hd__a22oi_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _01677_ vssd1 vssd1 vccd1 vccd1 _02982_ sky130_fd_sc_hd__clkbuf_4
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17416_ _07883_ _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__nand2_1
X_14628_ _04852_ _04854_ _04859_ vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__or3_4
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18396_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08956_ sky130_fd_sc_hd__or2_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ _06680_ _07812_ _07815_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__or3_1
X_14559_ _00107_ _05888_ vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _07606_ _07614_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19017_ clknet_4_9_0_clk _00002_ vssd1 vssd1 vccd1 vccd1 sel_op\[2\] sky130_fd_sc_hd__dfxtp_1
X_16229_ _06477_ _03029_ _02784_ _06333_ _06598_ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__a41o_1
XFILLER_0_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09603_ _04329_ _04613_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09534_ _04427_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__buf_8
XFILLER_0_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09465_ _03651_ _03662_ _03673_ _03618_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nand4_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _00305_ _00330_ _00331_ _00332_ vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__and4b_2
XFILLER_0_30_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _00262_ _00263_ vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13930_ _04095_ _04096_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or2_1
X_13861_ _00163_ _01678_ vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__nand2_1
X_15600_ _02998_ _04125_ _05832_ _05833_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a31o_1
X_12812_ _02903_ _02904_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__xor2_1
X_16580_ _06936_ _06979_ vssd1 vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__xnor2_1
X_13792_ _03938_ _03939_ _03944_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15531_ _05830_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12743_ _02776_ _02834_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__a21boi_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18250_ _08796_ _08797_ vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__xnor2_1
X_15462_ _05767_ _05768_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and2_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12674_ _02727_ _02730_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__xnor2_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _07654_ _07655_ vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__nor2_1
X_14413_ _04608_ _04609_ _04625_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11625_ _01708_ _01709_ _01610_ _01619_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__a211o_1
X_18181_ _08716_ _08722_ vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__xnor2_1
X_15393_ _05692_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__nand3_2
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17132_ _03920_ _07578_ _07580_ _06484_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__o211a_1
X_14344_ _04546_ _04547_ _04420_ _04397_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__o211a_1
X_11556_ _06982_ _05050_ _01647_ _01648_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__nand4_1
XFILLER_0_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10507_ _00537_ _00580_ _00581_ _00582_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__nor4_1
X_17063_ _07496_ _07505_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__xnor2_1
X_14275_ _00358_ _09172_ _04864_ _04143_ vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__and4_1
X_11487_ _01576_ _01579_ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16014_ _06363_ _06364_ _01041_ vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__a21bo_1
X_13226_ _03320_ _03328_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__xnor2_2
X_10438_ _00349_ _00350_ _00367_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__nand3_2
XFILLER_0_20_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _03252_ _03253_ _03248_ _03249_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__a211o_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _06460_ _00461_ _00296_ _00295_ vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _02200_ _09354_ _02139_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a21o_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _02257_ _03179_ _03040_ vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__o21ai_1
X_17965_ _07207_ _07623_ _08384_ _08386_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__a31o_1
X_12039_ _02123_ _02129_ _02130_ _02131_ vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__or4_4
X_16916_ _07283_ _07284_ _07344_ vssd1 vssd1 vccd1 vccd1 _07346_ sky130_fd_sc_hd__and3_1
X_17896_ _08218_ _08324_ _08325_ vssd1 vssd1 vccd1 vccd1 _08414_ sky130_fd_sc_hd__nand3_1
X_16847_ _03920_ _07268_ _07270_ _06484_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__o211a_1
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_125_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16778_ _07194_ vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18517_ _06416_ _06545_ _09085_ _06246_ vssd1 vssd1 vccd1 vccd1 _09086_ sky130_fd_sc_hd__a22o_1
X_15729_ _05989_ _05998_ _06057_ vssd1 vssd1 vccd1 vccd1 _06059_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18448_ _08915_ _08965_ _09010_ vssd1 vssd1 vccd1 vccd1 _09012_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18379_ _07474_ _08036_ _08937_ _06720_ vssd1 vssd1 vccd1 vccd1 _08938_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09517_ net169 ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel _04242_
+ net227 vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ cla_inst.in2\[17\] vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__buf_6
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11410_ _00108_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ _02435_ _02440_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11341_ _01421_ _01433_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14060_ _04237_ _04239_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11272_ _01338_ _01364_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13011_ _03028_ _02127_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__nor2_2
X_10223_ _00314_ _00315_ vssd1 vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10154_ _04067_ vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__clkbuf_8
X_17750_ _08215_ _08214_ vssd1 vssd1 vccd1 vccd1 _08254_ sky130_fd_sc_hd__or2b_1
X_14962_ _05208_ _05209_ _05222_ vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__nand3_1
X_10085_ _00177_ vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__buf_4
X_16701_ _07107_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13913_ _04077_ _04079_ _03081_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__mux2_1
X_17681_ _08173_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__xnor2_1
X_14893_ _00107_ _01223_ _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__a22o_1
X_13844_ _03811_ _03833_ _04002_ net239 vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__a211oi_2
X_16632_ _06560_ _06764_ _06951_ _07035_ vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13775_ _03123_ _03923_ _03928_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__or3_2
X_16563_ _06578_ _06961_ vssd1 vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__nor2_1
X_10987_ _07984_ _07973_ cla_inst.in1\[20\] net233 vssd1 vssd1 vccd1 vccd1 _01080_
+ sky130_fd_sc_hd__nand4_1
X_18302_ _07665_ _07516_ _08150_ _08625_ _08781_ vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__a41o_1
XFILLER_0_139_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15514_ _05728_ _05730_ _05824_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__nor3_1
X_12726_ _02804_ _02813_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_139_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16494_ _06868_ _06886_ vssd1 vssd1 vccd1 vccd1 _06887_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15445_ _05749_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__nand2_1
X_18233_ _08777_ _08779_ vssd1 vssd1 vccd1 vccd1 _08780_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12657_ _02748_ _02749_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11608_ _01699_ _01691_ _01690_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15376_ _05528_ _05531_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__and2_1
XFILLER_0_108_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18164_ _07751_ _07314_ _08260_ _08625_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__or4b_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ _02675_ _02679_ _02680_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14327_ _04529_ _04530_ _04511_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17115_ _02671_ _02842_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11539_ _01625_ _01626_ _01629_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__a21o_1
X_18095_ _08624_ _08628_ vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__nand2_1
Xmax_cap115 _08985_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_1
Xmax_cap126 _04670_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_1
XFILLER_0_111_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17046_ _07486_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__clkbuf_4
X_14258_ _04447_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__xnor2_2
Xmax_cap137 _02565_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__buf_1
XFILLER_0_150_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13209_ _03307_ _03309_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__xnor2_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14189_ _04378_ _04379_ _04161_ _04335_ vssd1 vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ clknet_4_3_0_clk _09363_ vssd1 vssd1 vccd1 vccd1 salida\[50\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _08368_ _08371_ _08369_ vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17879_ _08382_ _08287_ _08393_ vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09997_ _09338_ _09337_ _06873_ _06819_ vssd1 vssd1 vccd1 vccd1 _09340_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10910_ _01001_ _01002_ vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__and2b_1
X_11890_ _01978_ _01945_ _01976_ vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _03454_ _00129_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ _05921_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__clkbuf_4
X_10772_ _00863_ _00864_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12511_ _02556_ _02594_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__nand3_1
X_13491_ _03615_ _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__and2b_1
XFILLER_0_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15230_ _05426_ _05427_ _05515_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__or3_2
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12442_ _05747_ _00132_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15161_ _05439_ _05440_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12373_ _02320_ _02312_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__xnor2_1
X_14112_ _04283_ net133 _04295_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11324_ _09351_ vssd1 vssd1 vccd1 vccd1 _01417_ sky130_fd_sc_hd__clkbuf_4
X_15092_ _05364_ _05365_ vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14043_ _04218_ _04219_ _04221_ vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__nor3_1
X_18920_ clknet_4_13_0_clk _00074_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
X_11255_ _01344_ _01345_ _01346_ vssd1 vssd1 vccd1 vccd1 _01348_ sky130_fd_sc_hd__o21ba_1
X_10206_ _00292_ _00298_ vssd1 vssd1 vccd1 vccd1 _00299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18851_ clknet_4_6_0_clk net300 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__dfxtp_1
X_11186_ _01275_ _01276_ _01278_ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__a21oi_4
X_17802_ _08296_ _08310_ vssd1 vssd1 vccd1 vccd1 _08312_ sky130_fd_sc_hd__xnor2_1
X_10137_ _00168_ _00229_ vssd1 vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__xnor2_4
X_18782_ _09294_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__buf_1
X_15994_ _06084_ _00878_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__nand2_2
X_17733_ _03588_ _06383_ _06385_ vssd1 vssd1 vccd1 vccd1 _08237_ sky130_fd_sc_hd__nand3_1
X_14945_ _05190_ _05193_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__or2b_1
X_10068_ _00141_ _00160_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__or2b_1
X_17664_ _07042_ _07487_ _08056_ vssd1 vssd1 vccd1 vccd1 _08161_ sky130_fd_sc_hd__or3_1
X_14876_ _05128_ _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16615_ _06816_ vssd1 vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__clkbuf_4
X_13827_ _03816_ _03825_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__and2b_1
X_17595_ _07956_ _07961_ _08085_ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16546_ _05410_ _06812_ _03003_ _03004_ vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__or4_1
X_13758_ _03093_ _03096_ _03050_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__mux2_1
X_12709_ _02792_ _02793_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__nor2_1
X_13689_ _03649_ _03751_ _03832_ _03833_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16477_ _06653_ _06756_ vssd1 vssd1 vccd1 vccd1 _06868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18216_ _03201_ _08760_ _08761_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__and3_2
X_15428_ _05730_ _05731_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15359_ _01505_ _00495_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__nand2_1
X_18147_ _06425_ _06446_ _08686_ vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__or3_1
XFILLER_0_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18078_ _08609_ _08610_ _08611_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__a21oi_1
X_09920_ _08605_ _08626_ vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17029_ _03101_ _06436_ _00593_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09851_ _07690_ _07875_ vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__xnor2_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _06722_ vssd1 vssd1 vccd1 vccd1 _07134_ sky130_fd_sc_hd__buf_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11040_ _01126_ _01132_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12991_ _03026_ _03083_ _02783_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__a21bo_1
X_14730_ _02984_ _01520_ _00498_ _07015_ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nand4_1
X_11942_ _02032_ _02034_ vssd1 vssd1 vccd1 vccd1 _02035_ sky130_fd_sc_hd__nor2_2
XFILLER_0_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14661_ _04885_ _04768_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__a21oi_4
X_11873_ _00846_ _05921_ _01863_ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16400_ _02807_ _02822_ _03201_ vssd1 vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__o21ai_1
X_13612_ _03039_ _03565_ _03584_ _03121_ _03749_ vssd1 vssd1 vccd1 vccd1 _09379_ sky130_fd_sc_hd__o221ai_2
X_10824_ _00914_ _00915_ _00916_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17380_ _07822_ _07729_ _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__a21oi_1
X_14592_ _04818_ _04820_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13543_ _03671_ _03672_ _03434_ _03586_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16331_ _06707_ _06709_ _03060_ vssd1 vssd1 vccd1 vccd1 _06710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ _08191_ _00122_ _00847_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16262_ _03077_ _06632_ _06634_ vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__a21oi_1
X_13474_ _04088_ _03892_ _05617_ _05246_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__nand4_2
X_10686_ _00762_ _00763_ _00778_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__nand3_4
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _05460_ _05384_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__a21o_1
X_18001_ _07256_ _08515_ _08516_ _08527_ vssd1 vssd1 vccd1 vccd1 _08528_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ _02516_ _02483_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16193_ _06522_ _06525_ _01113_ vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ _05307_ _05419_ _05423_ _03039_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__o22ai_2
X_12356_ _02380_ _02381_ _02382_ _02352_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11307_ _00843_ _00841_ _00836_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15075_ _05132_ _05255_ vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__and2b_1
XFILLER_0_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ _02368_ _02376_ _02378_ _02379_ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14026_ _04201_ _04202_ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__xnor2_1
X_18903_ clknet_4_10_0_clk _00057_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[21\] sky130_fd_sc_hd__dfxtp_1
X_11238_ net325 _01328_ _01016_ _01014_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__o211a_1
X_18834_ net57 op_code\[2\] _09331_ vssd1 vssd1 vccd1 vccd1 _09335_ sky130_fd_sc_hd__mux2_1
X_11169_ _01243_ _01260_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__nor2_1
X_18765_ _02347_ net38 _09276_ vssd1 vssd1 vccd1 vccd1 _09282_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15977_ _05308_ _05306_ _03920_ vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ _08216_ _08217_ vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__xor2_1
X_14928_ _05065_ _05067_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__a21o_1
X_18696_ net48 _09189_ _09228_ vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _06381_ _06790_ _08142_ _03111_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__a22oi_1
X_14859_ _05110_ _05111_ vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17578_ _02347_ _06891_ _07943_ vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16529_ _06424_ _06432_ _06924_ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09903_ _04580_ vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09834_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _07700_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _05181_ _06181_ _06906_ _06928_ vssd1 vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__a211oi_1
X_09696_ _03356_ _03377_ _03903_ _03410_ vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__nand4_2
XFILLER_0_69_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer30 _01971_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__clkbuf_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer41 _01659_ vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer52 net342 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer63 net225 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer74 _02043_ vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer85 _04432_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer96 _06524_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _00620_ _00621_ _00631_ vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__or3_4
XFILLER_0_134_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10471_ _00175_ _00563_ _00211_ _00173_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_44_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ _02285_ _02287_ vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__nor2_1
X_13190_ _03268_ _03289_ vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__xnor2_2
X_12141_ _07363_ _04067_ _02232_ _02233_ vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12072_ _01990_ _02000_ vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__nand2_1
X_11023_ _01110_ _01111_ _01115_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__or3_1
X_15900_ _06211_ _06241_ vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__or2_1
X_16880_ _06874_ _06961_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__or2_1
X_15831_ _06167_ _06168_ vssd1 vssd1 vccd1 vccd1 _06169_ sky130_fd_sc_hd__and2_1
X_18550_ _09119_ _09120_ _09097_ vssd1 vssd1 vccd1 vccd1 _09121_ sky130_fd_sc_hd__o21ai_1
X_12974_ _09059_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__buf_2
X_15762_ _06088_ _06093_ vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17501_ _06875_ _07516_ vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14713_ _04946_ _04951_ _03202_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__o21a_1
X_11925_ net183 vssd1 vssd1 vccd1 vccd1 _02018_ sky130_fd_sc_hd__inv_2
X_18481_ _08969_ _08978_ _09011_ _09012_ _09046_ vssd1 vssd1 vccd1 vccd1 _09047_ sky130_fd_sc_hd__o311a_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _02974_ _04248_ _06020_ vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__o21a_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _02529_ _07906_ _07907_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__o21ai_2
X_14644_ _04869_ _04876_ vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__nand2_1
X_11856_ _07363_ _00715_ _01947_ _01948_ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__a31o_2
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _00893_ _00898_ _00430_ _00899_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14575_ _04758_ _04759_ _04801_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nand4_2
X_17363_ _07707_ _07832_ vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11787_ _01526_ _01539_ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16314_ _02810_ _03201_ _06679_ _06691_ vssd1 vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__a31o_1
X_13526_ _03654_ _00212_ _07526_ _03655_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__and4b_1
X_10738_ _08017_ _00830_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17294_ _07756_ _07757_ vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16245_ _06611_ _06616_ _03098_ vssd1 vssd1 vccd1 vccd1 _06617_ sky130_fd_sc_hd__mux2_1
X_13457_ _02982_ _03135_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__or2_1
X_10669_ _04296_ _04187_ _04285_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__nand3_2
XFILLER_0_141_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _02485_ _02499_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__xor2_1
X_13388_ _03276_ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__xor2_1
X_16176_ _07657_ net168 vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__and2_2
Xoutput106 net106 vssd1 vssd1 vccd1 vccd1 o_wb_data[30] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15127_ _05292_ _05294_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__and2b_1
X_12339_ _02422_ _02430_ _02431_ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a21oi_1
X_15058_ _05326_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__xnor2_1
X_14009_ _00877_ _05888_ _04182_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__a21o_1
X_18817_ _09322_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__clkbuf_1
X_09550_ _04537_ _04602_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__xor2_2
X_18748_ _03790_ net64 _09251_ vssd1 vssd1 vccd1 vccd1 _09268_ sky130_fd_sc_hd__mux2_1
X_09481_ _03848_ vssd1 vssd1 vccd1 vccd1 _03859_ sky130_fd_sc_hd__clkbuf_4
X_18679_ _02045_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09217_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ _07504_ vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__clkbuf_4
X_09748_ _05682_ vssd1 vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__inv_6
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _06008_ vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__clkbuf_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _01800_ _01801_ _01771_ _01781_ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a211o_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _00120_ _09219_ vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__nand2_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _01732_ _01731_ _01636_ _01633_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__o211a_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14360_ _02984_ _01520_ _07962_ _05964_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11572_ _01645_ _01664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _05834_ _08224_ _03417_ _03418_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_135_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput19 i_wb_addr[25] vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10523_ _00614_ _00615_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14291_ _04317_ _04327_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13242_ _00741_ _00743_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__nor2_1
X_16030_ _02988_ _03111_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10454_ _00109_ _09349_ _00171_ _00177_ vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__and4_1
X_13173_ _03270_ _00172_ _07537_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__and4b_1
X_10385_ _05649_ _07406_ _07112_ _06029_ vssd1 vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12124_ _06765_ _02214_ _02211_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__o22a_1
X_17981_ _08447_ _08419_ _08505_ vssd1 vssd1 vccd1 vccd1 _08506_ sky130_fd_sc_hd__o21a_1
X_12055_ _02143_ _02146_ _02065_ _02147_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__o211a_1
X_16932_ _06361_ _06360_ _06359_ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__a21oi_1
X_11006_ _00832_ _05617_ _01080_ _01083_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16863_ net331 _07194_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__nor2_1
X_18602_ _09113_ vssd1 vssd1 vccd1 vccd1 _09159_ sky130_fd_sc_hd__buf_2
X_15814_ _03537_ _04557_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16794_ _07114_ vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__inv_2
X_18533_ net32 net4 net3 net6 vssd1 vssd1 vccd1 vccd1 _09103_ sky130_fd_sc_hd__or4_1
X_15745_ _05947_ _05950_ _06015_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or3_1
X_12957_ _03049_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__clkbuf_4
X_11908_ _04493_ _04416_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _02001_ sky130_fd_sc_hd__and4_1
X_18464_ _03013_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _09030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15676_ _05968_ _06000_ _06001_ vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand3_1
XFILLER_0_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12888_ _02980_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__buf_4
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _07888_ _07889_ vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__xnor2_1
X_14627_ _04858_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11839_ _01928_ _01931_ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__and2_1
X_18395_ _08953_ _08954_ vssd1 vssd1 vccd1 vccd1 _08955_ sky130_fd_sc_hd__nand2_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17346_ _02972_ _07813_ _07814_ _06484_ vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14558_ _04782_ _04783_ vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13509_ _03631_ _03419_ _03635_ _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__o211ai_2
X_17277_ _07488_ _07612_ vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__and2b_1
X_14489_ _03651_ _03596_ _07004_ _06722_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__nand4_2
XFILLER_0_3_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19016_ clknet_4_9_0_clk _00001_ vssd1 vssd1 vccd1 vccd1 sel_op\[1\] sky130_fd_sc_hd__dfxtp_1
X_16228_ _06597_ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[9\].genblk1.mux.sel
+ sel_op\[0\] vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09602_ _04318_ _04766_ _05159_ _05170_ vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__a211o_2
XFILLER_0_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09533_ _04416_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__buf_6
XFILLER_0_64_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09464_ _03476_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10170_ _00261_ _00250_ _00251_ vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__or3_1
XFILLER_0_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13860_ _04018_ _04020_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__xnor2_2
X_12811_ _01470_ _01472_ _01483_ vssd1 vssd1 vccd1 vccd1 _02904_ sky130_fd_sc_hd__a21o_1
X_13791_ _03938_ _03939_ _03944_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__and3_2
XFILLER_0_97_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ _05841_ _05842_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__nor2_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _02777_ _02833_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__nand2_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _05760_ _05766_ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _02764_ _02765_ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__or2b_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _07652_ _07531_ _07653_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14412_ _04622_ _04623_ vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__and2_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _01713_ _01714_ _01715_ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__a21o_1
X_18180_ _08720_ _08721_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__nor2_1
X_15392_ _05674_ _05675_ _05692_ vssd1 vssd1 vccd1 vccd1 _05694_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17131_ _02973_ _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__nand2_1
X_11555_ _07254_ _00439_ _04384_ _07232_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__a22o_1
X_14343_ net342 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10506_ _00418_ _00421_ _00585_ _00586_ vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a211oi_2
X_14274_ _03005_ _00247_ vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17062_ _07502_ _07503_ vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _01577_ _01578_ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__and2b_1
XFILLER_0_100_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ _03326_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__xnor2_2
X_16013_ _08615_ _00399_ vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__or2_1
X_10437_ _00528_ _00527_ _00331_ _00326_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__o211a_2
XFILLER_0_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ _03248_ _03249_ _03252_ _03253_ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__o211ai_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _00460_ vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__clkbuf_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _02059_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__clkbuf_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _03028_ _02045_ vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__nor2_1
X_17964_ _07302_ _07303_ _07741_ _07861_ vssd1 vssd1 vccd1 vccd1 _08488_ sky130_fd_sc_hd__or4_2
X_10299_ _00386_ _00391_ vssd1 vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__xnor2_1
X_12038_ _02126_ _02128_ vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__nor2_1
X_16915_ _07283_ _07284_ _07344_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a21oi_2
X_17895_ _08320_ _08412_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16846_ _02973_ _07269_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__nand2_1
X_16777_ _00645_ _07105_ vssd1 vssd1 vccd1 vccd1 _07194_ sky130_fd_sc_hd__nand2_4
X_13989_ _04149_ _04150_ _04160_ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ _06200_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _09085_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15728_ _05989_ _05998_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18447_ _08915_ _08965_ _09010_ vssd1 vssd1 vccd1 vccd1 _09011_ sky130_fd_sc_hd__nor3_1
X_15659_ _05972_ _05982_ vssd1 vssd1 vccd1 vccd1 _05983_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18378_ _06405_ _06790_ _08936_ _03068_ vssd1 vssd1 vccd1 vccd1 _08937_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_44_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17329_ _03206_ _07795_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09516_ ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04242_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ _03465_ _03476_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__and2_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11340_ _01422_ _01432_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11271_ _01362_ _01363_ vssd1 vssd1 vccd1 vccd1 _01364_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13010_ _03040_ _03102_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__nand2_1
X_10222_ _05834_ _05986_ _08778_ _08768_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10153_ _00244_ _00157_ _00232_ vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__or3_1
X_14961_ _05208_ _05209_ _05222_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__a21o_1
X_10084_ _00176_ vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__buf_6
X_16700_ _06937_ _06961_ _07109_ _06542_ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__a2bb2o_1
X_13912_ _03062_ _03163_ vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__nor2_1
X_17680_ _08176_ _08177_ vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__xor2_1
X_14892_ _05147_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16631_ _07033_ _07034_ _00207_ vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o21ai_4
X_13843_ _03983_ _03984_ _04000_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16562_ _06880_ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__buf_2
X_10986_ _01020_ _01021_ _01078_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__or3_4
X_13774_ _03117_ _03927_ _03036_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__o21a_1
X_18301_ _08847_ _08852_ vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__xnor2_1
X_15513_ _05728_ _05730_ _05824_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__o21a_1
X_12725_ _02814_ _02817_ vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__nor2_1
X_16493_ _06876_ _06885_ vssd1 vssd1 vccd1 vccd1 _06886_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18232_ _07314_ _08260_ _08625_ vssd1 vssd1 vccd1 vccd1 _08779_ sky130_fd_sc_hd__or3_1
X_15444_ _03000_ _05652_ _05748_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ _02694_ _02708_ _02707_ vssd1 vssd1 vccd1 vccd1 _02749_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _01690_ _01691_ _01699_ vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__a21boi_1
X_18163_ _08701_ _08703_ vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xnor2_1
X_15375_ _05672_ _05673_ _05571_ _05629_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12587_ _02638_ _02637_ _02636_ vssd1 vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17114_ _02671_ _02842_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__or2_1
X_14326_ _04511_ _04529_ _04530_ vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__nor3_2
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11538_ _01547_ _01549_ _01546_ vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__a21o_1
X_18094_ _08624_ _08628_ vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap127 _04428_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__buf_1
X_17045_ _02188_ _06889_ vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__nand2_1
X_14257_ _04448_ _04454_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__xnor2_2
X_11469_ _01550_ _01561_ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__nor2_1
Xmax_cap138 _01843_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13208_ _00709_ _00710_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _04161_ _04335_ _04378_ _04379_ vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__a211oi_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13139_ _03226_ _03235_ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__xnor2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ clknet_4_6_0_clk _09362_ vssd1 vssd1 vccd1 vccd1 salida\[49\] sky130_fd_sc_hd__dfxtp_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _08467_ _08468_ vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__nor2_1
X_17878_ _08382_ _08287_ _08393_ vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16829_ _07157_ _07154_ vssd1 vssd1 vccd1 vccd1 _07251_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09996_ _06819_ _06873_ _09337_ _09338_ vssd1 vssd1 vccd1 vccd1 _09339_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_86_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10840_ _00916_ _00915_ _00914_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _00105_ _00117_ vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__xnor2_1
X_12510_ _02598_ _02601_ _02602_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__a21bo_1
X_13490_ _03613_ _03614_ _03610_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__a21o_1
X_12441_ _02533_ _09354_ vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15160_ _05320_ _05324_ vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__or2_1
X_12372_ _02462_ _02464_ vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14111_ _04286_ _04294_ vssd1 vssd1 vccd1 vccd1 _04295_ sky130_fd_sc_hd__xnor2_2
X_11323_ _01330_ _01332_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__or2b_1
X_15091_ _05348_ _05349_ _05363_ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__nor3_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14042_ _04004_ _04050_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__and2b_1
X_11254_ _01344_ _01345_ _01346_ vssd1 vssd1 vccd1 vccd1 _01347_ sky130_fd_sc_hd__nor3b_2
X_10205_ _00293_ _00297_ vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__xnor2_1
X_18850_ clknet_4_6_0_clk net298 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__dfxtp_1
X_11185_ _00768_ _01277_ vssd1 vssd1 vccd1 vccd1 _01278_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17801_ _08298_ _08309_ vssd1 vssd1 vccd1 vccd1 _08310_ sky130_fd_sc_hd__xnor2_1
X_10136_ _00227_ _00228_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__and2b_1
X_18781_ _09273_ _09293_ vssd1 vssd1 vccd1 vccd1 _09294_ sky130_fd_sc_hd__and2_1
X_15993_ _06339_ _06341_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__or2b_1
X_17732_ _08230_ _08231_ _08233_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__nand3_1
X_10067_ _00142_ _00159_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__xor2_2
X_14944_ _03125_ _05096_ _05099_ _03199_ _05205_ vssd1 vssd1 vccd1 vccd1 _09359_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ _07143_ _07487_ _08056_ vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__o21ai_1
X_14875_ _07635_ _05888_ _05129_ _05125_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16614_ _06940_ _06965_ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__nand2_1
X_13826_ _03786_ _03810_ _03981_ _03982_ vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__o211a_1
X_17594_ _07963_ _07955_ vssd1 vssd1 vccd1 vccd1 _08085_ sky130_fd_sc_hd__or2b_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16545_ _03313_ net150 _06805_ vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__or3_1
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13757_ _03103_ _03105_ _03090_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__mux2_1
X_10969_ _01060_ _01057_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12708_ _02776_ _02778_ _02798_ _02800_ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16476_ _06572_ _06756_ _06820_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__or3_2
X_13688_ _03811_ _03812_ _03831_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__nand3_2
XFILLER_0_122_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18215_ _02871_ _02172_ _02470_ _02851_ vssd1 vssd1 vccd1 vccd1 _08761_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15427_ _05728_ _05729_ _05634_ _05636_ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ _02693_ _02696_ _02699_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18146_ _04647_ _06445_ _03052_ vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15358_ _05654_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14309_ _04360_ _04366_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__and2b_1
XFILLER_0_151_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18077_ _08609_ _08610_ _06508_ vssd1 vssd1 vccd1 vccd1 _08611_ sky130_fd_sc_hd__o21ai_1
X_15289_ _05579_ _05580_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17028_ _06598_ _07466_ _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _07831_ _07842_ _07864_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__and3b_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _07112_ vssd1 vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__clkbuf_8
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ clknet_4_0_0_clk _09418_ vssd1 vssd1 vccd1 vccd1 salida\[32\] sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09979_ _09197_ _09205_ _07526_ _09219_ vssd1 vssd1 vccd1 vccd1 _09226_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12990_ _01248_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__clkbuf_4
X_11941_ _02032_ _02033_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel
+ _03476_ vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_98_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14660_ _04893_ _04894_ vssd1 vssd1 vccd1 vccd1 _04895_ sky130_fd_sc_hd__xor2_2
XFILLER_0_98_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11872_ _01864_ _01964_ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__nor2_1
X_13611_ _03747_ _03748_ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nand2_1
X_10823_ net229 net169 _00772_ _00129_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__nand4_2
X_14591_ _04819_ _04695_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16330_ _03089_ _02257_ _03181_ _06626_ _06708_ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__o311a_1
X_13542_ _03434_ _03586_ _03671_ _03672_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__o211ai_2
X_10754_ _00846_ _00322_ _08180_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ _03062_ _06470_ _06633_ _03913_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__a31o_1
X_13473_ _03782_ _08746_ _06613_ _03881_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__a22o_1
X_10685_ _00768_ _00776_ _00777_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__a21o_1
X_18000_ _08520_ _08522_ _08525_ _08526_ vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__nand4_1
X_15212_ _05480_ _05496_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__xnor2_1
X_12424_ _02484_ _02509_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__or2b_1
X_16192_ _03195_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15143_ _05420_ _05422_ _03536_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12355_ _02417_ _02446_ _02447_ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__nand3_2
XFILLER_0_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11306_ _00843_ _00836_ _00841_ vssd1 vssd1 vccd1 vccd1 _01399_ sky130_fd_sc_hd__and3_1
X_15074_ _05345_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__xnor2_1
X_12286_ _02264_ _02377_ _02344_ vssd1 vssd1 vccd1 vccd1 _02379_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14025_ _00106_ _01575_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__nand2_1
X_11237_ _01014_ _01016_ _01328_ net141 vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__a211oi_4
X_18902_ clknet_4_10_0_clk _00056_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[20\] sky130_fd_sc_hd__dfxtp_2
X_11168_ _01243_ _01260_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__and2_1
X_18833_ _09334_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _00211_ vssd1 vssd1 vccd1 vccd1 _00212_ sky130_fd_sc_hd__clkbuf_4
X_18764_ _09281_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__buf_1
X_11099_ _01187_ _01188_ _01191_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__nand3_4
X_15976_ _06314_ _06320_ _06322_ _02969_ vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__a31o_1
X_17715_ _08111_ _08112_ _08116_ vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__a21o_1
X_14927_ _05059_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__xnor2_1
X_18695_ _00813_ _09183_ _09191_ vssd1 vssd1 vccd1 vccd1 _09228_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17646_ _02988_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__a21o_1
X_14858_ _02989_ _04034_ _03455_ _00513_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__and4_2
X_13809_ _03800_ _03802_ vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__and2_1
X_17577_ _07106_ _07332_ _07957_ _07958_ vssd1 vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__o31a_1
X_14789_ _04892_ _04891_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__or2b_1
X_16528_ _03086_ _06851_ vssd1 vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16459_ _03920_ _06848_ vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18129_ _08665_ _08666_ vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__xnor2_1
X_09902_ _08420_ _08431_ vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__nor2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _07624_ _07679_ vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__nor2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _05181_ _06181_ _06906_ _06928_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__a211o_2
X_09695_ _04973_ _05137_ _05148_ vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__nand3_1
Xrebuffer20 _01950_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer31 _00941_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer42 _07062_ vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer53 _06232_ vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer64 _03520_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_6
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer75 _07615_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_1
Xrebuffer86 _04432_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer97 net343 vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _03476_ vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_150_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12140_ _07221_ _07243_ _00949_ _03421_ vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__and4_1
XFILLER_0_103_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12071_ _02161_ _02163_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__and2b_1
X_11022_ _00845_ _01112_ _01114_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__a21oi_4
X_15830_ _06104_ _06108_ _06166_ vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__nand3_1
X_15761_ _06091_ _06092_ vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__xor2_1
X_12973_ _03050_ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__or2_1
X_17500_ _07980_ _07981_ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__nand2_1
X_14712_ _04946_ _04951_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__nand2_1
X_11924_ _02011_ _02015_ vssd1 vssd1 vccd1 vccd1 _02017_ sky130_fd_sc_hd__xor2_1
X_18480_ _09044_ _09045_ vssd1 vssd1 vccd1 vccd1 _09046_ sky130_fd_sc_hd__nor2_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _03536_ _03912_ _04243_ vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__or3_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _02529_ _07906_ _04238_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__a21oi_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _04869_ _04876_ vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__or2_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel _03826_ vssd1 vssd1
+ vccd1 vccd1 _01948_ sky130_fd_sc_hd__and4_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _00427_ _00429_ _00428_ _00270_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17362_ _07829_ _07830_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__xnor2_2
X_14574_ _04798_ _04800_ _04667_ net126 vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__a211o_1
X_11786_ _01877_ _01878_ vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16313_ _06680_ _06684_ _06690_ vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__or3b_1
XFILLER_0_126_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13525_ cla_inst.in2\[29\] _00205_ _00171_ cla_inst.in2\[30\] vssd1 vssd1 vccd1 vccd1
+ _03655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10737_ _08104_ _08093_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__and2b_1
X_17293_ _07630_ _07332_ _07633_ _07631_ vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16244_ _06467_ _06615_ vssd1 vssd1 vccd1 vccd1 _06616_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _03180_ _03578_ _03048_ vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__mux2_1
X_10668_ _00597_ _00760_ vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12407_ _02485_ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__or2b_1
XFILLER_0_113_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16175_ _06531_ _06535_ _06540_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_140_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10599_ _00507_ _00528_ _00690_ _00691_ vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_23_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13387_ _03495_ _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 net107 vssd1 vssd1 vccd1 vccd1 o_wb_data[31] sky130_fd_sc_hd__clkbuf_4
X_15126_ _05402_ _05403_ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__xor2_2
XFILLER_0_23_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12338_ _02426_ _02429_ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _05111_ _05221_ _05327_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__a21bo_1
X_12269_ _07352_ _00563_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__nand2_1
X_14008_ _00877_ _01678_ _04182_ vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__nand3_1
XFILLER_0_37_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18816_ _09298_ _09321_ vssd1 vssd1 vccd1 vccd1 _09322_ sky130_fd_sc_hd__and2_1
X_18747_ _09267_ vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__buf_1
X_15959_ _06304_ _06305_ vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_616 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09480_ cla_inst.in2\[16\] vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__clkbuf_4
X_18678_ net39 _09189_ _09216_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17629_ _08121_ _08122_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09816_ cla_inst.in2\[29\] vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__clkbuf_4
X_09747_ _06678_ vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__inv_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ ApproximateM_inst.lob_16.lob2.genblk1\[7\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _06008_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _01633_ _01636_ _01731_ _01732_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11571_ _00832_ _00439_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13310_ _05224_ _08169_ _03417_ _03418_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__and4_2
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _03728_ _05486_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ _04376_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10453_ _00125_ _00218_ _00178_ _00151_ vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22oi_1
X_13241_ _03341_ _03342_ _00696_ _03204_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10384_ _05736_ _08224_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__nand2_1
X_13172_ _07504_ _00178_ _00147_ _00358_ vssd1 vssd1 vccd1 vccd1 _03271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _06040_ _00194_ _02215_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__a21oi_2
X_17980_ _08410_ _08504_ vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _02023_ _02063_ _02064_ vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__o21ai_1
X_16931_ _07356_ _07357_ _07360_ vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a21o_1
X_11005_ _04580_ _01064_ _01063_ _01066_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__o2bb2a_1
X_16862_ _07196_ _07197_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15813_ _04823_ _06140_ _06141_ _06142_ _06150_ vssd1 vssd1 vccd1 vccd1 _09371_ sky130_fd_sc_hd__a32o_1
X_18601_ _09097_ vssd1 vssd1 vccd1 vccd1 _09157_ sky130_fd_sc_hd__buf_2
X_16793_ _07209_ _07211_ vssd1 vssd1 vccd1 vccd1 _07212_ sky130_fd_sc_hd__xor2_1
X_18532_ net14 net17 net16 net19 vssd1 vssd1 vccd1 vccd1 _09102_ sky130_fd_sc_hd__or4_1
X_15744_ _05411_ _05415_ _05792_ _06075_ vssd1 vssd1 vccd1 vccd1 _06076_ sky130_fd_sc_hd__a211o_1
X_12956_ _03048_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__clkbuf_4
X_18463_ _06425_ _06451_ _09028_ vssd1 vssd1 vccd1 vccd1 _09029_ sky130_fd_sc_hd__or3_1
X_11907_ _01987_ _01989_ _01988_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__o21ai_1
X_15675_ _05998_ _05999_ _05912_ _05969_ vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _00494_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__buf_4
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _06750_ _07623_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _04855_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _01851_ _01930_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__nor2_1
X_18394_ _08848_ _08899_ _08901_ vssd1 vssd1 vccd1 vccd1 _08954_ sky130_fd_sc_hd__o21ai_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _02978_ _06999_ _02972_ vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__o21ai_1
X_14557_ _00148_ _00149_ _06471_ _08452_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11769_ _08452_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _03632_ _03633_ _03634_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17276_ _07629_ _07736_ _07737_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__o21ai_1
X_14488_ _03377_ _07004_ cla_inst.in1\[24\] _03356_ vssd1 vssd1 vccd1 vccd1 _04707_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19015_ clknet_4_9_0_clk _00000_ vssd1 vssd1 vccd1 vccd1 sel_op\[0\] sky130_fd_sc_hd__dfxtp_2
X_16227_ _02965_ _06418_ _06419_ vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__a21o_1
X_13439_ _03152_ _03127_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__or2_1
XFILLER_0_140_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16158_ _06518_ _06521_ _03313_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__a21o_2
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15109_ _05367_ _05383_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16089_ _04900_ _06446_ vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__and2_1
X_09601_ _04973_ _05148_ _05137_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a21oi_2
X_09532_ ApproximateM_inst.lob_16.lob2.genblk1\[12\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04416_ sky130_fd_sc_hd__buf_6
X_09463_ _03366_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12810_ _02901_ _02902_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__nor2_1
X_13790_ _03942_ _03943_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _02777_ _02833_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__xor2_2
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _05760_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__or2_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12672_ _02759_ _02760_ vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _04610_ _04611_ _04621_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__or3_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _01713_ _01714_ _01715_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nand3_2
XFILLER_0_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15391_ _05690_ _05691_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17130_ _02978_ _06843_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__or2_1
X_14342_ _04420_ _04397_ _04546_ _04547_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__a211o_4
X_11554_ _07232_ _07254_ _00439_ _04384_ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__nand4_2
XFILLER_0_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10505_ _00559_ _00574_ vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__or2b_1
X_17061_ _07393_ _07399_ _07501_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__and3_1
X_14273_ _04301_ _04311_ vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__and2_1
X_11485_ _05595_ _04886_ _03815_ _05573_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16012_ _06359_ _06360_ _06361_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a21bo_1
X_13224_ _00107_ _00166_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__nand2_1
X_10436_ _00326_ _00331_ _00527_ _00528_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13155_ _08724_ _08158_ _03250_ _03251_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__a22o_1
X_10367_ _00459_ vssd1 vssd1 vccd1 vccd1 _00460_ sky130_fd_sc_hd__buf_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _02197_ _02183_ _02187_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__nand3_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _00389_ _00390_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__nor2_1
X_13086_ _03172_ _03177_ _03060_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__mux2_1
X_17963_ _07207_ _07745_ _07859_ _06947_ vssd1 vssd1 vccd1 vccd1 _08487_ sky130_fd_sc_hd__a22o_1
X_12037_ _00845_ _02124_ _02125_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__a21oi_2
X_16914_ _07342_ _07343_ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__xor2_1
X_17894_ _08410_ _08411_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__or2_1
X_16845_ _02978_ _06617_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__or2_1
X_16776_ _07111_ _07137_ vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__or2_1
X_13988_ _04149_ _04150_ _04160_ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15727_ _06055_ _06056_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or2_1
X_18515_ _06246_ _06452_ vssd1 vssd1 vccd1 vccd1 _09084_ sky130_fd_sc_hd__or2_1
X_12939_ _03024_ _03031_ vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15658_ _05980_ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__nor2_1
X_18446_ _09007_ _09009_ vssd1 vssd1 vccd1 vccd1 _09010_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14609_ _01521_ _07015_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__nand4_4
XFILLER_0_145_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18377_ _02992_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _08936_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15589_ _05905_ _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17328_ _07792_ _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_154_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17259_ _07607_ _07609_ _07610_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09515_ _03454_ _04220_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ ApproximateM_inst.lob_16.lob1.genblk1\[9\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03476_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _01355_ _01361_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__and2_1
X_10221_ _00310_ _00313_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10152_ _00157_ _00232_ _00244_ vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__o21ai_2
X_14960_ _05111_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__xnor2_1
X_10083_ ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00176_ sky130_fd_sc_hd__buf_4
X_13911_ _03147_ _03159_ _03061_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__mux2_1
X_14891_ _00106_ _06094_ _05145_ _05146_ vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__and4_1
X_16630_ _01005_ _03184_ _06871_ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__a21oi_2
X_13842_ _03983_ _03984_ _04000_ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__nor3_2
X_16561_ _06952_ _06958_ vssd1 vssd1 vccd1 vccd1 _06959_ sky130_fd_sc_hd__xor2_1
X_13773_ _03913_ _03926_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10985_ _01053_ _01077_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15512_ _05767_ _05822_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__xnor2_1
X_18300_ _08849_ _08850_ _08851_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__and3_1
X_12724_ _02791_ _02816_ vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16492_ _06882_ _06883_ vssd1 vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18231_ _07650_ _07708_ vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__nand2_1
X_15443_ _03000_ _05652_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__nand3_1
XFILLER_0_128_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12655_ _02747_ _02666_ vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11606_ _01694_ _01697_ _01698_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__or3b_1
X_18162_ _06368_ _07390_ vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15374_ _05571_ _05629_ _05672_ _05673_ vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__a211o_1
X_12586_ _07591_ _02676_ _02677_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17113_ _07556_ _07557_ _07560_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__o21a_1
X_14325_ _04369_ _04372_ _04528_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__and3_1
XFILLER_0_135_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11537_ _01625_ _01626_ _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__nand3_2
X_18093_ _08625_ _08627_ vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__xor2_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ _06756_ _07318_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__or2_1
X_14256_ _04452_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__or2_1
X_11468_ _01551_ _01560_ vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__xnor2_1
Xmax_cap128 _02383_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
X_13207_ _00708_ _00707_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10419_ _00510_ _00511_ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__or2_1
X_14187_ _04376_ _04377_ _04354_ vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__a21oi_2
X_11399_ _01415_ _01454_ _01490_ _01491_ vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__o211a_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _03233_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__and2b_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ clknet_4_6_0_clk _09361_ vssd1 vssd1 vccd1 vccd1 salida\[48\] sky130_fd_sc_hd__dfxtp_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _02983_ vssd1 vssd1 vccd1 vccd1 _03161_ sky130_fd_sc_hd__buf_4
X_17946_ _08359_ net132 _08466_ vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__o21a_1
X_17877_ _08391_ _08392_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__and2_1
X_16828_ _07248_ _07249_ vssd1 vssd1 vccd1 vccd1 _07250_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16759_ _07173_ _06420_ _07174_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18429_ _06408_ _08991_ vssd1 vssd1 vccd1 vccd1 _08992_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09995_ _09152_ _09158_ _09333_ vssd1 vssd1 vccd1 vccd1 _09338_ sky130_fd_sc_hd__nor3_4
XFILLER_0_79_530 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ _00122_ _00862_ vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09429_ _03239_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12440_ _05834_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__buf_6
XFILLER_0_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12371_ _02397_ _02463_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ _04287_ _04293_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11322_ _01312_ _01378_ _01413_ _01414_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__a211oi_4
X_15090_ _05348_ _05349_ _05363_ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__o21a_1
X_14041_ _04169_ _04170_ _04216_ _04217_ vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__o22a_1
X_11253_ _01254_ _01256_ _01255_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _00295_ _00296_ vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__and2b_1
X_11184_ _00777_ _00776_ vssd1 vssd1 vccd1 vccd1 _01277_ sky130_fd_sc_hd__and2b_1
X_17800_ _08307_ _08308_ vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__nor2_1
X_10135_ _00226_ _00202_ _00209_ vssd1 vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__or3_1
X_18780_ _02988_ net43 _09276_ vssd1 vssd1 vccd1 vccd1 _09293_ sky130_fd_sc_hd__mux2_1
X_15992_ _03790_ _00207_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__or2_1
X_10066_ _00157_ _00158_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__or2_1
X_14943_ _05198_ _05202_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__o21a_1
X_17731_ _08230_ _08231_ _08233_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__a21o_1
X_14874_ _05127_ vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17662_ _08155_ _08157_ vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__xor2_1
X_13825_ _03981_ _03982_ _03786_ net189 vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__a211oi_2
X_16613_ _03169_ _06464_ _06987_ _07016_ vssd1 vssd1 vccd1 vccd1 _09414_ sky130_fd_sc_hd__o2bb2a_2
X_17593_ _07979_ _07989_ _07987_ vssd1 vssd1 vccd1 vccd1 _08084_ sky130_fd_sc_hd__a21o_1
X_16544_ _06876_ _06885_ vssd1 vssd1 vccd1 vccd1 _06941_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ _03906_ _03907_ _02980_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__mux2_1
X_10968_ _01057_ _01060_ vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12707_ _02762_ _02799_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__xor2_2
X_16475_ _06828_ _06831_ vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__and2b_1
X_13687_ _03811_ _03812_ _03831_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ _06008_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15426_ _05634_ _05636_ _05728_ _05729_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18214_ _08759_ _02871_ vssd1 vssd1 vccd1 vccd1 _08760_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12638_ _02727_ _02730_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15357_ _00190_ _00192_ _07744_ _08224_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__and4_1
X_18145_ _06598_ _08683_ _08684_ vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__or3_1
X_12569_ _02654_ _02660_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__and3_1
XFILLER_0_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14308_ _04509_ _04510_ vssd1 vssd1 vccd1 vccd1 _04511_ sky130_fd_sc_hd__xor2_4
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18076_ _08513_ _08514_ _08512_ vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__a21boi_2
X_15288_ _01505_ _00339_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _01041_ _06364_ _06363_ vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14239_ net201 _04433_ _04270_ _04271_ vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_150_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _07102_ vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__buf_6
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ clknet_4_3_0_clk _09410_ vssd1 vssd1 vccd1 vccd1 salida\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _08378_ _08379_ vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__and2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09978_ _09212_ vssd1 vssd1 vccd1 vccd1 _09219_ sky130_fd_sc_hd__buf_4
X_11940_ _05638_ _03421_ _03607_ _00992_ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_98_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11871_ _07711_ _01962_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__and3_2
X_13610_ _03741_ _03746_ _02969_ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__a21oi_1
X_10822_ net169 _00772_ _00129_ net227 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__a22o_1
X_14590_ _04688_ _04689_ vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13541_ _03649_ _03650_ _03670_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__or3_4
XFILLER_0_95_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10753_ _00845_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _01746_ _01503_ _03083_ _03166_ _06477_ _03161_ vssd1 vssd1 vccd1 vccd1 _06633_
+ sky130_fd_sc_hd__mux4_1
X_13472_ _03593_ _03594_ _03591_ _03592_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__o211ai_2
X_10684_ _00771_ _00775_ _00769_ _00770_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__o211a_1
X_15211_ _05494_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__xor2_2
XFILLER_0_124_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _02482_ vssd1 vssd1 vccd1 vccd1 _02516_ sky130_fd_sc_hd__inv_2
X_16191_ _03029_ _06464_ _06465_ _06557_ vssd1 vssd1 vccd1 vccd1 _09386_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15142_ _04254_ _04258_ _02780_ vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__mux2_1
X_12354_ _02443_ _02444_ _02433_ _02441_ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11305_ _00846_ _00119_ _00121_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__a21oi_2
X_15073_ _05227_ _05239_ _05226_ vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ _02264_ _02344_ _02377_ vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14024_ _04199_ _04200_ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__nor2_1
X_18901_ clknet_4_12_0_clk _00055_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[19\] sky130_fd_sc_hd__dfxtp_2
X_11236_ _01315_ _01327_ _01316_ _01318_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__nor4_1
X_18832_ net46 _03217_ _09331_ vssd1 vssd1 vccd1 vccd1 _09334_ sky130_fd_sc_hd__mux2_1
X_11167_ _01253_ _01259_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__xnor2_1
X_10118_ _00210_ vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__clkbuf_8
X_18763_ _09273_ _09280_ vssd1 vssd1 vccd1 vccd1 _09281_ sky130_fd_sc_hd__and2_1
X_11098_ _01189_ _01190_ vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__xnor2_4
X_15975_ _06314_ _06320_ _06322_ vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__a21oi_1
X_17714_ _08214_ _08215_ vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__xnor2_1
X_14926_ _05184_ _05185_ vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__xnor2_1
X_10049_ _00124_ _00137_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__nand2_2
X_18694_ net47 _09189_ _09227_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17645_ _08036_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__clkbuf_4
X_14857_ _04034_ _03456_ _00665_ _02989_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__a22oi_4
X_13808_ _03961_ _03962_ net236 _03931_ vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__a211o_4
X_17576_ _08063_ _08064_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__or2b_1
X_14788_ _05016_ _04917_ _05033_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__nor3_1
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13739_ net121 _03885_ _03887_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16527_ _06346_ _06790_ _06922_ _03086_ vssd1 vssd1 vccd1 vccd1 _06923_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16458_ _06469_ _06476_ _06498_ _06473_ _03079_ _03077_ vssd1 vssd1 vccd1 vccd1 _06848_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ _05614_ _05618_ _05612_ vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16389_ _06664_ _06772_ _06654_ vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18128_ _08577_ _08580_ _08576_ vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18059_ _06559_ _08590_ vssd1 vssd1 vccd1 vccd1 _08591_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09901_ _03859_ _04121_ _04460_ _04482_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__and4_1
XFILLER_0_6_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _07635_ _07646_ _07657_ _07668_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_67_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _06863_ _06873_ _06917_ _06548_ vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__o2bb2a_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _05181_ _06149_ _06159_ _06170_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__nand4_4
Xrebuffer10 _04094_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_1
Xrebuffer21 _00305_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__dlygate4sd1_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer32 net194 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__buf_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer43 _00772_ vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_2
Xrebuffer54 _04681_ vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_1
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer65 net227 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer76 _04003_ vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer87 _06560_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12070_ _02053_ _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__xnor2_1
X_11021_ _01113_ _06776_ vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__nor2_4
XFILLER_0_99_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15760_ _03015_ _03072_ vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__nand2_1
X_12972_ _09263_ _03064_ _03024_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14711_ _04410_ _04947_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__a21o_1
X_11923_ _02011_ _02015_ vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__and2_1
X_15691_ _06015_ _06016_ _04823_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _04872_ _04874_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__or2_1
X_17430_ _02589_ _02844_ _02587_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__o21ba_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ ApproximateM_inst.lob_16.lob2.genblk1\[3\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel
+ _03826_ ApproximateM_inst.lob_16.lob2.genblk1\[4\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _01947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _00893_ _00895_ _00897_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__nand3_2
X_14573_ _04667_ net126 _04798_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__o211ai_4
X_17361_ net331 _07706_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11785_ _01508_ _01513_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13524_ cla_inst.in2\[30\] cla_inst.in2\[29\] _00205_ _00171_ vssd1 vssd1 vccd1 vccd1
+ _03654_ sky130_fd_sc_hd__and4_1
X_16312_ _06687_ _06597_ _06688_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__or3_1
X_10736_ _00827_ _00828_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__nand2_1
X_17292_ _07753_ _07754_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16243_ _06612_ _06614_ _02982_ vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13455_ _03187_ vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__inv_2
X_10667_ _00594_ _00596_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ _02491_ _02498_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16174_ _06536_ _06538_ _06539_ _03313_ _06520_ vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__a2111o_1
X_13386_ _03496_ _03502_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ _00688_ _00689_ _00482_ _00487_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15125_ _03368_ _03067_ _05278_ _05276_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a31o_1
Xoutput108 net108 vssd1 vssd1 vccd1 vccd1 o_wb_data[3] sky130_fd_sc_hd__clkbuf_4
X_12337_ _02426_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15056_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12268_ _02357_ _02360_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__nor2_1
X_14007_ _04180_ _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ net220 _01020_ _01310_ _01311_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__o211ai_4
X_12199_ _02288_ _02289_ _02203_ vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__a21oi_1
Xoutput90 net90 vssd1 vssd1 vccd1 vccd1 o_wb_data[16] sky130_fd_sc_hd__clkbuf_4
X_18815_ _03016_ net55 _09301_ vssd1 vssd1 vccd1 vccd1 _09321_ sky130_fd_sc_hd__mux2_1
X_18746_ _09245_ _09266_ vssd1 vssd1 vccd1 vccd1 _09267_ sky130_fd_sc_hd__and2_1
X_15958_ _06272_ _06280_ _06278_ vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__o21ai_1
X_14909_ _05165_ _05166_ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__xnor2_1
X_18677_ _02127_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09216_ sky130_fd_sc_hd__a21oi_1
X_15889_ _06183_ _06225_ vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__or2_1
X_17628_ _08016_ _08018_ _08014_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__o21ba_1
X_17559_ _06655_ _07825_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09815_ _07472_ _07210_ _07319_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__nand3_2
X_09746_ _06678_ _06700_ _06711_ _06732_ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__and4b_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _05747_ _05986_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__nand2_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _04056_ net204 _01660_ _01662_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ _00443_ _00612_ _00613_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13240_ _00696_ _03204_ _03341_ _03342_ vssd1 vssd1 vccd1 vccd1 _03343_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ _07526_ _00132_ _00360_ _00359_ _07570_ vssd1 vssd1 vccd1 vccd1 _00545_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13171_ _09166_ _09172_ _00178_ _00181_ vssd1 vssd1 vccd1 vccd1 _03270_ sky130_fd_sc_hd__and4_1
X_10383_ _00474_ _00475_ vssd1 vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12122_ _06051_ _00172_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__and2_1
XFILLER_0_103_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12053_ _02144_ _02145_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__and2_1
X_16930_ _07356_ _07357_ _07360_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__nand3_1
X_11004_ _01094_ _01096_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__nand2_2
X_16861_ _06937_ _07130_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__nor2_1
X_18600_ net265 _09140_ _09156_ _09144_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__o211a_1
X_15812_ _03121_ _06148_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__nand2_1
X_16792_ _07018_ _06875_ vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__nor2_1
X_18531_ net18 net21 net20 net22 vssd1 vssd1 vccd1 vccd1 _09100_ sky130_fd_sc_hd__or4b_1
X_15743_ _05948_ _05875_ _05947_ _06015_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__or4_1
X_12955_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__clkbuf_4
X_11906_ _01997_ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__or2_1
X_18462_ _06408_ _06449_ _03073_ vssd1 vssd1 vccd1 vccd1 _09028_ sky130_fd_sc_hd__a21oi_1
X_15674_ _05912_ _05969_ _05998_ _05999_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12886_ _02978_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__clkbuf_4
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _07885_ _07887_ vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _04725_ _03455_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__and3_1
X_11837_ _06711_ _04045_ _01929_ _01850_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__a22oi_1
X_18393_ _08950_ _08952_ vssd1 vssd1 vccd1 vccd1 _08953_ sky130_fd_sc_hd__xor2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _03321_ _06471_ _04591_ _03322_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_23_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17344_ _06696_ _06701_ _06703_ _06707_ _03061_ _03079_ vssd1 vssd1 vccd1 vccd1 _07813_
+ sky130_fd_sc_hd__mux4_1
X_11768_ _01859_ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13507_ _03632_ _03633_ _03634_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10719_ _08060_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__inv_2
X_14487_ _01521_ _07962_ _04568_ _04570_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__and4_1
XFILLER_0_70_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17275_ _07637_ _07638_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__or2_1
X_11699_ _01764_ _01765_ _01767_ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_130_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19014_ clknet_4_3_0_clk _00104_ vssd1 vssd1 vccd1 vccd1 op_code\[3\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13438_ _03532_ _03559_ vssd1 vssd1 vccd1 vccd1 _09377_ sky130_fd_sc_hd__nand2_1
X_16226_ _02784_ _06333_ _03030_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_125_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer1 _00694_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__buf_1
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16157_ _03281_ _06519_ _06520_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13369_ _03482_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15108_ _05367_ _05383_ vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__nand2_1
X_16088_ _03052_ _04647_ _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__and3_1
X_15039_ _02976_ _03039_ _05306_ _05307_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__o32a_1
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09600_ _04973_ _05137_ _05148_ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ _04351_ _04373_ _04384_ _04395_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__and4_4
X_18729_ _09253_ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09462_ _03531_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__buf_8
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09729_ _05006_ _05104_ vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _02801_ _02831_ _02832_ vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a21o_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _08865_ _01357_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__nand2_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _04610_ _04611_ _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__o21ai_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11622_ _01625_ _01630_ vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15390_ _05536_ _05547_ _05534_ vssd1 vssd1 vccd1 vccd1 _05691_ sky130_fd_sc_hd__a21oi_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14341_ _04544_ _04545_ _04350_ _04422_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__o211a_1
X_11553_ _01643_ _01645_ vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ _00594_ _00596_ vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__or2_1
X_17060_ _07393_ _07399_ _07501_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__a21oi_1
X_14272_ _04468_ _04469_ _04299_ _04428_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a211o_2
XFILLER_0_123_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ _05573_ _05595_ _04886_ _03815_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16011_ _00644_ _00248_ vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13223_ _03323_ _03325_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__nor2_1
X_10435_ _00507_ _00508_ _00526_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__nor3_4
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13154_ _08724_ _08158_ _03250_ _03251_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__nand4_4
X_10366_ _06613_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__clkbuf_8
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _02183_ _02187_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__a21o_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _03174_ _03176_ _03047_ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__mux2_1
X_17962_ _08367_ _08375_ _08373_ vssd1 vssd1 vccd1 vccd1 _08486_ sky130_fd_sc_hd__a21o_1
X_10297_ cla_inst.in2\[25\] _00172_ _00387_ _00388_ vssd1 vssd1 vccd1 vccd1 _00390_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_20_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12036_ _02126_ _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__and2_1
X_16913_ _07233_ _07234_ _07237_ vssd1 vssd1 vccd1 vccd1 _07343_ sky130_fd_sc_hd__a21o_1
X_17893_ _08314_ _08347_ _08408_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__and3_1
X_16844_ _03912_ _06629_ _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16775_ _07152_ _07153_ vssd1 vssd1 vccd1 vccd1 _07192_ sky130_fd_sc_hd__and2b_1
X_13987_ _04158_ _04159_ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _06248_ _06414_ _09076_ vssd1 vssd1 vccd1 vccd1 _09083_ sky130_fd_sc_hd__or3b_1
X_15726_ _05917_ _06054_ vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__nor2_1
X_12938_ _03027_ _01746_ _03030_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18445_ _08961_ _09008_ vssd1 vssd1 vccd1 vccd1 _09009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15657_ _05978_ _05979_ _05973_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__a21oi_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _02958_ _02960_ _02961_ vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__a21oi_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14608_ _03651_ _03596_ cla_inst.in1\[27\] _07112_ vssd1 vssd1 vccd1 vccd1 _04838_
+ sky130_fd_sc_hd__nand4_4
X_18376_ _03068_ _06448_ vssd1 vssd1 vccd1 vccd1 _08935_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15588_ _05903_ _05904_ _05815_ _05817_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__o211a_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17327_ _07671_ _07558_ _07670_ _07793_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__o31a_4
X_14539_ _01504_ _06094_ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _07705_ _07717_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16209_ _06574_ _06576_ _03324_ vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a21o_1
X_17189_ _07619_ _07642_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09514_ ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04220_ sky130_fd_sc_hd__buf_6
XFILLER_0_149_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _03454_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_870 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _00311_ _00312_ vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__and2b_1
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _00233_ _00243_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _00174_ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__clkbuf_4
X_13910_ _02978_ _04075_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__nor2_1
X_14890_ _00148_ _00149_ _00459_ _05845_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__nand4_2
XFILLER_0_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13841_ _03985_ _03999_ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16560_ _06522_ _06525_ _06957_ _00515_ vssd1 vssd1 vccd1 vccd1 _06958_ sky130_fd_sc_hd__a211o_1
X_13772_ _03033_ _03924_ _03099_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__mux2_1
X_10984_ _01053_ _01074_ _01075_ _01076_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__and4b_1
XFILLER_0_85_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15511_ _05811_ _05821_ vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__xor2_1
XFILLER_0_139_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12723_ _02789_ _02815_ vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16491_ _06578_ _06816_ vssd1 vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18230_ _08774_ _08775_ vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__nand2_1
X_15442_ _05745_ _05746_ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__xnor2_1
X_12654_ _02611_ _02654_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11605_ _07853_ _01695_ _01696_ _01673_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__a31o_2
XFILLER_0_26_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18161_ _08699_ _08700_ vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__and2b_1
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15373_ _05651_ _05670_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__and2_1
X_12585_ _07243_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel ApproximateM_inst.lob_16.lob1.mux.sel
+ _07221_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17112_ _06559_ _07558_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__nor2_1
X_14324_ _04369_ _04372_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a21oi_2
X_11536_ _01627_ _01628_ vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18092_ _07332_ _08260_ _08459_ vssd1 vssd1 vccd1 vccd1 _08627_ sky130_fd_sc_hd__or3_1
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14255_ _06460_ _00502_ _04450_ _04451_ vssd1 vssd1 vccd1 vccd1 _04453_ sky130_fd_sc_hd__o2bb2a_1
X_17043_ _07392_ _07404_ vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap118 _05863_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_1
X_11467_ _01556_ _01559_ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap129 _02293_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_1
XFILLER_0_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13206_ _03305_ _03306_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10418_ cla_inst.in2\[31\] _07700_ _00509_ _07559_ vssd1 vssd1 vccd1 vccd1 _00511_
+ sky130_fd_sc_hd__and4_1
XFILLER_0_110_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14186_ _04354_ _04376_ _04377_ vssd1 vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__and3_2
X_11398_ _01468_ _01489_ _01488_ vssd1 vssd1 vccd1 vccd1 _01491_ sky130_fd_sc_hd__a21o_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _03231_ _03232_ _03227_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__a21o_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _03793_ _00440_ _00441_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__a21bo_1
X_18994_ clknet_4_0_0_clk _09360_ vssd1 vssd1 vccd1 vccd1 salida\[47\] sky130_fd_sc_hd__dfxtp_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _03159_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__inv_2
X_17945_ _08359_ net132 _08466_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__nor3_1
X_12019_ _05562_ _05584_ _04220_ _04242_ vssd1 vssd1 vccd1 vccd1 _02112_ sky130_fd_sc_hd__and4_1
X_17876_ _08389_ _08390_ vssd1 vssd1 vccd1 vccd1 _08392_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16827_ _07191_ _07192_ _07247_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16758_ _07172_ _06355_ _06354_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__a21o_1
X_15709_ _01417_ _00665_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16689_ _07096_ _07097_ _07098_ vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18428_ _03016_ _06592_ _06551_ vssd1 vssd1 vccd1 vccd1 _08991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18359_ _08862_ _08894_ _08914_ vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__or3_1
XFILLER_0_145_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09994_ _09152_ _09158_ _09333_ vssd1 vssd1 vccd1 vccd1 _09337_ sky130_fd_sc_hd__o21a_2
XFILLER_0_79_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09428_ sel_op\[1\] vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12370_ _02311_ _02396_ _02392_ _02395_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11321_ _01394_ _01395_ _01412_ vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_132_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _04169_ _04170_ _04216_ _04217_ vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__nor4_2
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11252_ _00169_ _00131_ _01342_ _01343_ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _00294_ _05322_ _05333_ _04504_ vssd1 vssd1 vccd1 vccd1 _00296_ sky130_fd_sc_hd__a22o_1
X_11183_ _00965_ _00961_ vssd1 vssd1 vccd1 vccd1 _01276_ sky130_fd_sc_hd__or2b_4
XFILLER_0_101_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10134_ _00202_ _00209_ _00226_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__o21a_1
X_15991_ _03790_ _00207_ vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__and2_1
X_17730_ _08025_ _08026_ _08132_ _08232_ vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__a31o_1
X_10065_ _08202_ _00143_ _00156_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__nor3_1
X_14942_ _05198_ _05202_ _04238_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a21oi_1
X_17661_ _08156_ _08051_ _08048_ vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__a21o_1
X_14873_ _05125_ _05888_ _07635_ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__and4b_1
X_16612_ _06992_ _06994_ _07011_ _07014_ vssd1 vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__a211o_1
X_13824_ _03963_ _03964_ _03980_ vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__nand3_2
X_17592_ _08079_ _08081_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16543_ _06937_ _06766_ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__nor2_1
X_10967_ _01058_ _01059_ vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__xnor2_4
X_13755_ _03110_ _03113_ _03090_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12706_ _02774_ _02773_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__and2b_1
X_16474_ _03166_ _06464_ _06865_ vssd1 vssd1 vccd1 vccd1 _09412_ sky130_fd_sc_hd__a21oi_2
X_13686_ _03814_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__xnor2_1
X_10898_ _05682_ _05388_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _02172_ _02470_ _02851_ vssd1 vssd1 vccd1 vccd1 _08759_ sky130_fd_sc_hd__nor3_1
X_15425_ _05720_ _05727_ vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ _02600_ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18144_ _08682_ _06397_ _06396_ vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15356_ _02996_ _00339_ _09059_ _02993_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_53_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12568_ _02534_ _02537_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14307_ _01873_ _03044_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__nand2_2
X_11519_ _04690_ _03673_ _01172_ _01173_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18075_ _08607_ _08608_ vssd1 vssd1 vccd1 vccd1 _08609_ sky130_fd_sc_hd__nand2_1
X_15287_ _05577_ _05578_ vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__nor2_1
X_12499_ _02582_ _02591_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17026_ _01041_ _06363_ _06364_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__and3_1
X_14238_ _04270_ _04271_ net200 _04433_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _00115_ _02124_ _04201_ _04200_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__a31o_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ clknet_4_6_0_clk _09409_ vssd1 vssd1 vccd1 vccd1 salida\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17928_ _08405_ _08407_ vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__and2b_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17859_ _08269_ _08271_ _08372_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09977_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _09212_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11870_ _00515_ _01862_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__nor2_2
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10821_ cla_inst.in2\[18\] _00179_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__and2_1
X_13540_ _03649_ _03650_ _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__o21ai_2
X_10752_ _07711_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__buf_4
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13471_ _03591_ _03592_ _03593_ _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__a211o_1
X_10683_ _00769_ _00770_ _00771_ _00775_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15210_ _01873_ _03071_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__nand2_1
X_12422_ _02448_ _02513_ _02514_ vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__and3_1
X_16190_ _06481_ _06484_ _06506_ _06556_ vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15141_ _02977_ _02980_ _03560_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__or3_1
X_12353_ _02445_ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11304_ _00122_ _00862_ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15072_ _05342_ _05343_ vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__nand2_1
X_12284_ _02261_ _02262_ _02263_ _02256_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14023_ cla_inst.in2\[27\] _09349_ _04657_ _04864_ vssd1 vssd1 vccd1 vccd1 _04200_
+ sky130_fd_sc_hd__and4_1
X_18900_ clknet_4_10_0_clk _00054_ vssd1 vssd1 vccd1 vccd1 cla_inst.in1\[18\] sky130_fd_sc_hd__dfxtp_2
X_11235_ _01315_ _01316_ _01318_ _01327_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__o31a_1
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18831_ _09332_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__clkbuf_1
X_11166_ _01241_ _01258_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10117_ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00210_ sky130_fd_sc_hd__buf_4
X_18762_ _08615_ net37 _09276_ vssd1 vssd1 vccd1 vccd1 _09280_ sky130_fd_sc_hd__mux2_1
X_11097_ _01123_ _01122_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__and2b_1
X_15974_ _06271_ _06307_ _06321_ vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__and3_1
X_17713_ _07978_ _08105_ _08108_ vssd1 vssd1 vccd1 vccd1 _08215_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14925_ _05014_ _05063_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__nand2_1
X_10048_ _00118_ _00139_ _00140_ vssd1 vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__a21oi_2
X_18693_ _01692_ _09183_ _09191_ vssd1 vssd1 vccd1 vccd1 _09227_ sky130_fd_sc_hd__a21oi_1
Xhold90 _00009_ vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17644_ _06425_ _06442_ _08139_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__or3_1
X_14856_ _05106_ _05108_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13807_ net236 _03931_ _03961_ _03962_ vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__o211ai_4
X_17575_ _08043_ _08044_ _08062_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__or3b_1
X_14787_ _05016_ _04917_ _05033_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__o21a_1
X_11999_ _02014_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16526_ _03036_ _06920_ _06921_ vssd1 vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__a21o_1
X_13738_ net121 _03885_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__nor3_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16457_ _06843_ _06846_ _03080_ vssd1 vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__mux2_1
X_13669_ _03809_ net326 _03622_ _03752_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_6_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15408_ _05710_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16388_ _06572_ _06664_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18127_ _08662_ _08664_ vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__xnor2_1
X_15339_ _09353_ _07025_ _05633_ _05634_ vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18058_ _08586_ _08589_ vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _03793_ _04460_ _08409_ _03859_ vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__a22oi_2
X_17009_ _07379_ _07380_ _07445_ _07446_ vssd1 vssd1 vccd1 vccd1 _07447_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _07515_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__clkbuf_4
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _06526_ _06537_ _04973_ _06191_ vssd1 vssd1 vccd1 vccd1 _06917_ sky130_fd_sc_hd__o211a_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _05159_ _05170_ _04318_ _04766_ vssd1 vssd1 vccd1 vccd1 _06170_ sky130_fd_sc_hd__o211ai_4
Xrebuffer11 net173 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__clkbuf_1
Xrebuffer22 _00772_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer33 _04741_ vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer44 net206 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer55 _04152_ vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer66 net227 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer77 _03376_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer88 _04458_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11020_ _00514_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__clkbuf_8
X_12971_ _03028_ _00516_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__nor2_1
X_14710_ _04817_ _04948_ _04949_ vssd1 vssd1 vccd1 vccd1 _04950_ sky130_fd_sc_hd__nand3_4
X_11922_ _02012_ _02014_ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__or2_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _06015_ _06016_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__and2_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _03014_ _05921_ _04873_ _04870_ vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__o2bb2a_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ _01848_ _01856_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__xnor2_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _00896_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__inv_2
X_17360_ _07824_ _07826_ _07827_ _07828_ vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__o22a_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14572_ _04796_ _04797_ _04622_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__o21ai_2
X_11784_ _01825_ _01824_ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16311_ _06685_ _06332_ _06686_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__a21oi_1
X_13523_ _03005_ _00223_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nand2_1
X_10735_ _00826_ _00825_ _00818_ _00801_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__o211ai_1
X_17291_ _06875_ _07318_ vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16242_ _07810_ _03069_ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10666_ _00757_ _00758_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__nor2_2
X_13454_ _03575_ _03576_ _03098_ vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12405_ _02491_ _02496_ _02497_ vssd1 vssd1 vccd1 vccd1 _02498_ sky130_fd_sc_hd__or3_1
X_13385_ _03500_ _03501_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__xnor2_1
X_16173_ _04449_ _04471_ _03281_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__o21a_1
X_10597_ _00482_ _00487_ _00688_ _00689_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__a211o_2
XFILLER_0_152_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15124_ _05398_ _05401_ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__xor2_2
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput109 net109 vssd1 vssd1 vccd1 vccd1 o_wb_data[4] sky130_fd_sc_hd__clkbuf_4
X_12336_ _02427_ _02428_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15055_ _05324_ _05325_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__nor2_1
X_12267_ _02357_ _02358_ _02359_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__and3b_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11218_ _01290_ _01309_ _01308_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__o21ai_2
X_14006_ _04008_ _04011_ _04009_ vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__o21ba_1
X_12198_ _02285_ _02286_ _02268_ _02275_ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__o211a_1
Xoutput80 net80 vssd1 vssd1 vccd1 vccd1 leds[8] sky130_fd_sc_hd__buf_2
Xoutput91 net91 vssd1 vssd1 vccd1 vccd1 o_wb_data[17] sky130_fd_sc_hd__clkbuf_4
X_18814_ _09320_ vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__clkbuf_1
X_11149_ _00169_ _09188_ _07591_ _00175_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18745_ _02728_ net63 _09251_ vssd1 vssd1 vccd1 vccd1 _09266_ sky130_fd_sc_hd__mux2_1
X_15957_ _06274_ _06302_ _06303_ vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__o21ba_1
X_14908_ _01504_ _01317_ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nand2_1
X_18676_ net38 _09189_ _09215_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__o21a_1
X_15888_ _06227_ _06228_ _06230_ vssd1 vssd1 vccd1 vccd1 _09373_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_144_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17627_ _08119_ _08120_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__or2_1
X_14839_ _03538_ _04241_ _03918_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__and3_1
X_17558_ _06755_ _07741_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16509_ _06902_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__inv_2
X_17489_ _07968_ _07969_ vssd1 vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09814_ _07210_ _07319_ _07472_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__a21o_2
X_09745_ _06722_ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__buf_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _05975_ vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__buf_4
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10520_ _03892_ _05333_ _05039_ _03881_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10451_ _00388_ _00389_ vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13170_ _03005_ _01248_ vssd1 vssd1 vccd1 vccd1 _03269_ sky130_fd_sc_hd__nand2_1
X_10382_ _08724_ _00309_ _00312_ _00311_ vssd1 vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12121_ _03607_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _02104_ _02103_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__xnor2_1
X_11003_ _07352_ _00459_ _01094_ _01095_ vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__nand4_2
X_16860_ _07245_ _07246_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__nand2_1
X_15811_ _02974_ _06144_ _06147_ vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__a21o_1
X_16791_ _07206_ _07208_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__nand2_1
X_18530_ net26 net25 net23 vssd1 vssd1 vccd1 vccd1 _09099_ sky130_fd_sc_hd__or3b_2
X_15742_ _06071_ _06072_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__and2_1
X_12954_ _01106_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18461_ _06328_ _06411_ _06410_ _06024_ vssd1 vssd1 vccd1 vccd1 _09026_ sky130_fd_sc_hd__a211o_1
X_11905_ _01810_ _01903_ vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__xnor2_4
X_15673_ _05991_ _05996_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__nand2_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _02977_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__clkbuf_4
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _07742_ _07747_ _07884_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__and3_1
X_14624_ _02188_ _00502_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__nand2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11836_ net182 vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__inv_2
X_18392_ _03107_ _07596_ vssd1 vssd1 vccd1 vccd1 _08952_ sky130_fd_sc_hd__nand2_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _06371_ _06545_ _07811_ _03311_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__a22o_1
X_14555_ _04614_ _04616_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__nor2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11767_ net175 net180 vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__nand2_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _05213_ cla_inst.in1\[28\] vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and2_2
X_10718_ _00805_ _00809_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__xor2_1
X_17274_ _07637_ _07638_ vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__and2_1
X_14486_ _02984_ _01520_ _07112_ _00308_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__and4_1
XFILLER_0_153_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ _01221_ _01693_ _01774_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__nor3_1
XFILLER_0_70_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19013_ clknet_4_3_0_clk _00103_ vssd1 vssd1 vccd1 vccd1 op_code\[2\] sky130_fd_sc_hd__dfxtp_4
X_16225_ _03161_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__a21o_1
X_13437_ _02976_ _03038_ _03534_ _03558_ _03121_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__o32a_1
XFILLER_0_130_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10649_ _00739_ _00740_ _00529_ _00699_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a211oi_2
Xrebuffer2 _00662_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16156_ sel_op\[3\] _03281_ sel_op\[2\] vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13368_ _03480_ _03481_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__nand2_1
X_15107_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__and2_1
X_12319_ _02410_ _02405_ _02409_ vssd1 vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__and3_1
X_16087_ _03044_ _06444_ vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__and2_1
X_13299_ _03393_ _03394_ _03405_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__or3_2
X_15038_ _04246_ _04249_ _04247_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16989_ _07409_ _07424_ vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09530_ ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _04395_ sky130_fd_sc_hd__buf_6
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18728_ _09245_ _09252_ vssd1 vssd1 vccd1 vccd1 _09253_ sky130_fd_sc_hd__and2_1
X_09461_ _03596_ _03476_ _03618_ _03629_ vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18659_ _09202_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__buf_1
XFILLER_0_94_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09728_ _04973_ _06191_ _06526_ _06537_ vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__a211oi_2
X_09659_ _05551_ _05791_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__xnor2_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12670_ _02733_ _02738_ _02737_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__a21o_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11621_ _01192_ _01712_ _01711_ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14340_ _04350_ _04422_ _04544_ _04545_ vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a211oi_2
X_11552_ _06971_ _04580_ _01643_ _01644_ vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nand4_2
XFILLER_0_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ _00589_ _00595_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__or2_2
X_14271_ _04299_ net127 _04468_ _04469_ vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__o211ai_4
X_11483_ _05736_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16010_ _00644_ _00248_ vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__or2_1
X_10434_ _00507_ _00508_ _00526_ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__o21a_1
X_13222_ _00148_ _09350_ _00212_ _00206_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__and4_1
XFILLER_0_150_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10365_ _00456_ _00457_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__and2b_1
X_13153_ _05453_ _00645_ _07156_ _06732_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__nand4_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _02195_ _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__nand2_1
X_13084_ _02563_ _03175_ _03022_ vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__o21ai_1
X_17961_ _08482_ _08483_ vssd1 vssd1 vccd1 vccd1 _08484_ sky130_fd_sc_hd__nand2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _00387_ _00388_ cla_inst.in2\[25\] _00172_ vssd1 vssd1 vccd1 vccd1 _00389_
+ sky130_fd_sc_hd__and4bb_1
X_12035_ _01106_ _00515_ _02045_ _02127_ vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__or4_4
X_16912_ _07339_ _07340_ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__xnor2_1
X_17892_ _08314_ _08347_ _08408_ vssd1 vssd1 vccd1 vccd1 _08410_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16843_ _02979_ _06642_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16774_ _07149_ _07151_ vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__and2_1
X_13986_ _04155_ _04157_ _04151_ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__o21ai_1
X_18513_ _06248_ _06414_ _09076_ vssd1 vssd1 vccd1 vccd1 _09082_ sky130_fd_sc_hd__o21bai_1
X_15725_ _05917_ _06054_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ _03028_ _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18444_ _08912_ _08965_ vssd1 vssd1 vccd1 vccd1 _09008_ sky130_fd_sc_hd__nor2_1
X_15656_ _05973_ _05978_ _05979_ vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _02949_ _02955_ _02954_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a21bo_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _03377_ cla_inst.in1\[27\] _07102_ _03356_ vssd1 vssd1 vccd1 vccd1 _04837_
+ sky130_fd_sc_hd__a22o_1
X_18375_ _08932_ _08933_ vssd1 vssd1 vccd1 vccd1 _08934_ sky130_fd_sc_hd__xnor2_4
X_11819_ _06460_ _00147_ _01911_ _01909_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__a31o_1
X_15587_ _05815_ _05817_ _05903_ _05904_ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__a211oi_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _02884_ _02886_ vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__or2_2
X_17326_ _07669_ vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__inv_2
X_14538_ _04760_ _04761_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17257_ _07710_ _07716_ vssd1 vssd1 vccd1 vccd1 _07717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14469_ net177 _04684_ _04685_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__o21ai_1
X_16208_ _03281_ _06575_ _06520_ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17188_ _07620_ _07641_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16139_ _06499_ _06500_ _03152_ vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09513_ _03684_ _03640_ _03585_ vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__a21o_1
XFILLER_0_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ cla_inst.in2\[18\] vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__buf_6
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10150_ _00234_ _00242_ vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__xnor2_1
X_10081_ cla_inst.in2\[23\] vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__buf_2
X_13840_ _03997_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__nor2_1
X_13771_ _03085_ _03088_ _03050_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _01051_ _01052_ _01039_ _01050_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15510_ _05819_ _05820_ vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12722_ _02759_ _02790_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16490_ _06877_ _06881_ vssd1 vssd1 vccd1 vccd1 _06882_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15441_ _05654_ _05657_ _05655_ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__o21ba_1
X_12653_ _02710_ _02745_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__or2_1
X_11604_ _00845_ _01695_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__a21oi_2
X_18160_ _06366_ _07592_ _07650_ _07596_ vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__a22o_1
X_15372_ _05651_ _05670_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ ApproximateM_inst.lob_16.lob2.genblk1\[2\].genblk1.mux.sel _01031_ vssd1
+ vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__and2_2
XFILLER_0_26_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17111_ _07345_ _07349_ _07447_ _07448_ _07556_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__o311a_4
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14323_ _04525_ _04527_ vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__nand2_1
X_11535_ _01212_ _01211_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__and2b_1
X_18091_ _07318_ _07706_ vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__nor2_2
XFILLER_0_151_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17042_ _07285_ _07295_ _07405_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__and3_1
X_14254_ _04450_ _04451_ _04558_ _00502_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_151_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11466_ _01557_ _01558_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__xor2_1
XFILLER_0_34_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ _01745_ _00716_ _03304_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10417_ _07788_ _00509_ _07570_ cla_inst.in2\[31\] vssd1 vssd1 vccd1 vccd1 _00510_
+ sky130_fd_sc_hd__a22oi_1
X_14185_ _04355_ _04356_ _04375_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nand3_1
X_11397_ _01468_ _01488_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__nand3_2
XFILLER_0_110_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _03227_ _03231_ _03232_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__and3_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _03892_ _05028_ _00439_ _03881_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__a22o_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18993_ clknet_4_6_0_clk _09359_ vssd1 vssd1 vccd1 vccd1 salida\[46\] sky130_fd_sc_hd__dfxtp_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _00370_ _00371_ _09152_ _09338_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__a211o_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _03090_ _03151_ _03158_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21ai_2
X_17944_ _08464_ _08465_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__and2_1
X_12018_ _07363_ _04045_ _02109_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__a31o_1
X_17875_ _08389_ _08390_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16826_ _07191_ _07192_ _07247_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__nor3_1
X_16757_ _07172_ _06354_ _06355_ vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__nand3_1
X_13969_ _04128_ _04129_ _04138_ vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15708_ _03015_ _03067_ _05960_ _05959_ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__a31o_1
X_16688_ _07096_ _07097_ _06836_ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15639_ _05959_ _03067_ _03015_ _05960_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__and4b_1
X_18427_ _06408_ _06449_ _08989_ vssd1 vssd1 vccd1 vccd1 _08990_ sky130_fd_sc_hd__o21ai_1
X_18358_ _08862_ _08894_ _08914_ vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_84_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_22 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17309_ _07773_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18289_ _08736_ _08739_ _08809_ vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09240_ _09326_ vssd1 vssd1 vccd1 vccd1 _09333_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09427_ sel_op\[3\] _03206_ _03260_ _03239_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _01394_ _01395_ _01412_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11251_ _00169_ _00130_ _01342_ _01343_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _04504_ _00294_ _08049_ _05377_ vssd1 vssd1 vccd1 vccd1 _00295_ sky130_fd_sc_hd__and4_1
X_11182_ _00964_ _00963_ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__or2b_1
XFILLER_0_101_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10133_ _00215_ _00225_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__xnor2_1
X_15990_ _06335_ _06336_ _06337_ vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__a21bo_1
X_10064_ _08202_ _00143_ _00156_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__o21a_1
X_14941_ _04951_ _05200_ _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a21boi_1
X_17660_ _08045_ _08046_ vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__nand2_1
X_14872_ _00678_ _06471_ _08452_ _00679_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__a22o_1
X_16611_ _02828_ _07012_ _03930_ _07013_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__o211a_1
X_13823_ _03963_ _03964_ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__a21o_1
X_17591_ _07954_ _07964_ _08080_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__a21o_1
X_16542_ _06653_ _06937_ _06886_ vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__nor3_1
X_13754_ _03043_ _03046_ _03090_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__mux2_1
X_10966_ _00987_ _00986_ vssd1 vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12705_ _02795_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__and2b_1
X_16473_ _06833_ _06835_ _06864_ vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__o21a_1
X_13685_ _03828_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__nand2_1
X_10897_ _00985_ _00988_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__xor2_1
X_18212_ _04900_ _06446_ vssd1 vssd1 vccd1 vccd1 _08758_ sky130_fd_sc_hd__nor2_1
X_15424_ _05720_ _05727_ vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12636_ _08865_ _01746_ _01357_ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ _08682_ _06396_ _06397_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__and3_1
X_15355_ _05582_ _05581_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ _02613_ _02653_ _02643_ _02652_ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14306_ _04507_ _04508_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11518_ _01552_ _01554_ _01553_ vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__a21bo_1
X_18074_ _04647_ _08428_ _02998_ vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__or3b_1
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15286_ _02993_ _02996_ _09059_ _00322_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12498_ _02580_ _02581_ _02574_ vssd1 vssd1 vccd1 vccd1 _02591_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17025_ _07462_ _07463_ _07464_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__a21o_1
X_14237_ _02986_ _00309_ _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__a22oi_4
X_11449_ _04427_ _03607_ _00217_ _04504_ vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__a22o_1
X_14168_ _04196_ _04204_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__and2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _03210_ _03211_ _03212_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a21o_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _04276_ _04281_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__xnor2_1
X_18976_ clknet_4_7_0_clk _09407_ vssd1 vssd1 vccd1 vccd1 salida\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _08320_ _08412_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__nor2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17858_ _08370_ _08371_ vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ _07193_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__or2_1
X_17789_ _08179_ _08172_ vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09976_ _09172_ _07559_ _07602_ _09166_ vssd1 vssd1 vccd1 vccd1 _09205_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10820_ _03454_ _00909_ _00910_ _00911_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _00836_ _00841_ _00843_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13470_ _03574_ _05039_ _03376_ _03378_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__and4_1
XFILLER_0_94_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ _00771_ _00773_ _03454_ _00774_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_137_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12421_ _02446_ _02447_ _02417_ vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15140_ _04259_ _04262_ _03081_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__mux2_1
X_12352_ _02433_ _02441_ _02443_ _02444_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ _00863_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__inv_2
X_15071_ _05330_ _05341_ vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__or2_1
X_12283_ _02369_ _02372_ _02374_ _02375_ vssd1 vssd1 vccd1 vccd1 _02376_ sky130_fd_sc_hd__or4_4
X_14022_ _00125_ _03750_ _04864_ _00151_ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11234_ _01324_ _01326_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18830_ net35 _03239_ _09331_ vssd1 vssd1 vccd1 vccd1 _09332_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ _01254_ _01257_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__xnor2_1
X_10116_ _00204_ _00207_ _00208_ vssd1 vssd1 vccd1 vccd1 _00209_ sky130_fd_sc_hd__and3_1
X_11096_ _06711_ _04591_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__nand2_2
X_18761_ _09278_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__clkbuf_1
X_15973_ _06282_ _06308_ vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__nand2_1
X_17712_ _08211_ _08212_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__xnor2_1
X_14924_ _05139_ _05183_ vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__xnor2_1
X_10047_ _00123_ _00138_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18692_ _09225_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 net254 sky130_fd_sc_hd__buf_1
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14855_ _05107_ _04972_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nor2_2
X_17643_ _03693_ _06441_ _03111_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__a21oi_1
X_13806_ _03949_ _03950_ _03960_ vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or3_4
XFILLER_0_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17574_ _08043_ _08044_ _08062_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__o21ba_1
X_14786_ _05030_ _05032_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__xnor2_1
X_11998_ _05213_ _00171_ _02012_ _02013_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__o2bb2a_1
X_16525_ _06550_ vssd1 vssd1 vccd1 vccd1 _06921_ sky130_fd_sc_hd__clkbuf_4
X_13737_ _03886_ _03722_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__nor2_1
X_10949_ _00951_ _00950_ vssd1 vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_888 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16456_ _06845_ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__inv_2
X_13668_ _03622_ _03752_ _03809_ net189 vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15407_ _05708_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_ sky130_fd_sc_hd__or2b_1
X_12619_ _02691_ _02711_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16387_ _06769_ _06770_ vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13599_ _03733_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__xor2_1
X_18126_ _08663_ _08570_ _08568_ vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__o21ai_1
X_15338_ _02991_ _09351_ _07123_ _00318_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__nand4_2
XFILLER_0_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _08418_ _08587_ _08588_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__o21a_1
X_15269_ _09351_ _00318_ _05758_ _03322_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17008_ _07443_ _07444_ _07381_ _07336_ vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__o211a_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _07613_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__buf_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _06895_ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__buf_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18959_ clknet_4_6_0_clk _09389_ vssd1 vssd1 vccd1 vccd1 salida\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _05943_ _06138_ _05812_ _05823_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a211o_1
Xrebuffer12 _01845_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_1
Xrebuffer23 _00336_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__buf_1
Xrebuffer34 _06076_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer45 ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel vssd1 vssd1
+ vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer56 net218 vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer67 _05311_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer78 _03376_ vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_1
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer89 _03759_ vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_138_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _08224_ vssd1 vssd1 vccd1 vccd1 _09059_ sky130_fd_sc_hd__buf_4
X_12970_ _03051_ _03059_ _03062_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__mux2_1
X_11921_ _02012_ _02013_ ApproximateM_inst.lob_16.lob2.genblk1\[8\].genblk1.mux.sel
+ _00217_ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__and4bb_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _04871_ vssd1 vssd1 vccd1 vccd1 _04873_ sky130_fd_sc_hd__inv_2
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _01944_ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__inv_2
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _00273_ _00892_ _00856_ _00891_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__a211oi_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _04622_ _04796_ _04797_ vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__or3_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _01872_ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ _06685_ _06332_ _06686_ vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__and3_1
X_13522_ _03449_ _03462_ _03460_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__a21o_1
X_10734_ _00801_ _00818_ _00825_ _00826_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17290_ _07750_ _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16241_ _03027_ _03056_ _00121_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__a21o_1
X_13453_ _03176_ _03182_ _03048_ vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10665_ _00756_ _00590_ _00597_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__and3_1
X_12404_ _02421_ _02490_ _02488_ vssd1 vssd1 vccd1 vccd1 _02497_ sky130_fd_sc_hd__o21a_1
X_16172_ _03739_ _03804_ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__or2_1
X_13384_ _00107_ _00247_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ _00676_ _00677_ _00687_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15123_ _05180_ _05291_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a21bo_2
X_12335_ _02355_ _02354_ vssd1 vssd1 vccd1 vccd1 _02428_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ _05312_ _05313_ _05323_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12266_ _05595_ _00180_ _00130_ _06019_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14005_ _04178_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__xnor2_1
X_11217_ _01290_ _01308_ _01309_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__or3_4
Xoutput70 net70 vssd1 vssd1 vccd1 vccd1 leds[0] sky130_fd_sc_hd__buf_2
X_12197_ _02288_ _02203_ _02289_ vssd1 vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput81 net81 vssd1 vssd1 vccd1 vccd1 leds[9] sky130_fd_sc_hd__clkbuf_4
X_18813_ _09298_ _09319_ vssd1 vssd1 vccd1 vccd1 _09320_ sky130_fd_sc_hd__and2_1
Xoutput92 net92 vssd1 vssd1 vccd1 vccd1 o_wb_data[18] sky130_fd_sc_hd__clkbuf_4
X_11148_ _00702_ _00169_ _07559_ _07602_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__and4_1
XFILLER_0_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18744_ _09265_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__clkbuf_1
X_11079_ _04646_ _04373_ _03432_ _00205_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__nand4_2
X_15956_ _06200_ _06246_ vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__nand2_1
X_14907_ _05163_ _05164_ vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nor2_1
X_18675_ _02259_ _09190_ _09191_ vssd1 vssd1 vccd1 vccd1 _09215_ sky130_fd_sc_hd__a21oi_1
X_15887_ _04828_ _05307_ _06229_ _03039_ vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__o22a_1
X_17626_ _08009_ _08042_ _08118_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__nor3_2
XFILLER_0_59_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14838_ _03539_ _05089_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17557_ _07942_ _07949_ vssd1 vssd1 vccd1 vccd1 _08044_ sky130_fd_sc_hd__nor2_1
X_14769_ _04867_ _04968_ _05012_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16508_ _06834_ _06900_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__or2b_1
X_17488_ _07965_ _07967_ vssd1 vssd1 vccd1 vccd1 _07969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16439_ _06825_ _06826_ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18109_ _08636_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09813_ _07330_ _07461_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__xnor2_2
X_09744_ cla_inst.in1\[24\] vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__clkbuf_4
X_09675_ _05964_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__clkbuf_8
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ _00356_ _00364_ _00355_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10381_ _00472_ _00473_ vssd1 vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12120_ _02211_ _02212_ _05671_ _00205_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__and4b_1
XFILLER_0_103_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12051_ _02140_ _02142_ vssd1 vssd1 vccd1 vccd1 _02144_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11002_ _07069_ net232 net221 _07984_ vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__a22o_1
X_15810_ _03536_ _06146_ _03123_ vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__a21o_1
X_16790_ _06762_ _06947_ _07207_ _06655_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__a22o_1
X_15741_ _06006_ _06010_ _06070_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__or3_1
X_12953_ _03024_ _03045_ vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
X_11904_ _01992_ _01994_ vssd1 vssd1 vccd1 vccd1 _01997_ sky130_fd_sc_hd__xnor2_4
X_15672_ _05991_ _05996_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__or2_2
X_18460_ _02938_ _09023_ _09024_ vssd1 vssd1 vccd1 vccd1 _09025_ sky130_fd_sc_hd__a21oi_2
X_12884_ _07091_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__buf_4
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _04714_ _04717_ _04715_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__o21ba_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _07742_ _07747_ _07884_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__a21oi_1
X_11835_ _01926_ _01927_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__nor2_1
X_18391_ _04853_ _08895_ _08896_ _08948_ _08949_ vssd1 vssd1 vccd1 vccd1 _08950_ sky130_fd_sc_hd__a221o_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17342_ _02200_ _06547_ _06550_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__a21o_1
X_14554_ _00115_ _01866_ _04658_ _04656_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__a31o_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11766_ _01845_ _01858_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__or2_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13505_ _05508_ _05366_ _07374_ _07406_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__nand4_2
X_10717_ _00805_ _00809_ vssd1 vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__and2_1
X_17273_ _07731_ _07734_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__or2b_1
X_14485_ _04584_ _04585_ _04595_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__nor3_1
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11697_ _01760_ _01769_ _01236_ _01789_ vssd1 vssd1 vccd1 vccd1 _01790_ sky130_fd_sc_hd__o211a_4
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19012_ clknet_4_9_0_clk _00102_ vssd1 vssd1 vccd1 vccd1 op_code\[1\] sky130_fd_sc_hd__dfxtp_1
X_16224_ _06551_ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__clkbuf_4
X_13436_ _03539_ _03548_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a21oi_1
X_10648_ _00529_ _00699_ _00739_ _00740_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer3 _06548_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_1
XFILLER_0_130_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ _01151_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel _04340_
+ _04362_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__or4_1
X_13367_ _03480_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__or2_1
X_10579_ _00667_ _00670_ _00671_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _01873_ _03149_ _05380_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__a21o_1
X_12318_ _02405_ _02409_ _02410_ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16086_ _04336_ _03041_ _06443_ vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__and3_1
X_13298_ _03393_ _03394_ _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__o21ai_2
X_15037_ _03117_ _03199_ vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__nand2_4
X_12249_ _02339_ _02341_ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16988_ _07415_ _07423_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18727_ _06477_ net35 _09251_ vssd1 vssd1 vccd1 vccd1 _09252_ sky130_fd_sc_hd__mux2_1
X_15939_ _06219_ _06260_ vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__or2_1
X_09460_ _03345_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__buf_4
X_18658_ _09176_ _09201_ vssd1 vssd1 vccd1 vccd1 _09202_ sky130_fd_sc_hd__and2_1
X_17609_ _08099_ _08100_ vssd1 vssd1 vccd1 vccd1 _08101_ sky130_fd_sc_hd__or2_1
X_18589_ salida\[14\] _09141_ _09142_ salida\[46\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09727_ _06373_ _06515_ _06504_ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09658_ _05725_ _05780_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _05028_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__buf_6
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _01192_ _01711_ _01712_ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__nand3_2
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ _07243_ ApproximateM_inst.lob_16.lob1.genblk2.mux_final.sel ApproximateM_inst.lob_16.lob1.genblk1\[14\].genblk1.mux.sel
+ _07221_ vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ _00587_ _00588_ _00427_ _00430_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__a211oi_1
X_14270_ _04461_ _04462_ _04467_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ _08409_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__buf_8
X_13221_ _03321_ _00212_ _00206_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__a22oi_1
X_10433_ _00524_ _00525_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__nand2_2
XFILLER_0_33_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13152_ _00645_ _07156_ _06732_ _05453_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10364_ _00453_ _00455_ _00454_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12103_ _02193_ _02194_ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__nand2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _03025_ _03101_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__and2_1
X_17960_ _08363_ _08450_ _08481_ vssd1 vssd1 vccd1 vccd1 _08483_ sky130_fd_sc_hd__nand3_1
X_10295_ _00109_ _09349_ _00177_ _00146_ vssd1 vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__and4_1
X_12034_ _00715_ vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__clkinv_4
X_16911_ _07231_ _07239_ _07229_ vssd1 vssd1 vccd1 vccd1 _07340_ sky130_fd_sc_hd__o21ai_1
X_17891_ _08405_ _08407_ vssd1 vssd1 vccd1 vccd1 _08408_ sky130_fd_sc_hd__xor2_1
X_16842_ _06358_ _06356_ _06357_ _07264_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__o31a_1
X_13985_ _04151_ _04155_ _04157_ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or3_1
X_16773_ _03094_ _06463_ _07190_ vssd1 vssd1 vccd1 vccd1 _09416_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18512_ _07256_ _09078_ _09079_ vssd1 vssd1 vccd1 vccd1 _09081_ sky130_fd_sc_hd__and3_1
X_15724_ _06052_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__nor2_1
X_12936_ _01357_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18443_ _09004_ _09006_ vssd1 vssd1 vccd1 vccd1 _09007_ sky130_fd_sc_hd__or2_1
X_15655_ _01356_ _00665_ _05974_ _05976_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__a22o_1
X_12867_ _02918_ _02937_ _02936_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__a21oi_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14606_ _01521_ _07112_ _04707_ _04708_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__and4_1
X_11818_ _01909_ _01910_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__nor2_1
X_15586_ _05895_ _05902_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__nor2_1
X_18374_ _02892_ _08878_ vssd1 vssd1 vccd1 vccd1 _08933_ sky130_fd_sc_hd__nand2_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _02172_ _02470_ _02851_ _02882_ _02890_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__o311a_4
XFILLER_0_56_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _00189_ _00191_ _05257_ _05486_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__and4_1
X_17325_ _07790_ _07791_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__and2b_1
X_11749_ _01676_ _01679_ _01680_ _01670_ vssd1 vssd1 vccd1 vccd1 _01842_ sky130_fd_sc_hd__o31a_1
XFILLER_0_154_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14468_ _04683_ _04684_ _04685_ vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__nor3_2
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17256_ _07714_ _07715_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16207_ _04121_ _03717_ _04351_ vssd1 vssd1 vccd1 vccd1 _06575_ sky130_fd_sc_hd__or3_4
X_13419_ _03538_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__clkbuf_4
X_17187_ _07502_ _07640_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__xnor2_1
X_14399_ _04464_ _04465_ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _01108_ _03136_ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16069_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09512_ _03684_ _03585_ _03640_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ _03356_ _03377_ _03410_ _03432_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nand4_1
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ cla_inst.in2\[24\] vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__clkbuf_4
X_13770_ _03538_ _03915_ _03922_ _06765_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__o211a_1
X_10982_ _01072_ _01073_ _01061_ _01068_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__a211o_1
X_12721_ _02804_ _02813_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15440_ _05743_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__xnor2_1
X_12652_ _02742_ _02744_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__and2_1
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ _00515_ _01692_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nor2_4
X_15371_ _05668_ _05669_ vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__or2_1
X_12583_ _01082_ _01081_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14322_ _04512_ _04513_ _04524_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__or3_1
X_17110_ _07345_ _07349_ _07447_ _07448_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__o31a_1
XFILLER_0_135_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11534_ _05736_ _01005_ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nand2_1
X_18090_ _08622_ _08623_ vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17041_ _07481_ vssd1 vssd1 vccd1 vccd1 _09388_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14253_ _04515_ _04438_ _07755_ _07722_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11465_ _01159_ _01508_ vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13204_ _01745_ _00716_ _03304_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10416_ cla_inst.in1\[31\] vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14184_ _04355_ _04356_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__a21o_1
X_11396_ _01466_ _01467_ _01394_ _01413_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13135_ _05017_ _00308_ _03229_ _03230_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__a22o_1
X_10347_ _03881_ _05028_ _00439_ vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ clknet_4_6_0_clk _09358_ vssd1 vssd1 vccd1 vccd1 salida\[45\] sky130_fd_sc_hd__dfxtp_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _03152_ _03157_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__or2_1
X_17943_ _08458_ _08462_ vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__or2_1
X_10278_ _00369_ _00368_ _08984_ _08930_ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__o211ai_2
X_12017_ _01082_ _01081_ _03388_ _00949_ vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__and4_1
X_17874_ _08301_ _08303_ _08299_ vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__a21bo_1
X_16825_ _07245_ _07246_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__xor2_1
Xmax_cap1 _04218_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_1
X_16756_ _02533_ _03094_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__nand2_1
X_13968_ _04128_ _04129_ _04138_ vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__a21oi_1
X_15707_ _05976_ _05978_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
X_12919_ _07668_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__buf_2
X_13899_ _03897_ _03899_ _04063_ vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__a21oi_1
X_16687_ _06990_ _06991_ _06989_ vssd1 vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ _06408_ _06449_ _06425_ vssd1 vssd1 vccd1 vccd1 _08989_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15638_ _03012_ _03142_ _03055_ _03010_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a22o_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _08912_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__and2_1
X_15569_ _05883_ _03142_ _03015_ _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__and4b_1
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17308_ _07641_ _07620_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__or2b_1
XFILLER_0_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18288_ _08835_ _08837_ _08838_ vssd1 vssd1 vccd1 vccd1 _08839_ sky130_fd_sc_hd__o21a_2
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17239_ _00786_ _06367_ _06369_ _07084_ _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__a311o_1
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09992_ _09287_ _09295_ _09318_ vssd1 vssd1 vccd1 vccd1 _09326_ sky130_fd_sc_hd__nand3_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ _03217_ op_code\[2\] op_code\[3\] vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ cla_inst.in2\[23\] _01031_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel
+ cla_inst.in2\[24\] vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10201_ _04416_ vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__buf_6
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11181_ _00967_ _00976_ _00977_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__nor3_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10132_ _00222_ _00224_ vssd1 vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _00144_ _00155_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__xor2_1
X_14940_ _05078_ _05074_ _05075_ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__a21o_1
X_14871_ _03008_ _07515_ _06471_ _04591_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__and4_1
XFILLER_0_98_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16610_ _02829_ _02828_ vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__nand2_1
X_13822_ _03965_ _03978_ vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__xnor2_1
X_17590_ _07950_ _07953_ vssd1 vssd1 vccd1 vccd1 _08080_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13753_ _03738_ _03747_ _03902_ _02969_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__a31o_1
X_16541_ _06756_ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__buf_2
X_10965_ _05213_ _04482_ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__nand2_2
X_12704_ _02772_ _02796_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ _03642_ _03644_ _03827_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__or3_1
X_16472_ _06836_ _06842_ _06860_ _06862_ vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__o211a_1
X_10896_ _00985_ _00988_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__and2_1
X_18211_ _08753_ _08754_ _08755_ vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__o21a_1
X_15423_ _05724_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__xnor2_1
X_12635_ _06084_ vssd1 vssd1 vccd1 vccd1 _02728_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15354_ _04125_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__clkbuf_4
X_18142_ _02997_ _03052_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ _02615_ _02619_ _02621_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14305_ _04494_ _04347_ _04506_ vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__and3_1
X_11517_ _01607_ _01608_ _01609_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__and3_2
X_15285_ _02996_ _09059_ _00322_ _02993_ vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__a22oi_2
X_18073_ _02998_ _06511_ _01136_ vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ _02531_ _02583_ vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__xnor2_2
X_14236_ _01521_ _05715_ _04430_ _04431_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17024_ _07462_ _07463_ _06507_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11448_ _04504_ _00294_ _00205_ _00217_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__nand4_2
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14167_ _04197_ _04203_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__and2b_1
XFILLER_0_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _00865_ _01471_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _03210_ _03211_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__nand3_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _04279_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__xor2_1
X_18975_ clknet_4_5_0_clk _09406_ vssd1 vssd1 vccd1 vccd1 salida\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _08422_ _08426_ _08446_ _06723_ _01692_ vssd1 vssd1 vccd1 vccd1 _09398_ sky130_fd_sc_hd__o32a_1
X_13049_ _01108_ _03140_ _03023_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__o21a_1
X_17857_ _07109_ _07780_ vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__nand2_1
X_16808_ _07205_ _07227_ vssd1 vssd1 vccd1 vccd1 _07228_ sky130_fd_sc_hd__xnor2_1
X_17788_ _08194_ _08195_ _08295_ vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16739_ _06749_ _06969_ _07055_ _07053_ vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18409_ _08968_ _08967_ vssd1 vssd1 vccd1 vccd1 _08970_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09975_ _09166_ _09172_ _09188_ _07591_ vssd1 vssd1 vccd1 vccd1 _09197_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _00842_ _00840_ _00837_ vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__or3b_1
XFILLER_0_137_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _00774_ sky130_fd_sc_hd__buf_4
XFILLER_0_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ _02510_ _02512_ vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12351_ _02376_ _02442_ _02411_ vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _01392_ _01393_ _01290_ _01379_ vssd1 vssd1 vccd1 vccd1 _01395_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ _05330_ _05341_ vssd1 vssd1 vccd1 vccd1 _05342_ sky130_fd_sc_hd__nand2_1
X_12282_ _02260_ _02371_ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _03987_ _03989_ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__nor2_1
X_11233_ _01085_ _01092_ _01325_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11164_ _01255_ _01256_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__nand2_1
X_10115_ _00188_ _00201_ vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__xnor2_1
X_18760_ _09273_ _09277_ vssd1 vssd1 vccd1 vccd1 _09278_ sky130_fd_sc_hd__and2_1
X_11095_ _01056_ _01182_ _01186_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__a21o_1
X_15972_ _06308_ _06310_ vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__nand2_1
X_17711_ _08102_ _08110_ _08101_ vssd1 vssd1 vccd1 vccd1 _08212_ sky130_fd_sc_hd__a21boi_2
X_14923_ _05180_ _05182_ vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nor2_1
X_10046_ _00123_ _00138_ vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__or2_1
X_18691_ _09209_ _09224_ vssd1 vssd1 vccd1 vccd1 _09225_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17642_ _06382_ _06380_ _06381_ _07084_ _08136_ vssd1 vssd1 vccd1 vccd1 _08138_ sky130_fd_sc_hd__a311o_1
Xhold92 net92 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ _02984_ _01520_ _07733_ _08158_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13805_ _03949_ _03950_ _03960_ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__o21ai_2
X_17573_ _08054_ _08061_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__xnor2_1
X_14785_ _04906_ _04914_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a21oi_1
X_11997_ _02088_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16524_ _06547_ vssd1 vssd1 vccd1 vccd1 _06920_ sky130_fd_sc_hd__clkbuf_4
X_13736_ _03434_ _03586_ _03671_ _03672_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o211a_1
X_10948_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _03837_ vssd1
+ vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__nand2_4
XFILLER_0_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16455_ _03098_ _06467_ _06501_ _06844_ vssd1 vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__a31o_1
X_13667_ _03786_ _03787_ _03807_ _03808_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__and4bb_1
X_10879_ _00970_ _00971_ vssd1 vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15406_ _05626_ _05628_ _05707_ vssd1 vssd1 vccd1 vccd1 _05709_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12618_ _02683_ _02684_ _02690_ vssd1 vssd1 vccd1 vccd1 _02711_ sky130_fd_sc_hd__o21ai_1
X_13598_ _03482_ _03483_ _03486_ _03734_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__a31oi_2
X_16386_ _06757_ _06768_ vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18125_ _08490_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15337_ _09351_ _07123_ _00318_ _02991_ vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__a22o_1
X_12549_ _02602_ _02601_ _02598_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18056_ _08410_ _08447_ _08504_ vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__o21ai_1
XANTENNA_1 _00042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15268_ _03322_ _09351_ _00309_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _07381_ _07336_ _07443_ _07444_ vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_1_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14219_ _03034_ _03100_ _03081_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__mux2_1
X_15199_ _05481_ _05482_ vssd1 vssd1 vccd1 vccd1 _05483_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _06548_ _06863_ _06873_ _06884_ vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__and4b_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18958_ clknet_4_6_0_clk _09388_ vssd1 vssd1 vccd1 vccd1 salida\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _07355_ vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__buf_2
X_09691_ _05812_ _05823_ _05943_ _06138_ vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__o211ai_2
X_18889_ clknet_4_9_0_clk _00043_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[7\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer13 _01957_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_1
Xrebuffer24 _02118_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_1
Xrebuffer35 _01769_ vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
Xrebuffer46 ApproximateM_inst.lob_16.lob1.genblk1\[11\].genblk1.mux.sel vssd1 vssd1
+ vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer57 _00980_ vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer68 net233 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer79 net172 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__buf_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _07330_ _07461_ vssd1 vssd1 vccd1 vccd1 _09048_ sky130_fd_sc_hd__nand2_1
X_09889_ _06906_ _06928_ _05181_ _06181_ vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__o211ai_1
X_11920_ _05290_ _00176_ _00145_ _00806_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _01919_ _01941_ _01943_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__a21oi_2
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _00231_ _00857_ _00894_ _00859_ _00888_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__a32o_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _04794_ _04795_ _04775_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11782_ _01742_ _01874_ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__nor2_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _03647_ _03648_ _03408_ _03433_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__o211a_1
X_10733_ _08126_ _08137_ _08256_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _06467_ _06610_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__nand2_1
X_13452_ _03171_ _03174_ _03048_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__mux2_1
X_10664_ _00590_ _00597_ _00756_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__a21oi_1
X_12403_ _02495_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13383_ _03497_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16171_ _03281_ sel_op\[3\] vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__or2b_1
X_10595_ _00676_ _00677_ _00687_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_152_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15122_ _05289_ _05288_ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__or2b_1
X_12334_ _07352_ _00211_ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15053_ _05312_ _05313_ _05323_ vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__a21oi_1
X_12265_ ApproximateM_inst.lob_16.lob2.genblk1\[5\].genblk1.mux.sel _00909_ vssd1
+ vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__and2_2
XFILLER_0_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14004_ _00253_ _06482_ vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__nand2_1
X_11216_ _01288_ _01289_ _00967_ _01274_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_121_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12196_ _02144_ _02145_ vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__or2_1
Xoutput71 net71 vssd1 vssd1 vccd1 vccd1 leds[10] sky130_fd_sc_hd__buf_2
Xoutput82 net82 vssd1 vssd1 vccd1 vccd1 o_wb_ack sky130_fd_sc_hd__clkbuf_4
X_18812_ _02992_ net54 _09301_ vssd1 vssd1 vccd1 vccd1 _09319_ sky130_fd_sc_hd__mux2_1
X_11147_ _01239_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__inv_2
Xoutput93 net93 vssd1 vssd1 vccd1 vccd1 o_wb_data[19] sky130_fd_sc_hd__clkbuf_4
X_18743_ _09245_ _09264_ vssd1 vssd1 vccd1 vccd1 _09265_ sky130_fd_sc_hd__and2_1
X_11078_ _01167_ _01170_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__xor2_2
X_15955_ _06248_ vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__inv_2
X_14906_ _00190_ _05986_ _05162_ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__and3_1
X_10029_ _07853_ _00119_ _00121_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__nand3_4
X_18674_ _09214_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15886_ _04826_ _04827_ _03537_ vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__mux2_1
X_17625_ _08009_ _08042_ _08118_ vssd1 vssd1 vccd1 vccd1 _08119_ sky130_fd_sc_hd__o21a_1
X_14837_ _05087_ _05088_ _03916_ vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ _07938_ _07941_ vssd1 vssd1 vccd1 vccd1 _08043_ sky130_fd_sc_hd__nor2_1
X_14768_ _04999_ _05000_ _05011_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16507_ _06866_ _06900_ vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13719_ _03865_ _03866_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__nor2_1
X_17487_ _07965_ _07967_ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__or2_1
X_14699_ _04936_ _04937_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16438_ _06749_ _06763_ vssd1 vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__nand2_2
XFILLER_0_144_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16369_ _04121_ _03281_ vssd1 vssd1 vccd1 vccd1 _06751_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18108_ _08641_ _08643_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18039_ _08477_ _08566_ _08567_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09812_ _07341_ _07450_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__xor2_2
XFILLER_0_10_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09743_ _05671_ vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__buf_4
X_09674_ _05606_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__buf_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10380_ _05235_ _07134_ _00470_ _00471_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ _02140_ _02142_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__and2b_1
X_11001_ _07036_ _07069_ _08049_ net221 vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__nand4_2
X_15740_ _06006_ _06010_ _06070_ vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__o21ai_2
X_12952_ _03027_ _03044_ _01696_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a21o_1
X_11903_ _01810_ _01903_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15671_ _05994_ _05995_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand2_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _02975_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__buf_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _07738_ _07764_ _07762_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__a21oi_1
X_14622_ _04849_ _04850_ _04851_ vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _01920_ _01921_ _01925_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__o21ba_1
X_18390_ _08896_ _08947_ vssd1 vssd1 vccd1 vccd1 _08949_ sky130_fd_sc_hd__nor2_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _06440_ _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__nor2_1
X_14553_ _04653_ _04661_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11765_ _01848_ _01856_ _01857_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a21oi_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13504_ _05301_ cla_inst.in1\[27\] _07004_ _05279_ vssd1 vssd1 vccd1 vccd1 _03632_
+ sky130_fd_sc_hd__a22o_1
X_10716_ _08724_ _06482_ _00807_ _00808_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17272_ _07703_ _07704_ _07732_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__or3b_1
X_14484_ _04586_ _04594_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__nand2_1
X_11696_ _01233_ _01234_ _01235_ _01204_ vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19011_ clknet_4_9_0_clk _00101_ vssd1 vssd1 vccd1 vccd1 op_code\[0\] sky130_fd_sc_hd__dfxtp_2
X_16223_ _06592_ vssd1 vssd1 vccd1 vccd1 _06593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ _00737_ _00738_ _00718_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_64_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13435_ _03538_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer4 net166 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_1
X_13366_ _00877_ _03311_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__nand2_1
X_16154_ _05213_ _03004_ _03019_ _06517_ vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__or4_1
X_10578_ _06982_ _00509_ _00668_ _00669_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__a22o_1
X_15105_ _00591_ _03149_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__nand3_1
XFILLER_0_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12317_ _02339_ _02341_ vssd1 vssd1 vccd1 vccd1 _02410_ sky130_fd_sc_hd__xnor2_1
X_13297_ _03395_ _03404_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__xnor2_2
X_16085_ _01678_ _06442_ vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12248_ _02340_ _02335_ vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15036_ _04243_ _04245_ _04247_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__mux2_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12179_ _01113_ _02045_ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__nor2_2
X_16987_ _07421_ _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__xnor2_1
X_18726_ _09250_ vssd1 vssd1 vccd1 vccd1 _09251_ sky130_fd_sc_hd__clkbuf_4
X_15938_ _06282_ _06283_ vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__or2_2
X_18657_ net63 _03169_ _09193_ vssd1 vssd1 vccd1 vccd1 _09201_ sky130_fd_sc_hd__mux2_1
X_15869_ _06095_ _06165_ _06167_ vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__o21a_1
X_17608_ _07969_ _07994_ _07968_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18588_ net299 _09140_ _09149_ _09144_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17539_ _08023_ _08024_ vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09726_ _06373_ _06504_ _06515_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09657_ _05747_ _05758_ _05769_ _05660_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__a22oi_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ cla_inst.in1\[17\] vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__buf_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11550_ _07984_ _07973_ _04449_ _04471_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nand4_2
XFILLER_0_107_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10501_ _00592_ _00593_ _00413_ _00412_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11481_ _01568_ _01569_ _01572_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_107_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13220_ _00151_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10432_ _00519_ _00523_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__or2_1
X_13151_ _08724_ _07123_ _00647_ _00648_ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__and4_1
XFILLER_0_20_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10363_ _00453_ _00454_ _00455_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__and3_1
X_12102_ _02193_ _02194_ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13082_ _02607_ _03173_ _03040_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__o21ai_1
X_10294_ _00125_ _00178_ _00181_ _00151_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a22oi_1
X_12033_ _07711_ _02124_ _02125_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__and3_2
X_16910_ _07331_ _07338_ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__xor2_1
X_17890_ _08296_ _08310_ _08406_ vssd1 vssd1 vccd1 vccd1 _08407_ sky130_fd_sc_hd__a21bo_1
X_16841_ _06598_ _07263_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__nor2_1
X_16772_ _07160_ _07161_ _07164_ _07188_ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__o211a_1
X_13984_ _03014_ _00399_ _04153_ _04156_ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__a22oi_1
X_18511_ _09075_ _09056_ _09077_ vssd1 vssd1 vccd1 vccd1 _09079_ sky130_fd_sc_hd__o21ai_1
X_15723_ _06048_ _06050_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ _02505_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18442_ _08955_ _08958_ _09003_ vssd1 vssd1 vccd1 vccd1 _09006_ sky130_fd_sc_hd__and3_1
X_15654_ _05977_ vssd1 vssd1 vccd1 vccd1 _05978_ sky130_fd_sc_hd__inv_2
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _01502_ _02891_ _02894_ _02940_ _02958_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__o311ai_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _02984_ _01520_ _07015_ _07962_ vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__and4_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11817_ _04362_ _00196_ _00871_ _04340_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a22oi_1
X_18373_ _01502_ _02888_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__nor2_2
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15585_ _05895_ _05902_ vssd1 vssd1 vccd1 vccd1 _05903_ sky130_fd_sc_hd__and2_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__inv_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17324_ _07701_ _07702_ _07789_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nand3_1
X_14536_ _00191_ _00460_ _05486_ _00189_ vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_56_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11748_ _01836_ _01839_ _01828_ _01840_ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_153_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17255_ _06766_ _07387_ vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__nor2_1
X_14467_ _04508_ _04510_ _04507_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__o21ba_1
X_11679_ _01733_ _01734_ _01736_ vssd1 vssd1 vccd1 vccd1 _01772_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16206_ net212 _03019_ _06517_ vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__or3_1
X_13418_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__clkbuf_4
X_17186_ _07629_ _07639_ vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__xnor2_1
X_14398_ _04461_ _04468_ _04606_ _04607_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a211o_4
XFILLER_0_12_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16137_ _01220_ _03134_ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__or2_1
X_13349_ _03460_ _03461_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16068_ _06423_ vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15019_ _05285_ _05286_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09511_ _04023_ _04176_ vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18709_ _09237_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__buf_1
XFILLER_0_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09442_ _03421_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__clkbuf_8
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09709_ _06267_ _06319_ _06329_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__nand3_2
X_10981_ _01061_ _01068_ _01072_ _01073_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _02810_ _02812_ vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nor2_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12651_ _02735_ _02742_ _02743_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__nand3_1
XFILLER_0_84_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _05856_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__buf_4
X_15370_ _00591_ _05652_ _05667_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__a21oi_1
X_12582_ _02638_ _02636_ _02637_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__nand3_1
XFILLER_0_154_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ _04512_ _04513_ _04524_ vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11533_ _01622_ _01623_ _01624_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__a21o_1
X_17040_ _00593_ _06463_ _07453_ _07480_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14252_ _02188_ _09303_ _00498_ _04515_ vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__a22oi_1
X_11464_ _01160_ _01161_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10415_ _00506_ _00492_ _00493_ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__and3_1
X_13203_ _03302_ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14183_ _04372_ _04374_ vssd1 vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__nand2_1
X_11395_ _01486_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__xor2_1
X_13134_ _04558_ _05715_ _03229_ _03230_ vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__nand4_1
X_10346_ cla_inst.in1\[16\] vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_4
X_18991_ clknet_4_6_0_clk _09357_ vssd1 vssd1 vccd1 vccd1 salida\[44\] sky130_fd_sc_hd__dfxtp_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _07766_ _03156_ _03024_ vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__o21ai_1
X_17942_ _08458_ _08462_ vssd1 vssd1 vccd1 vccd1 _08464_ sky130_fd_sc_hd__nand2_1
X_10277_ _08930_ _08984_ _00368_ _00369_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__a211o_2
X_12016_ _01081_ _03388_ _00949_ _01082_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__a22o_1
X_17873_ _08386_ _08388_ vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__nor2_1
X_16824_ _07140_ _07141_ _07146_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap2 _03204_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_1
X_16755_ _07168_ _07170_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__xor2_1
X_13967_ _04136_ _04137_ vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ _06032_ _06033_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__and2_1
X_12918_ _03010_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__clkbuf_4
X_16686_ _07094_ _07095_ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__and2b_1
X_13898_ _03896_ _03895_ vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18425_ _06024_ _06409_ _06407_ _06330_ vssd1 vssd1 vccd1 vccd1 _08988_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15637_ _03010_ _03012_ _03142_ _03055_ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__and4_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _00592_ _00167_ _00228_ _00227_ vssd1 vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18356_ _08856_ _08859_ _08911_ vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__or3_1
X_15568_ _07668_ _00119_ _01317_ _03009_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__a22o_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ _07502_ _07640_ vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__and2_1
X_14519_ _04598_ _04701_ _04739_ _04740_ vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__a211o_4
X_18287_ _08835_ _08837_ _06836_ vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__a21oi_1
X_15499_ _05685_ _05732_ vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17238_ _00786_ _06369_ _06367_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17169_ _00716_ _06889_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__nand2_4
XFILLER_0_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09991_ _07711_ _09311_ _09263_ vssd1 vssd1 vccd1 vccd1 _09318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09425_ _03184_ _03206_ _03228_ _03239_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10200_ _04558_ _05257_ vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _01238_ _01271_ _01272_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__nor3_1
XFILLER_0_101_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10131_ _00190_ _00192_ _00223_ _00193_ _00186_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a41o_1
XFILLER_0_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10062_ _00153_ _00154_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__and2_1
X_14870_ _03006_ _03107_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__nand2_1
X_13821_ _03967_ _03977_ vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16540_ _06749_ _06762_ _06893_ vssd1 vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__and3_1
X_13752_ _03738_ _03747_ _03902_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ _01054_ _01056_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12703_ _02769_ _02771_ vssd1 vssd1 vccd1 vccd1 _02796_ sky130_fd_sc_hd__nor2_1
X_16471_ _02826_ _02968_ _06861_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__or3_1
X_13683_ _03642_ _03644_ _03827_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10895_ _05224_ _08409_ _00986_ _00987_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__a31o_1
X_18210_ _08753_ _08754_ _06836_ vssd1 vssd1 vccd1 vccd1 _08755_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15422_ _00115_ _09059_ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12634_ _02712_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18141_ _08675_ _08679_ _08677_ vssd1 vssd1 vccd1 vccd1 _08680_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_143_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15353_ _05646_ _05650_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12565_ _02655_ _02657_ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14304_ _04494_ _04347_ _04506_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11516_ _01556_ _01559_ _01519_ _01557_ vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18072_ _06543_ _08599_ _08600_ _08604_ vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__a31o_1
X_15284_ _03000_ _00339_ _05489_ vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12496_ _02587_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__or2_2
XFILLER_0_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17023_ _07357_ _07360_ _07356_ vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__a21boi_2
X_14235_ _03651_ _03662_ _06722_ _06689_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__nand4_2
XFILLER_0_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11447_ _01526_ _01539_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__nand2_2
XFILLER_0_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14166_ _04195_ _04206_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__nand2_1
X_11378_ _00863_ _00864_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__and2_1
X_13117_ _00604_ _00606_ _00605_ vssd1 vssd1 vccd1 vccd1 _03212_ sky130_fd_sc_hd__a21bo_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _00418_ _00419_ _00420_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a21o_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _02059_ _07025_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__nand2_1
X_18974_ clknet_4_4_0_clk _09405_ vssd1 vssd1 vccd1 vccd1 salida\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _07256_ _08432_ _08433_ _08445_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__a31o_1
X_13048_ _02505_ _06776_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__nor2_1
X_17856_ _08368_ _08369_ vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__nor2_1
X_16807_ _07224_ _07226_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__xor2_1
X_17787_ _08188_ _08196_ vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__or2b_1
X_14999_ _00191_ _00318_ _05758_ _00189_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16738_ _07149_ _07151_ vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16669_ _03790_ _06593_ _06594_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18408_ _08967_ _08968_ vssd1 vssd1 vccd1 vccd1 _08969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18339_ _08864_ _08866_ vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09974_ _09179_ vssd1 vssd1 vccd1 vccd1 _09188_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10680_ net169 _04220_ _00772_ net228 vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_137_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _02376_ _02411_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__and3_2
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11301_ _01290_ _01379_ _01392_ _01393_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__o211a_2
XFILLER_0_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12281_ _00846_ _00399_ _02373_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14020_ _09353_ _00716_ _04033_ _04032_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a31o_1
X_11232_ _01086_ _01091_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11163_ _00174_ _07548_ _07581_ cla_inst.in2\[24\] vssd1 vssd1 vccd1 vccd1 _01256_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10114_ _00206_ vssd1 vssd1 vccd1 vccd1 _00207_ sky130_fd_sc_hd__buf_4
X_11094_ _01056_ _01182_ _01186_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__nand3_4
X_15971_ _06313_ _06315_ _06317_ _03124_ _06318_ vssd1 vssd1 vccd1 vccd1 _09376_ sky130_fd_sc_hd__a221o_1
X_17710_ _08208_ _08210_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__xor2_1
X_14922_ _05140_ _05056_ _05179_ vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__and3_1
X_10045_ _00124_ _00137_ vssd1 vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__xor2_1
X_18690_ net45 _03041_ _09193_ vssd1 vssd1 vccd1 vccd1 _09224_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold82 ApproximateM_inst.lob_16.lob1.mux.sel vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _06382_ _06381_ _06380_ vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__a21oi_1
X_14853_ _05103_ _05105_ vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__or2_2
Xhold93 _00022_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ _03951_ _03959_ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__xnor2_1
X_17572_ _08058_ _08059_ vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__nor2_1
X_14784_ _04913_ _04907_ vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11996_ _02017_ _02020_ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__xnor2_1
X_16523_ _02974_ _06915_ _06918_ _06645_ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__a211o_1
X_13735_ _03834_ _03835_ _03882_ _03883_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10947_ _04984_ _00206_ _01025_ _01024_ vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__a31o_2
XFILLER_0_133_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16454_ _03060_ _06492_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__nor2_1
X_13666_ _03786_ _03787_ _03807_ _03808_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10878_ _04438_ _04864_ _04143_ _04646_ vssd1 vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_128_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15405_ _05626_ _05628_ _05707_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__and3_1
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12617_ _02694_ _02709_ vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__xor2_1
X_16385_ _06757_ _06768_ vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13597_ _00592_ _03108_ _03488_ vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__and3_1
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _08660_ _08661_ vssd1 vssd1 vccd1 vccd1 _08662_ sky130_fd_sc_hd__or2_1
X_15336_ _05449_ _01139_ _05539_ _05538_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12548_ _02597_ _02639_ _02640_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__and3_1
X_18055_ _08413_ _08505_ vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__or2b_1
X_15267_ _09353_ _00119_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__nand2_2
XANTENNA_2 _00100_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _02566_ _02542_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__and2b_1
XFILLER_0_112_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17006_ _07382_ _07383_ _07442_ vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__and3_1
X_14218_ _03125_ _04257_ _04265_ _03199_ _04412_ vssd1 vssd1 vccd1 vccd1 _09383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15198_ _00190_ _00192_ _07025_ _08876_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__and4_1
XFILLER_0_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14149_ _01873_ _04336_ vssd1 vssd1 vccd1 vccd1 _04337_ sky130_fd_sc_hd__nand2_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ clknet_4_6_0_clk _09387_ vssd1 vssd1 vccd1 vccd1 salida\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _03368_ _06511_ _01692_ vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__a21o_1
X_09690_ _05943_ _05954_ _06127_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__nand3_4
X_18888_ clknet_4_12_0_clk _00042_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[6\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
Xrebuffer14 _04683_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_1
X_17839_ _07751_ _07489_ _07596_ _07039_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__a22o_1
Xrebuffer25 _04599_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_1
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer36 _01859_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__buf_1
Xrebuffer47 _01803_ vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__clkbuf_1
Xrebuffer58 _05377_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer69 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09957_ _07341_ _07450_ vssd1 vssd1 vccd1 vccd1 _09037_ sky130_fd_sc_hd__nand2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _08126_ _08267_ _07919_ _07930_ vssd1 vssd1 vccd1 vccd1 _08289_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_99_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _01884_ _01942_ vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__nand2_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _00162_ _00230_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__or2_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _01873_ _01357_ _01680_ vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13520_ _03408_ _03433_ _03647_ _03648_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__a211oi_4
X_10732_ _08126_ _08137_ _08256_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13451_ _03569_ _03572_ _03547_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__mux2_1
X_10663_ _00754_ _00755_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12402_ _02492_ _02493_ _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16170_ _00181_ _06532_ _06533_ _06534_ _03313_ vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__o32a_1
XFILLER_0_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13382_ _00112_ _03321_ _00165_ _00212_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__and4_1
X_10594_ _00684_ _00686_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__xor2_2
X_15121_ _05396_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12333_ _02423_ _02425_ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15052_ _05320_ _05321_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12264_ _06019_ _08039_ _00180_ _00130_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14003_ _04175_ _04177_ vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__nor2_1
X_11215_ _01306_ _01307_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__nand2_1
X_12195_ _02144_ _02145_ vssd1 vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput72 net72 vssd1 vssd1 vccd1 vccd1 leds[11] sky130_fd_sc_hd__buf_2
X_18811_ _09317_ vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__clkbuf_1
X_11146_ _00253_ cla_inst.in2\[21\] _07570_ _07613_ vssd1 vssd1 vccd1 vccd1 _01239_
+ sky130_fd_sc_hd__and4_1
Xoutput83 net83 vssd1 vssd1 vccd1 vccd1 o_wb_data[0] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 vssd1 vssd1 vccd1 vccd1 o_wb_data[1] sky130_fd_sc_hd__clkbuf_4
X_11077_ _01168_ _01169_ vssd1 vssd1 vccd1 vccd1 _01170_ sky130_fd_sc_hd__xnor2_2
X_18742_ _03036_ net62 _09251_ vssd1 vssd1 vccd1 vccd1 _09264_ sky130_fd_sc_hd__mux2_1
X_15954_ _06300_ vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__inv_2
X_14905_ _00190_ _05986_ _05162_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__a21oi_1
X_10028_ _00120_ _08158_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__and2_4
X_18673_ _09209_ _09213_ vssd1 vssd1 vccd1 vccd1 _09214_ sky130_fd_sc_hd__and2_1
X_15885_ _06192_ _06226_ _02969_ vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__a21o_1
X_17624_ _08116_ _08117_ vssd1 vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__nor2_1
X_14836_ _03051_ _03114_ _02981_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17555_ _08011_ _08012_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14767_ _04999_ _05000_ _05011_ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _01973_ _01974_ _01975_ _01944_ vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__o22a_1
X_16506_ _06826_ _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__xor2_2
X_13718_ cla_inst.in2\[27\] cla_inst.in2\[26\] _03837_ _03410_ vssd1 vssd1 vccd1 vccd1
+ _03866_ sky130_fd_sc_hd__and4_1
XFILLER_0_85_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17486_ _07840_ _07849_ _07966_ vssd1 vssd1 vccd1 vccd1 _07967_ sky130_fd_sc_hd__a21oi_1
X_14698_ _04807_ _04808_ _04805_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16437_ _06657_ _06749_ _06763_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__a21o_1
X_13649_ _06040_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__buf_4
XFILLER_0_144_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16368_ _06749_ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ _07106_ _07861_ _08642_ _08639_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__o22a_1
X_15319_ _05612_ _05613_ vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16299_ _06513_ _06587_ _06586_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _08477_ _08566_ _08567_ vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ _07395_ _07439_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__xnor2_2
X_09742_ _05649_ _05704_ _06689_ _06029_ vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09673_ _05529_ _05867_ _05932_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a21o_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11000_ _01085_ _01092_ vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ _01223_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11902_ _01992_ _01994_ vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__or2_1
X_15670_ _05920_ _05993_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _02974_ vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__buf_4
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _04849_ _04850_ _04851_ vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__and3_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _01920_ _01921_ _01925_ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__nor3b_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _06368_ _06438_ _03311_ vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__a21oi_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _04654_ _04660_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__and2b_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11764_ _01852_ _01855_ vssd1 vssd1 vccd1 vccd1 _01857_ sky130_fd_sc_hd__and2_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _03418_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__inv_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17271_ _07729_ _07730_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nand2_1
X_10715_ _00806_ _06591_ _04569_ _04449_ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__and4_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14483_ _04587_ _04593_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_153_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11695_ _01748_ _01778_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__and2b_1
X_19010_ clknet_4_1_0_clk _09378_ vssd1 vssd1 vccd1 vccd1 salida\[63\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16222_ _06547_ vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _03551_ _03555_ _02780_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__mux2_1
X_10646_ _00718_ _00737_ _00738_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__or3_2
XFILLER_0_153_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16153_ _03771_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel _03184_
+ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__or3b_2
Xrebuffer5 _06541_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__buf_1
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13365_ _03478_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__xor2_1
X_10577_ _07363_ _00509_ _00668_ _00669_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__nand4_1
XFILLER_0_134_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15104_ _05378_ _05379_ vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__xnor2_1
X_12316_ _02360_ _02406_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16084_ _03111_ _03693_ _06441_ vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__and3_1
X_13296_ _03402_ _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15035_ _05302_ _05303_ _04823_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__o21ai_1
X_12247_ _02208_ _02331_ vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12178_ _02128_ _02258_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ _01137_ _01221_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16986_ _07304_ _07306_ _07301_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__o21ba_1
X_18725_ _09110_ _09115_ _09178_ vssd1 vssd1 vccd1 vccd1 _09250_ sky130_fd_sc_hd__nor3_4
X_15937_ _06242_ _06254_ _06281_ vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__and3_1
X_15868_ _06207_ _06208_ vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__nand2_1
X_18656_ _09200_ vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17607_ _08083_ _08098_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__xnor2_1
X_14819_ _04932_ _04964_ _05067_ _05068_ vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__o211ai_4
X_15799_ _06134_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18587_ salida\[13\] _09141_ _09142_ salida\[45\] _09146_ vssd1 vssd1 vccd1 vccd1
+ _09149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17538_ _03693_ _07355_ _02989_ vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__or3b_1
XFILLER_0_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17469_ _07945_ _07946_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09725_ _06340_ _06351_ _06362_ vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__a21o_1
X_09656_ _05627_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__inv_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05017_ sky130_fd_sc_hd__buf_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10500_ _00399_ vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11480_ _01568_ _01569_ _01572_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__nand3_1
XFILLER_0_135_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10431_ _00519_ _00523_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _00644_ _00645_ _07134_ _00309_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__and4_1
X_10362_ _04690_ _08757_ _00451_ _00452_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__a22o_1
X_12101_ _02098_ _02101_ vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__xnor2_1
X_10293_ _09197_ _09226_ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__nor2_1
X_13081_ _03025_ _03094_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__and2_1
X_12032_ _00514_ _02044_ vssd1 vssd1 vccd1 vccd1 _02125_ sky130_fd_sc_hd__nor2_2
X_16840_ _06358_ _06357_ _06356_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__o21a_1
X_16771_ _06508_ _07171_ _07187_ vssd1 vssd1 vccd1 vccd1 _07188_ sky130_fd_sc_hd__a21oi_1
X_13983_ net218 vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__inv_2
X_15722_ _06048_ _06050_ vssd1 vssd1 vccd1 vccd1 _06052_ sky130_fd_sc_hd__nor2_1
X_18510_ _09075_ _09056_ _09077_ vssd1 vssd1 vccd1 vccd1 _09078_ sky130_fd_sc_hd__or3_1
X_12934_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15653_ _00115_ _00665_ _05974_ _05976_ vssd1 vssd1 vccd1 vccd1 _05977_ sky130_fd_sc_hd__and4_1
X_18441_ _08955_ _08958_ _09003_ vssd1 vssd1 vccd1 vccd1 _09004_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12865_ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__inv_2
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _04723_ _04724_ _04734_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__nor3_2
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _08927_ _08928_ vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__nand2_1
X_11816_ _04493_ _04416_ _00129_ ApproximateM_inst.lob_16.lob1.genblk1\[2\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__and4_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _05900_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__xnor2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12796_ _02887_ _01502_ _02888_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__or3_4
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17323_ _07701_ _07702_ _07789_ vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__a21oi_1
X_14535_ _04754_ _04757_ _04609_ _04699_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__o211ai_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _01820_ _01826_ _01827_ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__nand3_2
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17254_ _07712_ _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__nor2_1
X_14466_ _04681_ _04682_ _04564_ _04565_ vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__o211a_2
XFILLER_0_50_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11678_ _01721_ _01739_ net198 _01770_ vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_126_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16205_ _06084_ _06711_ _06524_ vssd1 vssd1 vccd1 vccd1 _06573_ sky130_fd_sc_hd__or3_1
XFILLER_0_52_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13417_ _03536_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10629_ _00544_ _00551_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__nand2_1
X_17185_ _07637_ _07638_ vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__xor2_1
X_14397_ _04606_ _04607_ _04461_ _04468_ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16136_ _02983_ _06495_ _06497_ _06467_ vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__o211a_1
X_13348_ _03450_ _03451_ _03459_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16067_ _06418_ _06422_ vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__or2_1
X_13279_ _03892_ _06613_ _08049_ _03881_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15018_ _05161_ _05178_ _05158_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16969_ _07288_ _07291_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__a21o_1
X_09510_ _04110_ _04165_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__nor2_2
X_18708_ _09209_ _09236_ vssd1 vssd1 vccd1 vccd1 _09237_ sky130_fd_sc_hd__and2_1
X_09441_ ApproximateM_inst.lob_16.lob1.genblk1\[8\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _03421_ sky130_fd_sc_hd__buf_6
X_18639_ net46 _01746_ _09183_ vssd1 vssd1 vccd1 vccd1 _09186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _06234_ _06245_ _06256_ vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__a21o_1
X_10980_ _01069_ _01070_ _01071_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09639_ ApproximateM_inst.lob_16.lob2.genblk1\[6\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _05584_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12650_ _02740_ _02741_ _02733_ _02739_ vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _01693_ _01673_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__and2b_1
X_12581_ _02597_ _02639_ _02640_ vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__nand3_1
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _04325_ _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11532_ _01622_ _01623_ _01624_ vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nand3_2
XFILLER_0_93_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _02059_ _07025_ _04278_ _04277_ _08876_ vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__a32o_1
X_11463_ _01552_ _01555_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13202_ _01505_ _00399_ _00705_ _00704_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a31o_1
X_10414_ _00492_ _00493_ _00506_ vssd1 vssd1 vccd1 vccd1 _00507_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14182_ _04357_ _04358_ _04371_ vssd1 vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or3_1
X_11394_ _01358_ _01420_ _01434_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ _04646_ _04373_ _05606_ _05617_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__nand4_2
X_10345_ _00435_ _00436_ _00437_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__nand3_1
X_18990_ clknet_4_3_0_clk _09356_ vssd1 vssd1 vccd1 vccd1 salida\[43\] sky130_fd_sc_hd__dfxtp_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _03026_ _03155_ vssd1 vssd1 vccd1 vccd1 _03156_ sky130_fd_sc_hd__and2_1
X_17941_ _08459_ _08461_ vssd1 vssd1 vccd1 vccd1 _08462_ sky130_fd_sc_hd__xnor2_1
X_10276_ _00349_ _00350_ _00367_ vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__and3_1
X_12015_ _02031_ _02039_ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__xnor2_1
X_17872_ _07630_ _07861_ _08385_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__o21a_1
X_16823_ _07240_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__xor2_1
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13966_ _03970_ _03973_ _03971_ vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__o21ba_1
X_16754_ _06990_ _06991_ _07096_ _07169_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__a31o_1
Xmax_cap3 _03884_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__clkbuf_1
X_12917_ _03009_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__buf_2
X_15705_ _03007_ _03055_ _06031_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__a21o_1
X_16685_ _00881_ _06673_ _03790_ vssd1 vssd1 vccd1 vccd1 _07095_ sky130_fd_sc_hd__or3b_1
X_13897_ _04060_ _04061_ vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__xor2_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18424_ _02920_ net115 _08986_ vssd1 vssd1 vccd1 vccd1 _08987_ sky130_fd_sc_hd__a21o_1
X_12848_ _02928_ _02929_ _02931_ vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__and3_1
X_15636_ _03007_ _04900_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__nand2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15567_ _03009_ _07668_ _00119_ _01317_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18355_ _08856_ _08859_ _08911_ vssd1 vssd1 vccd1 vccd1 _08912_ sky130_fd_sc_hd__o21ai_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _02853_ _02865_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _04737_ _04738_ _04702_ _04703_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17306_ _07769_ _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__xnor2_1
X_15498_ _05773_ _05757_ _05759_ vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__nand3_1
X_18286_ _08753_ _08754_ _08815_ _08836_ vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ _04651_ _04652_ _04663_ vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__or3_1
X_17237_ _03198_ _05086_ _07693_ _07695_ vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17168_ _07518_ _07528_ _07525_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16119_ _06470_ _06478_ _03077_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__a21o_1
X_09990_ _09303_ vssd1 vssd1 vccd1 vccd1 _09311_ sky130_fd_sc_hd__buf_4
X_17099_ _07543_ _07544_ vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ op_code\[0\] vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10130_ _00194_ vssd1 vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10061_ _00106_ _00147_ _00150_ _00152_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ _03969_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ _03900_ _03901_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__xnor2_2
X_10963_ _05213_ _04657_ _01054_ _01055_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__nand4_4
X_12702_ _02758_ _02791_ _02794_ vssd1 vssd1 vccd1 vccd1 _02795_ sky130_fd_sc_hd__a21oi_2
X_16470_ _02823_ _02825_ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__nor2_1
X_13682_ _03816_ _03825_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10894_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel _05290_ ApproximateM_inst.lob_16.lob1.genblk1\[13\].genblk1.mux.sel
+ ApproximateM_inst.lob_16.lob1.genblk1\[12\].genblk1.mux.sel vssd1 vssd1 vccd1 vccd1
+ _00987_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15421_ _05722_ _05723_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__nor2_1
X_12633_ _02716_ _02718_ _02719_ _02725_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15352_ _05647_ _05648_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__or2_1
X_18140_ _08676_ vssd1 vssd1 vccd1 vccd1 _08679_ sky130_fd_sc_hd__inv_2
X_12564_ _02611_ _02654_ vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ _04503_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ _01164_ _01163_ _01156_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__a21o_1
X_18071_ _06462_ _08602_ _08603_ vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__or3_1
Xwire131 _03265_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
X_15283_ _05370_ _05487_ _05485_ vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire142 _00850_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_1
X_12495_ _02584_ _02586_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__nor2_1
X_17022_ _08615_ _07459_ _07460_ vssd1 vssd1 vccd1 vccd1 _07462_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14234_ _03596_ _06722_ _05606_ _03629_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _01535_ _01538_ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ _03993_ _04205_ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__or2_1
X_11377_ _01315_ _01419_ vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__and2_1
X_13116_ _03207_ _03208_ _03209_ vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__a21o_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _00418_ _00419_ _00420_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__nand3_2
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _07123_ _04277_ _04278_ vssd1 vssd1 vccd1 vccd1 _04279_ sky130_fd_sc_hd__a21bo_1
X_18973_ clknet_4_5_0_clk _09404_ vssd1 vssd1 vccd1 vccd1 salida\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _08444_ vssd1 vssd1 vccd1 vccd1 _08445_ sky130_fd_sc_hd__inv_2
X_13047_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__inv_2
X_10259_ _07799_ cla_inst.in1\[31\] _09256_ ApproximateM_inst.lob_16.lob2.genblk1\[1\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__a22o_1
X_17855_ _07394_ _07604_ _07665_ _07649_ vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__and4_1
X_16806_ _07122_ _07132_ _07225_ vssd1 vssd1 vccd1 vccd1 _07226_ sky130_fd_sc_hd__a21o_1
X_17786_ _08292_ _08293_ vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__or2_1
X_14998_ _05163_ _05166_ _05164_ vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_88_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16737_ _07049_ _07057_ _07150_ vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__a21o_1
X_13949_ _03954_ _03955_ _04116_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16668_ _00881_ _06433_ vssd1 vssd1 vccd1 vccd1 _07076_ sky130_fd_sc_hd__nor2_1
X_18407_ _08868_ _08917_ vssd1 vssd1 vccd1 vccd1 _08968_ sky130_fd_sc_hd__and2_1
X_15619_ _05938_ _05939_ vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16599_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18338_ _08807_ _08870_ vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_802 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18269_ _02869_ _08760_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09973_ ApproximateM_inst.lob_16.lob1.genblk1\[1\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 _09179_ sky130_fd_sc_hd__buf_4
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11300_ _01389_ _01390_ _01391_ _01382_ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ _01113_ _02259_ vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__nor2_2
XFILLER_0_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11231_ _01319_ _01323_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11162_ cla_inst.in2\[24\] _00174_ _07548_ _07581_ vssd1 vssd1 vccd1 vccd1 _01255_
+ sky130_fd_sc_hd__nand4_1
X_10113_ _00205_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__clkbuf_8
X_11093_ _01183_ _01184_ _01185_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__a21bo_1
X_15970_ _04241_ _04079_ _05623_ vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__and3_1
X_14921_ _05140_ _05056_ _05179_ vssd1 vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__a21oi_2
X_10044_ _00133_ _00136_ vssd1 vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ _08132_ _08133_ _08134_ vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__o21ai_1
X_14852_ _01521_ _00498_ _05101_ _05102_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__and4_1
Xhold83 ApproximateM_inst.lob_16.lob1.genblk1\[3\].genblk1.mux.sel vssd1 vssd1 vccd1
+ vccd1 net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 net96 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _03952_ _03958_ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__xor2_1
X_14783_ _04877_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__xnor2_1
X_17571_ _07143_ _07387_ _08055_ _08057_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__o22a_1
X_11995_ _02083_ _02087_ vssd1 vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__or2_1
X_13734_ _03834_ _03835_ _03882_ _03883_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nor4_1
X_16522_ _02974_ _06916_ vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__nor2_1
X_10946_ _01022_ _01023_ _01038_ vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__and3_4
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13665_ _03805_ _03806_ _03788_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a21o_1
X_16453_ _02980_ _06488_ vssd1 vssd1 vccd1 vccd1 _06843_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10877_ _04351_ _04373_ _03815_ _03837_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _05703_ _05706_ vssd1 vssd1 vccd1 vccd1 _05707_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12616_ _02707_ _02708_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16384_ _06763_ _06767_ vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__nor2_1
X_13596_ _03731_ _03732_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ _01356_ _03055_ _05559_ _05558_ _04900_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18123_ _08616_ _08573_ _08658_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__and3_1
X_12547_ _00832_ _00180_ _02595_ _02596_ vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ _05467_ _05468_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__or2_1
X_18054_ _08502_ _08585_ vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__xnor2_1
X_12478_ _02540_ _02541_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__or2b_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_3 _00166_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ _04401_ _04410_ _04411_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__a21oi_2
X_17005_ _07382_ _07383_ _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ _01520_ _07559_ _07602_ _01521_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_112_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15197_ _02996_ _07025_ _00119_ _02993_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14148_ _00461_ vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18956_ clknet_4_1_0_clk _09417_ vssd1 vssd1 vccd1 vccd1 salida\[9\] sky130_fd_sc_hd__dfxtp_1
X_14079_ _02979_ _04259_ vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__or2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ _02173_ _08423_ _08425_ vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__a21oi_4
X_18887_ clknet_4_11_0_clk _00041_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[5\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17838_ _08265_ _08273_ vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer15 _04574_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_1
Xrebuffer26 _03810_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_107_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer37 _04432_ vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_1
Xrebuffer48 _03004_ vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_1
X_17769_ _08259_ _08166_ _08274_ vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__o21a_1
Xrebuffer59 _05377_ vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09956_ net166 _06906_ _09005_ _09016_ vssd1 vssd1 vccd1 vccd1 _09027_ sky130_fd_sc_hd__o211a_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _07919_ _07930_ _08126_ _08267_ vssd1 vssd1 vccd1 vccd1 _08278_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _00856_ _00891_ _00273_ _00892_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__o211ai_4
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11780_ _00164_ vssd1 vssd1 vccd1 vccd1 _01873_ sky130_fd_sc_hd__buf_6
XFILLER_0_138_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10731_ _00797_ _00821_ _06181_ _00822_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_137_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13450_ _03164_ _03571_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__or2_1
X_10662_ _00752_ _00753_ _00572_ _00598_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12401_ _07984_ _07973_ _00909_ _00145_ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__nand4_2
XFILLER_0_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ _03321_ _00165_ _00212_ _03322_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10593_ _00685_ _00108_ _00511_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15120_ _05310_ _05395_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ _02423_ _02424_ _05671_ _00146_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__and4b_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15051_ _05212_ _05314_ _05319_ vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__nor3_1
X_12263_ _06993_ _00213_ _02354_ _02355_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a31o_1
X_14002_ _00195_ _00702_ _08452_ _04700_ vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__and4_1
X_11214_ _01304_ _01305_ _01291_ _01292_ vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12194_ _02268_ _02275_ _02285_ _02286_ vssd1 vssd1 vccd1 vccd1 _02287_ sky130_fd_sc_hd__a211oi_2
X_18810_ _09298_ _09316_ vssd1 vssd1 vccd1 vccd1 _09317_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11145_ _01147_ _01148_ _01237_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__and3_1
Xoutput73 net73 vssd1 vssd1 vccd1 vccd1 leds[1] sky130_fd_sc_hd__buf_2
Xoutput84 net84 vssd1 vssd1 vccd1 vccd1 o_wb_data[10] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 vssd1 vssd1 vccd1 vccd1 o_wb_data[20] sky130_fd_sc_hd__clkbuf_4
X_18741_ _09262_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__buf_1
X_11076_ _01046_ _01045_ vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__and2b_1
X_15953_ _06284_ _06285_ _06287_ _06269_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__a2bb2o_1
X_14904_ _00191_ _05715_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__and2_1
X_10027_ _07799_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__clkbuf_4
X_18672_ net37 _00593_ _09193_ vssd1 vssd1 vccd1 vccd1 _09213_ sky130_fd_sc_hd__mux2_1
X_15884_ _06192_ _06226_ vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__nor2_1
X_17623_ _08113_ _08114_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__nor2_1
X_14835_ _03059_ _03076_ _03164_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17554_ _08020_ _08022_ _08041_ _06723_ _01862_ vssd1 vssd1 vccd1 vccd1 _09393_ sky130_fd_sc_hd__o32a_1
X_14766_ _05009_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__and2_1
X_11978_ _01944_ _01973_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 _02071_ sky130_fd_sc_hd__nor4_1
X_16505_ _06897_ _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__xor2_2
X_13717_ _00125_ _04143_ _04154_ _00151_ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a22oi_1
X_10929_ _00939_ _00931_ _00938_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__nand3_1
X_14697_ _04934_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__xor2_2
X_17485_ _07823_ _07839_ vssd1 vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16436_ _06822_ _06823_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13648_ _03609_ _03616_ _03615_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13579_ _03697_ _03698_ _03712_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16367_ _06660_ _06663_ _00494_ vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__o21a_4
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ _08640_ vssd1 vssd1 vccd1 vccd1 _08642_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15318_ _05524_ _05525_ _05611_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__nand3_1
X_16298_ _02489_ _00108_ _06673_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__or3_1
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18037_ _07303_ _07861_ _08384_ vssd1 vssd1 vccd1 vccd1 _08567_ sky130_fd_sc_hd__or3_1
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15249_ _03006_ _01695_ vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09810_ _07417_ _07428_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ cla_inst.in1\[22\] vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__buf_4
X_18939_ clknet_4_2_0_clk _00093_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09672_ _05529_ _05867_ _05932_ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__nand3_4
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09939_ _05649_ _06722_ _05704_ _05573_ vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ _03040_ _03042_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__nand2_1
X_11901_ _01747_ _01993_ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__xor2_2
X_12881_ _02973_ vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__clkbuf_4
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _04713_ _04718_ _04712_ vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__a21bo_1
X_11832_ _01922_ _01923_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__a21bo_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _04480_ _04662_ vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__or2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _01852_ _01855_ vssd1 vssd1 vccd1 vccd1 _01856_ sky130_fd_sc_hd__xor2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _03627_ _03628_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__xnor2_1
X_10714_ _06591_ _04569_ _04449_ _00806_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__a22o_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _07703_ _07704_ _07729_ _07730_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__o211a_1
X_14482_ _04598_ _04599_ _04605_ vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand3_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11694_ _01751_ _01785_ _01783_ _01786_ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16221_ _06513_ _06586_ _06587_ _06588_ _06589_ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__a311o_1
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13433_ _03552_ _03554_ _02489_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__mux2_1
X_10645_ _00735_ _00736_ _00719_ _00720_ vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16152_ op_code\[2\] op_code\[3\] vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__and2_2
X_13364_ _01505_ _00557_ _03300_ _03299_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__a31o_1
X_10576_ _07047_ _07080_ _09256_ _09303_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__nand4_2
Xrebuffer6 _03498_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__buf_4
XFILLER_0_24_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15103_ _05273_ _05274_ _05271_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__o21ai_1
X_12315_ _02407_ _02359_ _02358_ vssd1 vssd1 vccd1 vccd1 _02408_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16083_ _03107_ _06440_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__and2_1
X_13295_ _03400_ _03401_ _03396_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__a21o_1
X_15034_ _05302_ _05303_ vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__and2_1
X_12246_ _02246_ _02338_ vssd1 vssd1 vccd1 vccd1 _02339_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12177_ _02268_ _02269_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__nand2_1
X_11128_ _07700_ _05257_ _01220_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__and3_2
X_16985_ _07419_ _07420_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ net59 _09190_ _09249_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11059_ _04078_ _01151_ _00176_ _00145_ vssd1 vssd1 vccd1 vccd1 _01152_ sky130_fd_sc_hd__and4_1
X_15936_ _06242_ _06254_ _06281_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__a21oi_1
X_18655_ _09176_ _09199_ vssd1 vssd1 vccd1 vccd1 _09200_ sky130_fd_sc_hd__and2_1
X_15867_ _06157_ _06205_ _06206_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17606_ _08084_ _08097_ vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__xnor2_1
X_14818_ _05065_ _05066_ _04965_ _04966_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__a211o_1
X_18586_ net297 _09140_ _09148_ _09144_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15798_ _06065_ _06068_ _06133_ vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _02989_ _06510_ _01862_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__a21o_1
X_14749_ _04989_ _04990_ _04991_ vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__nand3_1
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17468_ _07945_ _07946_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16419_ _01151_ ApproximateM_inst.lob_16.lob2.genblk1\[14\].genblk1.mux.sel _03184_
+ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17399_ _07753_ _07754_ _07750_ vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _06450_ _06493_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__xnor2_2
X_09655_ _05715_ vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__buf_4
X_09586_ _04995_ _03935_ _03925_ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__a21oi_2
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_307 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ _00521_ _00522_ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10361_ _00282_ _00285_ _00283_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12100_ _02190_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__or2_1
X_13080_ _03168_ _03171_ _03048_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10292_ _09353_ _00223_ _00238_ _00237_ vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__a31o_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12031_ _01575_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16770_ _03198_ _04257_ _07182_ _07186_ vssd1 vssd1 vccd1 vccd1 _07187_ sky130_fd_sc_hd__a211o_1
X_13982_ _04152_ _00398_ _07526_ _04153_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__and4b_1
X_15721_ _06049_ _05985_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__or2_1
X_12933_ _03025_ vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__clkbuf_4
X_18440_ _08999_ _09002_ vssd1 vssd1 vccd1 vccd1 _09003_ sky130_fd_sc_hd__xnor2_1
X_15652_ _02991_ _09351_ _00495_ _07744_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__nand4_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _02951_ _02956_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__or2b_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14603_ _04726_ _04732_ vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__nand2_2
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _08927_ _08928_ vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__or2_1
X_11815_ _01905_ _01907_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__xnor2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15583_ _00115_ _00495_ vssd1 vssd1 vccd1 vccd1 _05901_ sky130_fd_sc_hd__nand2_1
X_12795_ _01500_ _01499_ _01450_ _01447_ vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__o211a_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _07786_ _07787_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__or2b_1
X_14534_ _04609_ _04699_ _04754_ _04757_ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a211o_1
X_11746_ _01837_ _01838_ vssd1 vssd1 vccd1 vccd1 _01839_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17253_ _06653_ _07486_ _07593_ net331 vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_154_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14465_ _04564_ _04565_ net217 _04682_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__a211oi_4
X_11677_ _01760_ _01761_ _01768_ vssd1 vssd1 vccd1 vccd1 _01770_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ _06571_ vssd1 vssd1 vccd1 vccd1 _06572_ sky130_fd_sc_hd__clkbuf_4
X_10628_ _00545_ _00550_ vssd1 vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__nand2_1
X_13416_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__buf_4
XFILLER_0_126_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14396_ _04598_ net188 _04605_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a21oi_2
X_17184_ _07630_ _07130_ _07521_ _07519_ vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__o31a_1
XFILLER_0_52_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13347_ _03450_ _03451_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__a21oi_1
X_16135_ _03089_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__or2_1
X_10559_ _00649_ _00650_ _00646_ _00472_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13278_ _03881_ _03782_ _08049_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__and3_1
X_16066_ _03239_ _03217_ vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__nand2_2
X_15017_ _05283_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__nand2_1
X_12229_ _02160_ _02159_ vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16968_ _06657_ _07108_ _07292_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__and3_1
X_18707_ net53 _03143_ _09182_ vssd1 vssd1 vccd1 vccd1 _09236_ sky130_fd_sc_hd__mux2_1
X_15919_ _06232_ _06235_ _06263_ vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16899_ _07324_ _07326_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__xnor2_1
X_09440_ _03399_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__buf_6
X_18638_ _09185_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18569_ net261 _09098_ _09135_ _09126_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09707_ _06277_ _06309_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09638_ _05562_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__buf_2
XFILLER_0_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09569_ _04777_ _04799_ _04788_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__a21o_1
X_11600_ _01105_ _00514_ _01692_ _05845_ vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__or4b_4
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12580_ _02644_ _02645_ _02651_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ _01566_ _01567_ _01565_ vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14250_ _04289_ _04291_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _01553_ _01554_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13201_ _03300_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _00496_ _00505_ vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__xnor2_2
X_14181_ _04357_ _04358_ _04371_ vssd1 vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11393_ _01469_ _01485_ vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__xnor2_1
X_13132_ _00294_ _05606_ _05617_ _04351_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10344_ _00276_ _00277_ _00275_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__a21bo_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ _03154_ vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17940_ _08357_ _08460_ vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__nand2_1
X_10275_ _00349_ _00350_ _00367_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a21oi_1
X_12014_ _02090_ _02105_ _02106_ _02050_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__o211a_4
X_17871_ _07630_ _07861_ _08385_ vssd1 vssd1 vccd1 vccd1 _08386_ sky130_fd_sc_hd__nor3_1
X_16822_ _07241_ _07148_ _07242_ vssd1 vssd1 vccd1 vccd1 _07244_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _06989_ _07094_ _07095_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__o21a_1
X_13965_ _04134_ _04135_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__xnor2_1
Xmax_cap4 _02293_ vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__clkbuf_1
X_15704_ _03007_ _03055_ _06031_ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__nand3_1
X_12916_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__buf_2
X_16684_ _03790_ _06509_ _02214_ vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__a21oi_1
X_13896_ _03847_ _03849_ _03852_ _03854_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__a31oi_2
X_18423_ _02920_ net115 _03201_ vssd1 vssd1 vccd1 vccd1 _08986_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15635_ _05929_ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__inv_2
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ _02939_ vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__inv_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _08909_ _08910_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__xnor2_1
X_15566_ _03007_ _01112_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__nand2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _02869_ _02870_ vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17305_ _07618_ _07642_ _07617_ vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__o21ba_1
X_14517_ _04702_ _04703_ _04737_ _04738_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_84_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18285_ _08751_ _08813_ _08814_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__o21ba_1
X_11729_ ApproximateM_inst.lob_16.lob2.genblk1\[11\].genblk1.mux.sel _00177_ vssd1
+ vssd1 vccd1 vccd1 _01822_ sky130_fd_sc_hd__nand2_1
X_15497_ _02975_ _05805_ _05806_ vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17236_ _06368_ _06438_ _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14448_ _04651_ _04652_ _04663_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17167_ _07617_ _07618_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14379_ _02188_ _09256_ _07755_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16118_ _03029_ _01746_ _01503_ _03083_ _06477_ _03161_ vssd1 vssd1 vccd1 vccd1 _06478_
+ sky130_fd_sc_hd__mux4_1
X_17098_ _06665_ _07314_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16049_ _01417_ _03143_ vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__or2_2
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _03217_ _03206_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10060_ _09352_ _00147_ _00150_ _00152_ vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__nand4_1
X_13750_ _03732_ _03735_ _03731_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__o21ba_2
X_10962_ _06591_ _03804_ _03826_ _00806_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _02792_ _02793_ vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__and2_1
X_13681_ _03823_ _03824_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__and2_1
X_10893_ _05290_ _03739_ _03804_ ApproximateM_inst.lob_16.lob2.genblk1\[10\].genblk1.mux.sel
+ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__a22o_1
X_15420_ _02991_ _08876_ _05721_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12632_ _02722_ _02723_ _02724_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15351_ _05569_ _05567_ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _02618_ _02625_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14302_ _01745_ _04336_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__nand2_1
X_11514_ _01164_ _01156_ _01163_ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__nand3_1
XFILLER_0_80_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18070_ _07002_ _08036_ _03197_ _05881_ vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__a2bb2o_1
X_15282_ _05571_ _05572_ vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__nand2_1
X_12494_ _02584_ _02586_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire132 _08451_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17021_ _07386_ _07355_ _00399_ vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__o21a_1
X_14233_ _04283_ net133 _04295_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__nor3_2
X_11445_ _06460_ _00878_ _01536_ _01537_ _00193_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__a32o_1
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14164_ _04337_ _04353_ vssd1 vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11376_ _01409_ _01411_ _01407_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ _03207_ _03208_ _03209_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__nand3_1
X_10327_ _00245_ _00267_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__nand2_1
X_14095_ _04132_ _07156_ _06732_ _04099_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a22o_1
X_18972_ clknet_4_5_0_clk _09403_ vssd1 vssd1 vccd1 vccd1 salida\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _08434_ _08436_ _08439_ _08443_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__and4b_1
X_13046_ _03135_ _03137_ _03048_ vssd1 vssd1 vccd1 vccd1 _03138_ sky130_fd_sc_hd__mux2_1
X_10258_ _07700_ _07799_ cla_inst.in1\[31\] _09256_ vssd1 vssd1 vccd1 vccd1 _00351_
+ sky130_fd_sc_hd__nand4_1
X_17854_ _07608_ _07314_ _07516_ _07195_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__o22a_1
X_10189_ _04121_ _04580_ _04460_ _04088_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a22oi_2
X_16805_ _07121_ _07119_ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__and2b_1
X_17785_ _08257_ _08258_ _08291_ vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__and3_1
X_14997_ _05168_ _05167_ vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__or2b_1
X_16736_ _07017_ _07048_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nor2_1
X_13948_ _03954_ _03955_ _04116_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16667_ _02800_ _07073_ _07074_ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__o21a_1
X_13879_ _04025_ _04026_ _04040_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__and3_1
XFILLER_0_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18406_ _08965_ _08966_ vssd1 vssd1 vccd1 vccd1 _08967_ sky130_fd_sc_hd__xor2_1
X_15618_ _05861_ net118 _05937_ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16598_ _06696_ _06701_ _03060_ vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18337_ _03143_ _06464_ _08839_ _08892_ vssd1 vssd1 vccd1 vccd1 _09404_ sky130_fd_sc_hd__o2bb2a_1
X_15549_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18268_ _08815_ _08816_ _08817_ vssd1 vssd1 vccd1 vccd1 _08818_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17219_ _02669_ _02670_ _07562_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__o21a_1
X_18199_ _08587_ _08742_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ cla_inst.in2\[29\] vssd1 vssd1 vccd1 vccd1 _09172_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11230_ _01320_ _01322_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ cla_inst.in2\[22\] _09212_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10112_ _04220_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__clkbuf_8
X_11092_ _05508_ _05464_ _04143_ _04056_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__nand4_1
X_14920_ _05161_ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__xnor2_1
X_10043_ _09353_ _00134_ _00135_ _00128_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__a22oi_1
X_14851_ _02986_ _07733_ _05101_ _05102_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__a22oi_4
Xhold84 op_code\[1\] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_1
Xhold95 _00025_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _03955_ _03956_ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _07143_ _07387_ _08055_ _08057_ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__nor4_1
X_14782_ _05018_ _05027_ vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11994_ _02084_ _02085_ _02086_ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__o21ba_1
X_16521_ _06639_ _06632_ _06627_ _06641_ _03080_ _03077_ vssd1 vssd1 vccd1 vccd1 _06916_
+ sky130_fd_sc_hd__mux4_2
X_13733_ _03879_ _03880_ _03836_ _03715_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10945_ _01028_ _01036_ _01037_ vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16452_ _06839_ _06840_ vssd1 vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__xnor2_1
X_13664_ _03788_ _03805_ _03806_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__nand3_2
X_10876_ _05017_ _03750_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ _05705_ _05591_ _05588_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12615_ _02705_ _02706_ _02701_ _02704_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__o211a_1
X_16383_ _06579_ _06653_ _06766_ _06561_ vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__o22a_1
X_13595_ _03518_ _03521_ _03730_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_93_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ _08616_ _08573_ _08658_ vssd1 vssd1 vccd1 vccd1 _08660_ sky130_fd_sc_hd__a21oi_1
X_15334_ _05556_ _05565_ vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ _02636_ _02637_ _02638_ vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18053_ _08582_ _08584_ vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__or2_1
X_15265_ _05476_ _05473_ vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__and2b_1
X_12477_ _02568_ _02569_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__or2_1
XFILLER_0_151_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _00181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _07434_ _07441_ vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__xnor2_1
X_14216_ _04401_ _04410_ _03202_ vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__o21ai_1
X_11428_ _03574_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__buf_4
X_15196_ _05478_ _05479_ vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14147_ _04148_ _04163_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__nand2_1
X_11359_ _01436_ _01416_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18955_ clknet_4_1_0_clk _09416_ vssd1 vssd1 vccd1 vccd1 salida\[8\] sky130_fd_sc_hd__dfxtp_1
X_14078_ _03567_ _03581_ _02980_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__mux2_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _02976_ _03035_ _03039_ _03118_ _03121_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__o32a_1
X_17906_ _04238_ _08424_ vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__or2_1
X_18886_ clknet_4_13_0_clk _00040_ vssd1 vssd1 vccd1 vccd1 ApproximateM_inst.lob_16.lob1.genblk1\[4\].genblk1.mux.sel
+ sky130_fd_sc_hd__dfxtp_1
X_17837_ _08263_ _08264_ vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer16 _04574_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_1
Xrebuffer27 net337 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_1
Xrebuffer38 _04432_ vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_1
XFILLER_0_107_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17768_ _08265_ _08273_ vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xrebuffer49 _03004_ vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_1
XFILLER_0_107_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16719_ _06579_ _07130_ vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17699_ _08074_ _08076_ _08197_ vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__nor3_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09955_ _08973_ _08984_ _08995_ _08681_ vssd1 vssd1 vccd1 vccd1 _09016_ sky130_fd_sc_hd__a22o_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _08126_ _08137_ _08256_ vssd1 vssd1 vccd1 vccd1 _08267_ sky130_fd_sc_hd__nand3_2
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10730_ _00797_ _00821_ _06181_ _00822_ vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__o211a_2
XFILLER_0_138_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ _00572_ _00598_ _00752_ _00753_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_138_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _07243_ _00176_ _00145_ _07221_ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__a22o_1
X_13380_ _03270_ _03272_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10592_ cla_inst.in2\[31\] _00108_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12331_ _08039_ _00196_ _09212_ _00992_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15050_ _05212_ _05314_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__o21a_1
X_12262_ _07984_ _07243_ _04220_ _00774_ vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__and4_1
X_11213_ _01291_ _01292_ _01304_ _01305_ vssd1 vssd1 vccd1 vccd1 _01306_ sky130_fd_sc_hd__o211ai_2
X_14001_ _00702_ _08452_ _01005_ _00195_ vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__a22oi_2
X_12193_ _02195_ _02198_ _02284_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11144_ _01204_ _01236_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__or2b_1
Xoutput74 net74 vssd1 vssd1 vccd1 vccd1 leds[2] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 vssd1 vssd1 vccd1 vccd1 o_wb_data[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput96 net96 vssd1 vssd1 vccd1 vccd1 o_wb_data[21] sky130_fd_sc_hd__clkbuf_4
X_18740_ _09245_ _09261_ vssd1 vssd1 vccd1 vccd1 _09262_ sky130_fd_sc_hd__and2_1
X_11075_ _04548_ _04056_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__nand2_1
X_15952_ _06232_ _06235_ _06263_ _06297_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__a211o_1
X_14903_ _05158_ _05160_ vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__nor2_1
X_10026_ _08876_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__buf_4
X_18671_ _09211_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__buf_1
X_15883_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__inv_2
X_17622_ _08113_ _08114_ vssd1 vssd1 vccd1 vccd1 _08116_ sky130_fd_sc_hd__and2_1
X_14834_ _03921_ _05085_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17553_ _07256_ _08027_ _08029_ _08040_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__a31o_1
X_14765_ _05001_ _05008_ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11977_ _02052_ _02068_ _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__or3_2
X_16504_ _06824_ _06827_ _06822_ vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__o21a_1
X_13716_ _03654_ _03656_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17484_ _07954_ _07964_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__xnor2_1
X_10928_ _00980_ _01019_ _01018_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14696_ _04798_ _04801_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16435_ _06769_ _06821_ vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__nand2_1
X_13647_ _03637_ _03639_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nand2_1
X_10859_ _04558_ _04045_ _00950_ _00951_ vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _03539_ _06734_ _06747_ _06484_ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__o211a_1
X_13578_ _03697_ _03698_ _03712_ vssd1 vssd1 vccd1 vccd1 _03713_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18105_ _08639_ _07859_ _07109_ _08640_ vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__and4b_1
XFILLER_0_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _05524_ _05525_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__a21o_1
X_12529_ _02615_ _02619_ _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__and3_1
X_16297_ _06585_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__buf_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18036_ _08470_ _08479_ vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__or2b_1
X_15248_ _05534_ _05535_ vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15179_ _05237_ _05359_ vssd1 vssd1 vccd1 vccd1 _05461_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09740_ _05573_ _05595_ _05693_ _05606_ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__and4_1
X_18938_ clknet_4_11_0_clk _00092_ vssd1 vssd1 vccd1 vccd1 cla_inst.in2\[24\] sky130_fd_sc_hd__dfxtp_2
.ends

