* NGSPICE file created from egd_top_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

.subckt egd_top_wrapper la_data_in_58_43[0] la_data_in_58_43[10] la_data_in_58_43[11]
+ la_data_in_58_43[12] la_data_in_58_43[13] la_data_in_58_43[14] la_data_in_58_43[15]
+ la_data_in_58_43[1] la_data_in_58_43[2] la_data_in_58_43[3] la_data_in_58_43[4]
+ la_data_in_58_43[5] la_data_in_58_43[6] la_data_in_58_43[7] la_data_in_58_43[8]
+ la_data_in_58_43[9] la_data_in_60_59[0] la_data_in_60_59[1] la_data_in_65 la_data_out_23_16[0]
+ la_data_out_23_16[1] la_data_out_23_16[2] la_data_out_23_16[3] la_data_out_23_16[4]
+ la_data_out_23_16[5] la_data_out_23_16[6] la_data_out_23_16[7] la_data_out_26_24[0]
+ la_data_out_26_24[1] la_data_out_26_24[2] la_data_out_30_27[0] la_data_out_30_27[1]
+ la_data_out_30_27[2] la_data_out_30_27[3] vccd1 vssd1 wb_clk_i
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6914_ net35 _0317_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__dfxtp_2
X_6845_ net43 _0248_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[31\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3988_ _0473_ vssd1 vssd1 vccd1 vccd1 _0474_ sky130_fd_sc_hd__buf_4
XFILLER_0_64_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6776_ net130 _0179_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5727_ _0708_ _0385_ _2199_ vssd1 vssd1 vccd1 vccd1 _2200_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5658_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1 vccd1
+ _2132_ sky130_fd_sc_hd__inv_2
X_4609_ _0334_ _0380_ vssd1 vssd1 vccd1 vccd1 _1091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5589_ _0634_ _3349_ vssd1 vssd1 vccd1 vccd1 _2063_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4960_ _3258_ _0804_ vssd1 vssd1 vccd1 vccd1 _1439_ sky130_fd_sc_hd__nand2_1
X_4891_ _1360_ _1364_ _1367_ _1370_ vssd1 vssd1 vccd1 vccd1 _1371_ sky130_fd_sc_hd__and4_1
X_3911_ _0396_ vssd1 vssd1 vccd1 vccd1 _0397_ sky130_fd_sc_hd__clkbuf_4
X_3842_ _0327_ vssd1 vssd1 vccd1 vccd1 _0328_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6561_ _2894_ _2713_ vssd1 vssd1 vccd1 vccd1 _2895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5512_ _0482_ _0488_ _0535_ _0492_ _1986_ vssd1 vssd1 vccd1 vccd1 _1987_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3773_ _3306_ vssd1 vssd1 vccd1 vccd1 _3307_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6492_ _1652_ _2707_ _2827_ vssd1 vssd1 vccd1 vccd1 _2828_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5443_ _0554_ _3218_ _0745_ _3221_ vssd1 vssd1 vccd1 vccd1 _1918_ sky130_fd_sc_hd__o22ai_1
X_5374_ _0416_ _3095_ vssd1 vssd1 vccd1 vccd1 _1850_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4325_ _3318_ _3281_ _3322_ _3285_ _0808_ vssd1 vssd1 vccd1 vccd1 _0809_ sky130_fd_sc_hd__a221oi_1
X_4256_ _0727_ _0731_ _0736_ _0740_ vssd1 vssd1 vccd1 vccd1 _0741_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4187_ _0671_ _3350_ vssd1 vssd1 vccd1 vccd1 _0672_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6828_ net182 _0231_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[48\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6759_ net113 _0162_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[94\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6657__145 clknet_1_1__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__inv_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6692__21 clknet_1_1__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__inv_2
X_5090_ _1444_ _3289_ _3348_ _3293_ vssd1 vssd1 vccd1 vccd1 _1568_ sky130_fd_sc_hd__o22ai_1
X_4110_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _0596_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4041_ _0526_ vssd1 vssd1 vccd1 vccd1 _0527_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5992_ net13 _0475_ _2415_ vssd1 vssd1 vccd1 vccd1 _2435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4943_ _1410_ _1413_ _1417_ _1421_ vssd1 vssd1 vccd1 vccd1 _1422_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4874_ _0394_ _0386_ _1353_ vssd1 vssd1 vccd1 vccd1 _1354_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3825_ _3358_ vssd1 vssd1 vccd1 vccd1 _3359_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6544_ _2831_ _2877_ vssd1 vssd1 vccd1 vccd1 _2878_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3756_ egd_top.BitStream_buffer.BS_buffer\[93\] vssd1 vssd1 vccd1 vccd1 _3290_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6475_ _2812_ _2815_ vssd1 vssd1 vccd1 vccd1 _2816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5426_ _3128_ _3149_ vssd1 vssd1 vccd1 vccd1 _1901_ sky130_fd_sc_hd__nand2_1
X_3687_ _3220_ vssd1 vssd1 vccd1 vccd1 _3221_ sky130_fd_sc_hd__clkbuf_4
X_5357_ _0338_ _0429_ vssd1 vssd1 vccd1 vccd1 _1833_ sky130_fd_sc_hd__nand2_1
X_5288_ _0867_ _0561_ _1762_ _1763_ _1764_ vssd1 vssd1 vccd1 vccd1 _1765_ sky130_fd_sc_hd__o2111a_1
X_4308_ _0607_ _3212_ _0577_ _3215_ _0791_ vssd1 vssd1 vccd1 vccd1 _0792_ sky130_fd_sc_hd__a221oi_1
X_4239_ _0474_ _0479_ vssd1 vssd1 vccd1 vccd1 _0724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6729__55 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__inv_2
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6744__69 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__inv_2
X_4590_ _1060_ _1065_ _1068_ _1071_ vssd1 vssd1 vccd1 vccd1 _1072_ sky130_fd_sc_hd__and4_1
X_3610_ egd_top.BitStream_buffer.BS_buffer\[78\] vssd1 vssd1 vccd1 vccd1 _3144_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3541_ _3074_ vssd1 vssd1 vccd1 vccd1 _3075_ sky130_fd_sc_hd__buf_4
XFILLER_0_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3472_ _3018_ vssd1 vssd1 vccd1 vccd1 _0310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6260_ _2617_ vssd1 vssd1 vccd1 vccd1 _0175_ sky130_fd_sc_hd__clkbuf_1
X_6191_ net15 _3335_ _2557_ vssd1 vssd1 vccd1 vccd1 _2572_ sky130_fd_sc_hd__mux2_1
X_5211_ _3271_ _3282_ _3274_ _3318_ vssd1 vssd1 vccd1 vccd1 _1688_ sky130_fd_sc_hd__a22o_1
X_5142_ _0474_ _0363_ vssd1 vssd1 vccd1 vccd1 _1620_ sky130_fd_sc_hd__nand2_1
X_5073_ _0607_ _3184_ _0577_ _3187_ _1550_ vssd1 vssd1 vccd1 vccd1 _1551_ sky130_fd_sc_hd__a221oi_1
X_4024_ _0508_ _0509_ vssd1 vssd1 vccd1 vccd1 _0510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5975_ _2422_ _2423_ vssd1 vssd1 vccd1 vccd1 _2424_ sky130_fd_sc_hd__and2_1
X_4926_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] vssd1 vssd1 vccd1 vccd1
+ _1406_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4857_ _3365_ _3019_ vssd1 vssd1 vccd1 vccd1 _1337_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3808_ _3340_ _3341_ vssd1 vssd1 vccd1 vccd1 _3342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6527_ _2831_ _2859_ _2829_ vssd1 vssd1 vccd1 vccd1 _2862_ sky130_fd_sc_hd__nand3_1
X_4788_ _0750_ _0545_ _1266_ _1267_ _1268_ vssd1 vssd1 vccd1 vccd1 _1269_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3739_ _3122_ _3228_ vssd1 vssd1 vccd1 vccd1 _3273_ sky130_fd_sc_hd__and2_1
X_6458_ _2796_ _2798_ vssd1 vssd1 vccd1 vccd1 _2799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5409_ _0516_ _0561_ _1882_ _1883_ _1884_ vssd1 vssd1 vccd1 vccd1 _1885_ sky130_fd_sc_hd__o2111a_1
X_6389_ _2727_ _2731_ _2710_ vssd1 vssd1 vccd1 vccd1 _2732_ sky130_fd_sc_hd__nand3_1
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5760_ _0329_ _0523_ _0376_ _0527_ _2232_ vssd1 vssd1 vccd1 vccd1 _2233_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4711_ _1188_ _1189_ _1190_ _1191_ vssd1 vssd1 vccd1 vccd1 _1192_ sky130_fd_sc_hd__and4_1
X_5691_ _3257_ _3282_ vssd1 vssd1 vccd1 vccd1 _2164_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4642_ _0474_ _0531_ vssd1 vssd1 vccd1 vccd1 _1124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _3025_ _3198_ _3028_ _3201_ _1054_ vssd1 vssd1 vccd1 vccd1 _1055_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_21_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3524_ _2961_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _3058_ sky130_fd_sc_hd__nand2_2
X_6312_ _2654_ _1282_ vssd1 vssd1 vccd1 vccd1 _2655_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6243_ _2607_ vssd1 vssd1 vccd1 vccd1 _0180_ sky130_fd_sc_hd__inv_2
X_3455_ _2978_ _3004_ vssd1 vssd1 vccd1 vccd1 _3005_ sky130_fd_sc_hd__or2_1
X_6174_ _2560_ _2554_ vssd1 vssd1 vccd1 vccd1 _2561_ sky130_fd_sc_hd__and2_1
X_3386_ _2939_ _2941_ vssd1 vssd1 vccd1 vccd1 _2942_ sky130_fd_sc_hd__nor2_1
X_5125_ _0399_ _0461_ vssd1 vssd1 vccd1 vccd1 _1603_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ _3259_ _3068_ _3251_ _3075_ _1533_ vssd1 vssd1 vccd1 vccd1 _1534_ sky130_fd_sc_hd__a221oi_1
X_4007_ egd_top.BitStream_buffer.BS_buffer\[18\] vssd1 vssd1 vccd1 vccd1 _0493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5958_ _2411_ vssd1 vssd1 vccd1 vccd1 _0265_ sky130_fd_sc_hd__clkbuf_1
X_4909_ _1377_ _1380_ _1384_ _1388_ vssd1 vssd1 vccd1 vccd1 _1389_ sky130_fd_sc_hd__and4_1
X_5889_ _0723_ _0560_ _2358_ _2359_ _2360_ vssd1 vssd1 vccd1 vccd1 _2361_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6708__36 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__inv_2
XFILLER_0_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _2369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6861_ net59 _0264_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[15\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6792_ net146 _0195_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[100\]
+ sky130_fd_sc_hd__dfxtp_1
X_5812_ _2280_ _2281_ _2282_ _2283_ vssd1 vssd1 vccd1 vccd1 _2284_ sky130_fd_sc_hd__and4_1
X_5743_ _3085_ _0449_ _3057_ _0453_ _2215_ vssd1 vssd1 vccd1 vccd1 _2216_ sky130_fd_sc_hd__a221oi_1
X_5674_ _2135_ _2138_ _2142_ _2146_ vssd1 vssd1 vccd1 vccd1 _2147_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4625_ _0403_ _0417_ vssd1 vssd1 vccd1 vccd1 _1107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4556_ _3128_ _3076_ vssd1 vssd1 vccd1 vccd1 _1038_ sky130_fd_sc_hd__nand2_1
X_3507_ net10 _3044_ _3006_ vssd1 vssd1 vccd1 vccd1 _3045_ sky130_fd_sc_hd__mux2_1
X_4487_ _0371_ _0353_ vssd1 vssd1 vccd1 vccd1 _0970_ sky130_fd_sc_hd__nand2_1
X_3438_ _2949_ _2951_ vssd1 vssd1 vccd1 vccd1 _2991_ sky130_fd_sc_hd__nor2_1
X_6226_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2598_ sky130_fd_sc_hd__or2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _2548_ vssd1 vssd1 vccd1 vccd1 _0203_ sky130_fd_sc_hd__clkbuf_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _1574_ _1578_ _1582_ _1585_ vssd1 vssd1 vccd1 vccd1 _1586_ sky130_fd_sc_hd__and4_1
X_6088_ net15 _0701_ _2486_ vssd1 vssd1 vccd1 vccd1 _2501_ sky130_fd_sc_hd__mux2_1
X_5039_ _0563_ _0489_ vssd1 vssd1 vccd1 vccd1 _1518_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[0] sky130_fd_sc_hd__buf_12
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[0] sky130_fd_sc_hd__buf_12
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4410_ _0861_ _0879_ _0893_ vssd1 vssd1 vccd1 vccd1 _0894_ sky130_fd_sc_hd__and3_1
X_5390_ _0498_ _0531_ vssd1 vssd1 vccd1 vccd1 _1866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4341_ _0634_ _3363_ _0824_ vssd1 vssd1 vccd1 vccd1 _0825_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4272_ _0596_ _0595_ _0756_ _0598_ vssd1 vssd1 vccd1 vccd1 _0757_ sky130_fd_sc_hd__o22ai_1
X_6011_ _2932_ vssd1 vssd1 vccd1 vccd1 _2448_ sky130_fd_sc_hd__buf_2
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6913_ net111 _0316_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_76_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6844_ net42 _0247_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[32\]
+ sky130_fd_sc_hd__dfxtp_1
X_3987_ _3090_ _0470_ vssd1 vssd1 vccd1 vccd1 _0473_ sky130_fd_sc_hd__and2_1
X_6775_ net129 _0178_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5726_ _0387_ _0411_ vssd1 vssd1 vccd1 vccd1 _2199_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5657_ _2069_ _2129_ _2130_ vssd1 vssd1 vccd1 vccd1 _2131_ sky130_fd_sc_hd__nand3_2
X_6611__102 clknet_1_0__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__inv_2
X_5588_ _3343_ _3013_ vssd1 vssd1 vccd1 vccd1 _2062_ sky130_fd_sc_hd__nand2_1
X_4608_ _1046_ _1058_ _1072_ _1089_ vssd1 vssd1 vccd1 vccd1 _1090_ sky130_fd_sc_hd__and4_1
XFILLER_0_7_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4539_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1022_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6209_ _2584_ vssd1 vssd1 vccd1 vccd1 _0187_ sky130_fd_sc_hd__clkbuf_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_524 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3910_ _3139_ _0395_ vssd1 vssd1 vccd1 vccd1 _0396_ sky130_fd_sc_hd__nand2_1
X_4890_ _3095_ _0450_ _3102_ _0454_ _1369_ vssd1 vssd1 vccd1 vccd1 _1370_ sky130_fd_sc_hd__a221oi_1
X_3841_ _0326_ vssd1 vssd1 vccd1 vccd1 _0327_ sky130_fd_sc_hd__buf_1
X_6560_ _2891_ _2893_ vssd1 vssd1 vccd1 vccd1 _2894_ sky130_fd_sc_hd__nand2_1
X_3772_ _3305_ vssd1 vssd1 vccd1 vccd1 _3306_ sky130_fd_sc_hd__buf_1
X_5511_ _1249_ _0496_ _1985_ vssd1 vssd1 vccd1 vccd1 _1986_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_502 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6491_ _2707_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1
+ vccd1 _2827_ sky130_fd_sc_hd__nand2_1
X_6634__124 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__inv_2
X_5442_ _3047_ _3198_ _3050_ _3201_ _1916_ vssd1 vssd1 vccd1 vccd1 _1917_ sky130_fd_sc_hd__a221oi_1
X_5373_ _0456_ _0397_ _1846_ _1847_ _1848_ vssd1 vssd1 vccd1 vccd1 _1849_ sky130_fd_sc_hd__o2111a_1
X_4324_ _0656_ _3289_ _0807_ _3293_ vssd1 vssd1 vccd1 vccd1 _0808_ sky130_fd_sc_hd__o22ai_1
X_4255_ _0525_ _0524_ _0359_ _0528_ _0739_ vssd1 vssd1 vccd1 vccd1 _0740_ sky130_fd_sc_hd__a221oi_1
X_4186_ _3345_ vssd1 vssd1 vccd1 vccd1 _0671_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6827_ net181 _0230_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[49\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6758_ net112 _0161_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[95\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5709_ _0786_ _3349_ vssd1 vssd1 vccd1 vccd1 _2182_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4040_ _2964_ _0469_ vssd1 vssd1 vccd1 vccd1 _0526_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__2919_ clknet_0__2919_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2919_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5991_ _2434_ vssd1 vssd1 vccd1 vccd1 _0255_ sky130_fd_sc_hd__clkbuf_1
X_4942_ _3265_ _3148_ _3272_ _3152_ _1420_ vssd1 vssd1 vccd1 vccd1 _1421_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4873_ _0388_ _0404_ vssd1 vssd1 vccd1 vccd1 _1353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3824_ _3153_ _3299_ vssd1 vssd1 vccd1 vccd1 _3358_ sky130_fd_sc_hd__and2_1
X_6543_ _2859_ _2828_ vssd1 vssd1 vccd1 vccd1 _2877_ sky130_fd_sc_hd__nor2_1
X_3755_ _3288_ vssd1 vssd1 vccd1 vccd1 _3289_ sky130_fd_sc_hd__clkbuf_4
X_6474_ _2790_ _2788_ _2814_ vssd1 vssd1 vccd1 vccd1 _2815_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3686_ _3153_ _3167_ vssd1 vssd1 vccd1 vccd1 _3220_ sky130_fd_sc_hd__nand2_1
X_5425_ _3156_ _3101_ _3144_ _3106_ _1899_ vssd1 vssd1 vccd1 vccd1 _1900_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5356_ _0334_ _0433_ vssd1 vssd1 vccd1 vccd1 _1832_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5287_ _0494_ _0570_ vssd1 vssd1 vccd1 vccd1 _1764_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4307_ _0638_ _3218_ _0790_ _3221_ vssd1 vssd1 vccd1 vccd1 _0791_ sky130_fd_sc_hd__o22ai_1
X_4238_ _0475_ vssd1 vssd1 vccd1 vccd1 _0723_ sky130_fd_sc_hd__inv_2
X_4169_ _3271_ _3275_ _3274_ _0653_ vssd1 vssd1 vccd1 vccd1 _0654_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6663__150 clknet_1_1__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__inv_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3540_ _3073_ vssd1 vssd1 vccd1 vccd1 _3074_ sky130_fd_sc_hd__buf_1
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3471_ _3017_ _2933_ vssd1 vssd1 vccd1 vccd1 _3018_ sky130_fd_sc_hd__and2_1
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5210_ _3291_ _3264_ _0656_ _3268_ vssd1 vssd1 vccd1 vccd1 _1687_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6190_ _2571_ vssd1 vssd1 vccd1 vccd1 _0193_ sky130_fd_sc_hd__clkbuf_1
X_5141_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _1619_ sky130_fd_sc_hd__inv_2
X_5072_ _0582_ _3190_ _1549_ vssd1 vssd1 vccd1 vccd1 _1550_ sky130_fd_sc_hd__o21ai_1
X_4023_ egd_top.BitStream_buffer.BS_buffer\[22\] vssd1 vssd1 vccd1 vccd1 _0509_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5974_ _2932_ vssd1 vssd1 vccd1 vccd1 _2423_ sky130_fd_sc_hd__buf_2
X_4925_ _1341_ _1403_ _1404_ vssd1 vssd1 vccd1 vccd1 _1405_ sky130_fd_sc_hd__nand3_1
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4856_ _1332_ _3338_ _1333_ _1334_ _1335_ vssd1 vssd1 vccd1 vccd1 _1336_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _3341_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6526_ _2858_ _2860_ vssd1 vssd1 vccd1 vccd1 _2861_ sky130_fd_sc_hd__nand2_1
X_4787_ _0593_ _0556_ vssd1 vssd1 vccd1 vccd1 _1268_ sky130_fd_sc_hd__or2_1
X_3738_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _3272_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6457_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] _2707_ _2797_ vssd1
+ vssd1 vccd1 vccd1 _2798_ sky130_fd_sc_hd__o21ai_1
X_3669_ _3109_ _3167_ vssd1 vssd1 vccd1 vccd1 _3203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5408_ _0728_ _0570_ vssd1 vssd1 vccd1 vccd1 _1884_ sky130_fd_sc_hd__or2_1
X_6388_ _2709_ _2730_ vssd1 vssd1 vccd1 vccd1 _2731_ sky130_fd_sc_hd__nand2_1
X_5339_ _3309_ _3016_ vssd1 vssd1 vccd1 vccd1 _1815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4710_ _3258_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _1191_
+ sky130_fd_sc_hd__nand2_1
X_5690_ _3253_ _3290_ vssd1 vssd1 vccd1 vccd1 _2163_ sky130_fd_sc_hd__nand2_1
X_4641_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _1123_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4572_ _3174_ _3204_ _1053_ vssd1 vssd1 vccd1 vccd1 _1054_ sky130_fd_sc_hd__o21ai_1
X_6311_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] _2653_ vssd1 vssd1
+ vccd1 vccd1 _2654_ sky130_fd_sc_hd__nor2_1
X_3523_ egd_top.BitStream_buffer.BS_buffer\[74\] vssd1 vssd1 vccd1 vccd1 _3057_ sky130_fd_sc_hd__clkbuf_4
X_6242_ _2989_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _2607_ sky130_fd_sc_hd__nand2_1
X_3454_ _2971_ _3003_ vssd1 vssd1 vccd1 vccd1 _3004_ sky130_fd_sc_hd__or2_1
X_6173_ net6 _3322_ _2557_ vssd1 vssd1 vccd1 vccd1 _2560_ sky130_fd_sc_hd__mux2_1
X_3385_ _2930_ _2940_ vssd1 vssd1 vccd1 vccd1 _2941_ sky130_fd_sc_hd__nor2_1
X_5124_ _1591_ _1595_ _1598_ _1601_ vssd1 vssd1 vccd1 vccd1 _1602_ sky130_fd_sc_hd__and4_1
X_5055_ _1408_ _3084_ _1532_ _3092_ vssd1 vssd1 vccd1 vccd1 _1533_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4006_ _0491_ vssd1 vssd1 vccd1 vccd1 _0492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5957_ _2410_ _2396_ vssd1 vssd1 vccd1 vccd1 _2411_ sky130_fd_sc_hd__and2_1
X_4908_ _0691_ _0524_ _0346_ _0528_ _1387_ vssd1 vssd1 vccd1 vccd1 _1388_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5888_ _0504_ _0569_ vssd1 vssd1 vccd1 vccd1 _2360_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4839_ _1317_ _1318_ vssd1 vssd1 vccd1 vccd1 _1319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6509_ _2842_ _2844_ _2713_ vssd1 vssd1 vccd1 vccd1 _2845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6860_ net58 _0263_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[16\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_88_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6791_ net145 _0194_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[101\]
+ sky130_fd_sc_hd__dfxtp_1
X_5811_ _3257_ _3318_ vssd1 vssd1 vccd1 vccd1 _2283_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5742_ _0900_ _0457_ _2214_ vssd1 vssd1 vccd1 vccd1 _2215_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5673_ _3232_ _3147_ _3286_ _3151_ _2145_ vssd1 vssd1 vccd1 vccd1 _2146_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_44_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4624_ _0399_ _0421_ vssd1 vssd1 vccd1 vccd1 _1106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4555_ _3134_ _3101_ _3119_ _3106_ _1036_ vssd1 vssd1 vccd1 vccd1 _1037_ sky130_fd_sc_hd__a221oi_1
X_3506_ egd_top.BitStream_buffer.BS_buffer\[124\] vssd1 vssd1 vccd1 vccd1 _3044_ sky130_fd_sc_hd__clkbuf_4
X_4486_ _0967_ _0968_ vssd1 vssd1 vccd1 vccd1 _0969_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3437_ _2952_ _2988_ _2989_ _2990_ vssd1 vssd1 vccd1 vccd1 _0317_ sky130_fd_sc_hd__o211a_1
X_6225_ _2594_ _2595_ _2596_ vssd1 vssd1 vccd1 vccd1 _2597_ sky130_fd_sc_hd__a21bo_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _2547_ _2529_ vssd1 vssd1 vccd1 vccd1 _2548_ sky130_fd_sc_hd__and2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5107_ _3019_ _3356_ _3022_ _3360_ _1584_ vssd1 vssd1 vccd1 vccd1 _1585_ sky130_fd_sc_hd__a221oi_1
X_6087_ _2500_ vssd1 vssd1 vccd1 vccd1 _0225_ sky130_fd_sc_hd__clkbuf_1
X_5038_ _0593_ _0545_ _1514_ _1515_ _1516_ vssd1 vssd1 vccd1 vccd1 _1517_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[1] sky130_fd_sc_hd__buf_12
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[1] sky130_fd_sc_hd__buf_12
XFILLER_0_53_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6699__28 clknet_1_0__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__inv_2
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _3365_ _2998_ vssd1 vssd1 vccd1 vccd1 _0824_ sky130_fd_sc_hd__nand2_1
X_4271_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _0756_ sky130_fd_sc_hd__inv_2
X_6010_ net1 _0525_ _2414_ vssd1 vssd1 vccd1 vccd1 _2447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6912_ net110 _0315_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6843_ net41 _0246_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[33\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3986_ _0471_ vssd1 vssd1 vccd1 vccd1 _0472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6774_ net128 _0177_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5725_ _0380_ _0361_ _0389_ _0365_ _2197_ vssd1 vssd1 vccd1 vccd1 _2198_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5656_ _0605_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _2130_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4607_ _1076_ _1080_ _1085_ _1088_ vssd1 vssd1 vccd1 vccd1 _1089_ sky130_fd_sc_hd__and4_1
X_5587_ _3339_ _2998_ vssd1 vssd1 vccd1 vccd1 _2061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4538_ _0541_ _0576_ _0753_ _0580_ _1020_ vssd1 vssd1 vccd1 vccd1 _1021_ sky130_fd_sc_hd__o221a_1
X_4469_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _0952_ sky130_fd_sc_hd__inv_2
X_6208_ _2583_ _2581_ vssd1 vssd1 vccd1 vccd1 _2584_ sky130_fd_sc_hd__and2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ _2536_ vssd1 vssd1 vccd1 vccd1 _0209_ sky130_fd_sc_hd__clkbuf_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3840_ _3061_ _0325_ vssd1 vssd1 vccd1 vccd1 _0326_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3771_ _3072_ _3300_ vssd1 vssd1 vccd1 vccd1 _3305_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5510_ _0498_ _0521_ vssd1 vssd1 vccd1 vccd1 _1985_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6490_ _2798_ _2764_ vssd1 vssd1 vccd1 vccd1 _2826_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5441_ _3188_ _3204_ _1915_ vssd1 vssd1 vccd1 vccd1 _1916_ sky130_fd_sc_hd__o21ai_1
X_5372_ _0614_ _0408_ vssd1 vssd1 vccd1 vccd1 _1848_ sky130_fd_sc_hd__or2_1
X_4323_ _3282_ vssd1 vssd1 vccd1 vccd1 _0807_ sky130_fd_sc_hd__inv_2
X_4254_ _0737_ _0738_ vssd1 vssd1 vccd1 vccd1 _0739_ sky130_fd_sc_hd__nand2_1
X_4185_ _3344_ _3335_ vssd1 vssd1 vccd1 vccd1 _0670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6826_ net180 _0229_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[50\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ egd_top.BitStream_buffer.BS_buffer\[63\] vssd1 vssd1 vccd1 vccd1 _0455_ sky130_fd_sc_hd__clkbuf_4
X_5708_ _3343_ _3016_ vssd1 vssd1 vccd1 vccd1 _2181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6688_ clknet_1_1__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2923_ sky130_fd_sc_hd__buf_1
X_5639_ _2111_ _2112_ vssd1 vssd1 vccd1 vccd1 _2113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6618__109 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__inv_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2918_ clknet_0__2918_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2918_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5990_ _2433_ _2423_ vssd1 vssd1 vccd1 vccd1 _2434_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4941_ _1418_ _1419_ vssd1 vssd1 vccd1 vccd1 _1420_ sky130_fd_sc_hd__nand2_1
X_4872_ _0353_ _0362_ _0356_ _0366_ _1351_ vssd1 vssd1 vccd1 vccd1 _1352_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3823_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _3357_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6542_ _2874_ _2875_ vssd1 vssd1 vccd1 vccd1 _2876_ sky130_fd_sc_hd__nand2_1
X_3754_ _3158_ _3228_ vssd1 vssd1 vccd1 vccd1 _3288_ sky130_fd_sc_hd__nand2_1
X_6473_ _2813_ _2959_ vssd1 vssd1 vccd1 vccd1 _2814_ sky130_fd_sc_hd__nand2_1
X_3685_ _3047_ vssd1 vssd1 vccd1 vccd1 _3219_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5424_ _0764_ _3111_ _1898_ vssd1 vssd1 vccd1 vccd1 _1899_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5355_ _1790_ _1801_ _1814_ _1830_ vssd1 vssd1 vccd1 vccd1 _1831_ sky130_fd_sc_hd__and4_1
X_5286_ _0566_ _0489_ vssd1 vssd1 vccd1 vccd1 _1763_ sky130_fd_sc_hd__nand2_1
X_4306_ _3053_ vssd1 vssd1 vccd1 vccd1 _0790_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4237_ _0699_ _0721_ vssd1 vssd1 vccd1 vccd1 _0722_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4168_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _0653_ sky130_fd_sc_hd__clkbuf_4
X_4099_ _0582_ _0584_ vssd1 vssd1 vccd1 vccd1 _0585_ sky130_fd_sc_hd__or2_1
X_6589__82 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__inv_2
XFILLER_0_92_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6809_ net163 _0212_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[67\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3470_ net4 _3016_ _3007_ vssd1 vssd1 vccd1 vccd1 _3017_ sky130_fd_sc_hd__mux2_1
X_5140_ _1602_ _1617_ vssd1 vssd1 vccd1 vccd1 _1618_ sky130_fd_sc_hd__and2_1
X_5071_ _3192_ _0573_ vssd1 vssd1 vccd1 vccd1 _1549_ sky130_fd_sc_hd__nand2_1
X_4022_ _0507_ vssd1 vssd1 vccd1 vccd1 _0508_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5973_ net4 _0499_ _2415_ vssd1 vssd1 vccd1 vccd1 _2422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4924_ _0606_ _0548_ vssd1 vssd1 vccd1 vccd1 _1404_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4855_ _1081_ _3350_ vssd1 vssd1 vccd1 vccd1 _1335_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3806_ _3339_ vssd1 vssd1 vccd1 vccd1 _3340_ sky130_fd_sc_hd__clkbuf_4
X_4786_ _0551_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _1267_
+ sky130_fd_sc_hd__nand2_1
X_6525_ _2859_ vssd1 vssd1 vccd1 vccd1 _2860_ sky130_fd_sc_hd__inv_2
X_3737_ _3270_ vssd1 vssd1 vccd1 vccd1 _3271_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3668_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _3202_ sky130_fd_sc_hd__inv_2
X_6456_ _2707_ _2013_ vssd1 vssd1 vccd1 vccd1 _2797_ sky130_fd_sc_hd__nand2_1
X_5407_ _0566_ _0493_ vssd1 vssd1 vccd1 vccd1 _1883_ sky130_fd_sc_hd__nand2_1
X_6387_ _2728_ _2729_ vssd1 vssd1 vccd1 vccd1 _2730_ sky130_fd_sc_hd__nand2_1
X_3599_ _3132_ vssd1 vssd1 vccd1 vccd1 _3133_ sky130_fd_sc_hd__clkbuf_4
X_5338_ _1803_ _1808_ _1811_ _1813_ vssd1 vssd1 vccd1 vccd1 _1814_ sky130_fd_sc_hd__and4_1
X_5269_ _0498_ _0535_ vssd1 vssd1 vccd1 vccd1 _1746_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6734__60 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__inv_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4640_ _1105_ _1121_ vssd1 vssd1 vccd1 vccd1 _1122_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4571_ _3206_ _3022_ vssd1 vssd1 vccd1 vccd1 _1053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6310_ _1029_ _1157_ vssd1 vssd1 vccd1 vccd1 _2653_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3522_ _2996_ vssd1 vssd1 vccd1 vccd1 _3056_ sky130_fd_sc_hd__clkbuf_4
X_6241_ _2606_ _2597_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[3\] sky130_fd_sc_hd__xnor2_4
X_3453_ _3002_ net201 vssd1 vssd1 vccd1 vccd1 _3003_ sky130_fd_sc_hd__nand2_1
X_6172_ _2559_ vssd1 vssd1 vccd1 vccd1 _0199_ sky130_fd_sc_hd__clkbuf_1
X_5123_ _0404_ _0379_ _0703_ _0383_ _1600_ vssd1 vssd1 vccd1 vccd1 _1601_ sky130_fd_sc_hd__a221oi_1
X_3384_ net33 net32 vssd1 vssd1 vccd1 vccd1 _2940_ sky130_fd_sc_hd__nor2_1
X_5054_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _1532_ sky130_fd_sc_hd__inv_2
X_4005_ _0490_ vssd1 vssd1 vccd1 vccd1 _0491_ sky130_fd_sc_hd__buf_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5956_ net8 egd_top.BitStream_buffer.BS_buffer\[14\] _2379_ vssd1 vssd1 vccd1 vccd1
+ _2410_ sky130_fd_sc_hd__mux2_1
X_4907_ _1385_ _1386_ vssd1 vssd1 vccd1 vccd1 _1387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5887_ _0565_ _0509_ vssd1 vssd1 vccd1 vccd1 _2359_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4838_ _3271_ _3286_ _3274_ _3290_ vssd1 vssd1 vccd1 vccd1 _1318_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4769_ _0474_ _0521_ vssd1 vssd1 vccd1 vccd1 _1250_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6508_ _2788_ _2843_ vssd1 vssd1 vccd1 vccd1 _2844_ sky130_fd_sc_hd__nor2_1
X_6439_ _2694_ vssd1 vssd1 vccd1 vccd1 _2781_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_7 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6790_ net144 _0193_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[102\]
+ sky130_fd_sc_hd__dfxtp_1
X_5810_ _3253_ _3278_ vssd1 vssd1 vccd1 vccd1 _2282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _0459_ _3069_ vssd1 vssd1 vccd1 vccd1 _2214_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5672_ _2143_ _2144_ vssd1 vssd1 vccd1 vccd1 _2145_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4623_ _1094_ _1098_ _1101_ _1104_ vssd1 vssd1 vccd1 vccd1 _1105_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6713__41 clknet_1_1__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__inv_2
X_4554_ _1034_ _3111_ _1035_ vssd1 vssd1 vccd1 vccd1 _1036_ sky130_fd_sc_hd__o21ai_1
X_3505_ _3043_ vssd1 vssd1 vccd1 vccd1 _0302_ sky130_fd_sc_hd__clkbuf_1
X_4485_ _0352_ _0335_ _0355_ _0323_ vssd1 vssd1 vccd1 vccd1 _0968_ sky130_fd_sc_hd__a22o_1
X_6224_ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3436_ _2988_ _2948_ vssd1 vssd1 vccd1 vccd1 _2990_ sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ net10 _3161_ _2520_ vssd1 vssd1 vccd1 vccd1 _2547_ sky130_fd_sc_hd__mux2_1
X_6086_ _2499_ _2475_ vssd1 vssd1 vccd1 vccd1 _2500_ sky130_fd_sc_hd__and2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5106_ _0780_ _3363_ _1583_ vssd1 vssd1 vccd1 vccd1 _1584_ sky130_fd_sc_hd__o21ai_1
X_5037_ _0756_ _0556_ vssd1 vssd1 vccd1 vccd1 _1516_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5939_ _2398_ _2396_ vssd1 vssd1 vccd1 vccd1 _2399_ sky130_fd_sc_hd__and2_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[2] sky130_fd_sc_hd__buf_12
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[2] sky130_fd_sc_hd__buf_12
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4270_ _0582_ _0576_ _0574_ _0580_ _0754_ vssd1 vssd1 vccd1 vccd1 _0755_ sky130_fd_sc_hd__o221a_1
X_6911_ net109 _0314_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_valid_n
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6842_ net40 _0245_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[34\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _3082_ _0470_ vssd1 vssd1 vccd1 vccd1 _0471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6773_ net127 _0176_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[80\]
+ sky130_fd_sc_hd__dfxtp_1
X_5724_ _0384_ _0368_ _2196_ vssd1 vssd1 vccd1 vccd1 _2197_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5655_ _2099_ _2115_ _2128_ vssd1 vssd1 vccd1 vccd1 _2129_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4606_ _2998_ _3356_ _3010_ _3360_ _1087_ vssd1 vssd1 vccd1 vccd1 _1088_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5586_ _3353_ _3320_ _3357_ _3323_ _2059_ vssd1 vssd1 vccd1 vccd1 _2060_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_25_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4537_ _0742_ _0584_ vssd1 vssd1 vccd1 vccd1 _1020_ sky130_fd_sc_hd__or2_1
X_4468_ _3327_ _3321_ _3341_ _3324_ _0950_ vssd1 vssd1 vccd1 vccd1 _0951_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6207_ net10 _3353_ net197 vssd1 vssd1 vccd1 vccd1 _2583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3419_ _2971_ _2972_ net200 vssd1 vssd1 vccd1 vccd1 _2973_ sky130_fd_sc_hd__and3_2
X_4399_ _0554_ _0545_ _0880_ _0881_ _0882_ vssd1 vssd1 vccd1 vccd1 _0883_ sky130_fd_sc_hd__o2111a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ _2535_ _2529_ vssd1 vssd1 vccd1 vccd1 _2536_ sky130_fd_sc_hd__and2_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _2488_ vssd1 vssd1 vccd1 vccd1 _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3770_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _3304_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5440_ _3206_ _3044_ vssd1 vssd1 vccd1 vccd1 _1915_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5371_ _0403_ _0461_ vssd1 vssd1 vccd1 vccd1 _1847_ sky130_fd_sc_hd__nand2_1
X_4322_ _0803_ _0805_ vssd1 vssd1 vccd1 vccd1 _0806_ sky130_fd_sc_hd__nor2_1
X_4253_ _0534_ _0531_ vssd1 vssd1 vccd1 vccd1 _0738_ sky130_fd_sc_hd__nand2_1
X_4184_ _3340_ _3347_ vssd1 vssd1 vccd1 vccd1 _0669_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6825_ net179 _0228_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[51\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3968_ _0453_ vssd1 vssd1 vccd1 vccd1 _0454_ sky130_fd_sc_hd__clkbuf_4
X_5707_ _3339_ _3010_ vssd1 vssd1 vccd1 vccd1 _2180_ sky130_fd_sc_hd__nand2_1
X_3899_ _2964_ _0325_ vssd1 vssd1 vccd1 vccd1 _0385_ sky130_fd_sc_hd__nand2_1
X_5638_ _0533_ _0339_ vssd1 vssd1 vccd1 vccd1 _2112_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5569_ _3249_ _3282_ vssd1 vssd1 vccd1 vccd1 _2043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2917_ clknet_0__2917_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2917_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4940_ _3160_ _3251_ vssd1 vssd1 vccd1 vccd1 _1419_ sky130_fd_sc_hd__nand2_1
X_4871_ _0966_ _0369_ _1350_ vssd1 vssd1 vccd1 vccd1 _1351_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6610_ clknet_1_1__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2917_ sky130_fd_sc_hd__buf_1
X_3822_ _3355_ vssd1 vssd1 vccd1 vccd1 _3356_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6541_ _2786_ _2755_ _2814_ vssd1 vssd1 vccd1 vccd1 _2875_ sky130_fd_sc_hd__nor3_1
X_6679__9 clknet_1_1__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__inv_2
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _3286_ vssd1 vssd1 vccd1 vccd1 _3287_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6472_ _2800_ _2810_ vssd1 vssd1 vccd1 vccd1 _2813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3684_ _3217_ vssd1 vssd1 vccd1 vccd1 _3218_ sky130_fd_sc_hd__clkbuf_4
X_5423_ _3114_ _3161_ vssd1 vssd1 vccd1 vccd1 _1898_ sky130_fd_sc_hd__nand2_1
X_5354_ _1818_ _1822_ _1826_ _1829_ vssd1 vssd1 vccd1 vccd1 _1830_ sky130_fd_sc_hd__and4_1
X_4305_ _3019_ _3198_ _3022_ _3201_ _0788_ vssd1 vssd1 vccd1 vccd1 _0789_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6683__13 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__inv_2
X_5285_ _0563_ _0499_ vssd1 vssd1 vccd1 vccd1 _1762_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4236_ _0707_ _0713_ _0717_ _0720_ vssd1 vssd1 vccd1 vccd1 _0721_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _3266_ _3264_ _0651_ _3268_ vssd1 vssd1 vccd1 vccd1 _0652_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4098_ _0583_ vssd1 vssd1 vccd1 vccd1 _0584_ sky130_fd_sc_hd__buf_2
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6808_ net162 _0211_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[68\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6624__114 clknet_1_0__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__inv_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5070_ _3050_ _3170_ _3053_ _3173_ _1547_ vssd1 vssd1 vccd1 vccd1 _1548_ sky130_fd_sc_hd__a221oi_1
X_4021_ _3131_ _0470_ vssd1 vssd1 vccd1 vccd1 _0507_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5972_ _2421_ vssd1 vssd1 vccd1 vccd1 _0261_ sky130_fd_sc_hd__clkbuf_1
X_4923_ _1372_ _1389_ _1402_ vssd1 vssd1 vccd1 vccd1 _1403_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4854_ _3344_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1334_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _3126_ _3300_ vssd1 vssd1 vccd1 vccd1 _3339_ sky130_fd_sc_hd__and2_1
X_4785_ _0547_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1266_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3736_ _3131_ _3228_ vssd1 vssd1 vccd1 vccd1 _3270_ sky130_fd_sc_hd__and2_1
X_6524_ _2707_ _1774_ _1530_ vssd1 vssd1 vccd1 vccd1 _2859_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_27_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6455_ _2709_ _2764_ _2726_ vssd1 vssd1 vccd1 vccd1 _2796_ sky130_fd_sc_hd__nand3_1
X_3667_ _3200_ vssd1 vssd1 vccd1 vccd1 _3201_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6386_ _2701_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] _2668_ vssd1
+ vssd1 vccd1 vccd1 _2729_ sky130_fd_sc_hd__nand3_1
X_3598_ _3131_ _3065_ vssd1 vssd1 vccd1 vccd1 _3132_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5406_ _0563_ _0513_ vssd1 vssd1 vccd1 vccd1 _1882_ sky130_fd_sc_hd__nand2_1
X_5337_ _3314_ _3281_ _3310_ _3285_ _1812_ vssd1 vssd1 vccd1 vccd1 _1813_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_2_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5268_ _1741_ _0472_ _1742_ _1744_ vssd1 vssd1 vccd1 vccd1 _1745_ sky130_fd_sc_hd__o211a_1
X_6647__136 clknet_1_1__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__inv_2
X_4219_ _0403_ _0703_ vssd1 vssd1 vccd1 vccd1 _0704_ sky130_fd_sc_hd__nand2_1
X_5199_ _3040_ _3198_ _3044_ _3201_ _1675_ vssd1 vssd1 vccd1 vccd1 _1676_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2919_ _2919_ vssd1 vssd1 vccd1 vccd1 clknet_0__2919_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _3044_ _3184_ _3047_ _3187_ _1051_ vssd1 vssd1 vccd1 vccd1 _1052_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3521_ _3055_ vssd1 vssd1 vccd1 vccd1 _0298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3452_ _2999_ _3000_ _2945_ _3001_ vssd1 vssd1 vccd1 vccd1 _3002_ sky130_fd_sc_hd__a22o_4
X_6240_ _2598_ _2599_ vssd1 vssd1 vccd1 vccd1 _2606_ sky130_fd_sc_hd__nand2_2
X_6171_ _2558_ _2554_ vssd1 vssd1 vccd1 vccd1 _2559_ sky130_fd_sc_hd__and2_1
X_3383_ net31 vssd1 vssd1 vccd1 vccd1 _2939_ sky130_fd_sc_hd__inv_2
X_5122_ _0406_ _0386_ _1599_ vssd1 vssd1 vccd1 vccd1 _1600_ sky130_fd_sc_hd__o21ai_1
X_5053_ _3056_ _1529_ _1531_ vssd1 vssd1 vccd1 vccd1 _0290_ sky130_fd_sc_hd__o21a_1
X_4004_ _3112_ _0470_ vssd1 vssd1 vccd1 vccd1 _0490_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5955_ _2409_ vssd1 vssd1 vccd1 vccd1 _0266_ sky130_fd_sc_hd__clkbuf_1
X_4906_ _0534_ _0689_ vssd1 vssd1 vccd1 vccd1 _1386_ sky130_fd_sc_hd__nand2_1
X_5886_ _0562_ _0467_ vssd1 vssd1 vccd1 vccd1 _2358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4837_ _0642_ _3264_ _0794_ _3268_ vssd1 vssd1 vccd1 vccd1 _1317_ sky130_fd_sc_hd__o22ai_1
X_4768_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _1249_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4699_ _3206_ _3025_ vssd1 vssd1 vccd1 vccd1 _1180_ sky130_fd_sc_hd__nand2_1
X_6507_ _2840_ _2814_ vssd1 vssd1 vccd1 vccd1 _2843_ sky130_fd_sc_hd__nand2_1
X_3719_ _3109_ _3228_ vssd1 vssd1 vccd1 vccd1 _3253_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6438_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2745_ vssd1 vssd1 vccd1
+ vccd1 _2780_ sky130_fd_sc_hd__nor2_1
X_6369_ _2699_ _2705_ _2711_ vssd1 vssd1 vccd1 vccd1 _2712_ sky130_fd_sc_hd__nand3_2
XFILLER_0_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 net4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5740_ _0455_ _0431_ _3107_ _0435_ _2212_ vssd1 vssd1 vccd1 vccd1 _2213_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5671_ _3159_ _0804_ vssd1 vssd1 vccd1 vccd1 _2144_ sky130_fd_sc_hd__nand2_1
X_4622_ _0437_ _0379_ _0443_ _0383_ _1103_ vssd1 vssd1 vccd1 vccd1 _1104_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4553_ _3114_ _3136_ vssd1 vssd1 vccd1 vccd1 _1035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4484_ _0833_ _0345_ _0966_ _0349_ vssd1 vssd1 vccd1 vccd1 _0967_ sky130_fd_sc_hd__o22ai_1
X_3504_ _3041_ _3042_ vssd1 vssd1 vccd1 vccd1 _3043_ sky130_fd_sc_hd__and2_1
X_3435_ _2932_ vssd1 vssd1 vccd1 vccd1 _2989_ sky130_fd_sc_hd__clkbuf_4
X_6223_ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ vssd1 vssd1 vccd1 vccd1 _2595_ sky130_fd_sc_hd__or2_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _2546_ vssd1 vssd1 vccd1 vccd1 _0204_ sky130_fd_sc_hd__clkbuf_1
X_6085_ net16 _0400_ _2486_ vssd1 vssd1 vccd1 vccd1 _2499_ sky130_fd_sc_hd__mux2_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _3365_ _3025_ vssd1 vssd1 vccd1 vccd1 _1583_ sky130_fd_sc_hd__nand2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5036_ _0551_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1515_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5938_ net14 egd_top.BitStream_buffer.BS_buffer\[8\] _2380_ vssd1 vssd1 vccd1 vccd1
+ _2398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5869_ _0685_ _0471_ _2338_ _2340_ vssd1 vssd1 vccd1 vccd1 _2341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 la_data_out_30_27[3] sky130_fd_sc_hd__buf_12
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[3] sky130_fd_sc_hd__buf_12
XFILLER_0_85_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6910_ net108 _0313_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[112\]
+ sky130_fd_sc_hd__dfxtp_1
X_6841_ net195 _0244_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[35\]
+ sky130_fd_sc_hd__dfxtp_1
X_3984_ _0469_ vssd1 vssd1 vccd1 vccd1 _0470_ sky130_fd_sc_hd__buf_2
X_6772_ net126 _0175_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[81\]
+ sky130_fd_sc_hd__dfxtp_1
X_5723_ _0370_ _0437_ vssd1 vssd1 vccd1 vccd1 _2196_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5654_ _2119_ _2123_ _2125_ _2127_ vssd1 vssd1 vccd1 vccd1 _2128_ sky130_fd_sc_hd__and4_1
XFILLER_0_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4605_ _0922_ _3363_ _1086_ vssd1 vssd1 vccd1 vccd1 _1087_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5585_ _2057_ _2058_ vssd1 vssd1 vccd1 vccd1 _2059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4536_ _0756_ _0561_ _1016_ _1017_ _1018_ vssd1 vssd1 vccd1 vccd1 _1019_ sky130_fd_sc_hd__o2111a_1
X_4467_ _0948_ _0949_ vssd1 vssd1 vccd1 vccd1 _0950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6206_ _2582_ vssd1 vssd1 vccd1 vccd1 _0188_ sky130_fd_sc_hd__clkbuf_1
X_3418_ net196 vssd1 vssd1 vccd1 vccd1 _2972_ sky130_fd_sc_hd__inv_2
X_4398_ _0568_ _0556_ vssd1 vssd1 vccd1 vccd1 _0882_ sky130_fd_sc_hd__or2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6137_ net16 _3134_ _2521_ vssd1 vssd1 vccd1 vccd1 _2535_ sky130_fd_sc_hd__mux2_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _2487_ _2475_ vssd1 vssd1 vccd1 vccd1 _2488_ sky130_fd_sc_hd__and2_1
X_5019_ _0474_ _0359_ vssd1 vssd1 vccd1 vccd1 _1498_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5370_ _0399_ _3107_ vssd1 vssd1 vccd1 vccd1 _1846_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4321_ _3271_ _0653_ _3274_ _0804_ vssd1 vssd1 vccd1 vccd1 _0805_ sky130_fd_sc_hd__a22o_1
X_4252_ _0530_ _0521_ vssd1 vssd1 vccd1 vccd1 _0737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4183_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _0668_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6824_ net178 _0227_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[52\]
+ sky130_fd_sc_hd__dfxtp_1
X_6604__96 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__inv_2
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3967_ _0452_ vssd1 vssd1 vccd1 vccd1 _0453_ sky130_fd_sc_hd__buf_1
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5706_ _3357_ _3320_ _0674_ _3323_ _2178_ vssd1 vssd1 vccd1 vccd1 _2179_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3898_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _0384_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5637_ _0529_ _0335_ vssd1 vssd1 vccd1 vccd1 _2111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5568_ _3245_ _3290_ vssd1 vssd1 vccd1 vccd1 _2042_ sky130_fd_sc_hd__nand2_1
X_4519_ _0499_ _0488_ _0513_ _0492_ _1001_ vssd1 vssd1 vccd1 vccd1 _1002_ sky130_fd_sc_hd__a221oi_1
X_5499_ _0412_ _0440_ _1973_ vssd1 vssd1 vccd1 vccd1 _1974_ sky130_fd_sc_hd__o21ai_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2916_ clknet_0__2916_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2916_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _0371_ _0335_ vssd1 vssd1 vccd1 vccd1 _1350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3821_ _3354_ vssd1 vssd1 vccd1 vccd1 _3355_ sky130_fd_sc_hd__buf_1
X_6540_ _2873_ vssd1 vssd1 vccd1 vccd1 _2874_ sky130_fd_sc_hd__inv_2
X_3752_ egd_top.BitStream_buffer.BS_buffer\[92\] vssd1 vssd1 vccd1 vccd1 _3286_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6471_ _2791_ _2811_ vssd1 vssd1 vccd1 vccd1 _2812_ sky130_fd_sc_hd__nand2_1
X_3683_ _3158_ _3167_ vssd1 vssd1 vccd1 vccd1 _3217_ sky130_fd_sc_hd__nand2_1
X_5422_ _3265_ _3068_ _3272_ _3075_ _1896_ vssd1 vssd1 vccd1 vccd1 _1897_ sky130_fd_sc_hd__a221oi_1
X_5353_ _3025_ _3356_ _3028_ _3360_ _1828_ vssd1 vssd1 vccd1 vccd1 _1829_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4304_ _0786_ _3204_ _0787_ vssd1 vssd1 vccd1 vccd1 _0788_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5284_ _0756_ _0545_ _1758_ _1759_ _1760_ vssd1 vssd1 vccd1 vccd1 _1761_ sky130_fd_sc_hd__o2111a_1
X_4235_ _0451_ _0450_ _0461_ _0454_ _0719_ vssd1 vssd1 vccd1 vccd1 _0720_ sky130_fd_sc_hd__a221oi_1
X_4166_ egd_top.BitStream_buffer.BS_buffer\[86\] vssd1 vssd1 vccd1 vccd1 _0651_ sky130_fd_sc_hd__inv_2
X_4097_ _3103_ _0542_ vssd1 vssd1 vccd1 vccd1 _0583_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6807_ net161 _0210_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[69\]
+ sky130_fd_sc_hd__dfxtp_1
X_4999_ _0700_ _0386_ _1477_ vssd1 vssd1 vccd1 vccd1 _1478_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670__157 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__inv_2
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _0505_ vssd1 vssd1 vccd1 vccd1 _0506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5971_ _2420_ _2396_ vssd1 vssd1 vccd1 vccd1 _2421_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4922_ _1393_ _1397_ _1399_ _1401_ vssd1 vssd1 vccd1 vccd1 _1402_ sky130_fd_sc_hd__and4_1
XFILLER_0_74_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4853_ _3340_ _3297_ vssd1 vssd1 vccd1 vccd1 _1333_ sky130_fd_sc_hd__nand2_1
X_4784_ _1253_ _1256_ _1260_ _1264_ vssd1 vssd1 vccd1 vccd1 _1265_ sky130_fd_sc_hd__and4_1
X_3804_ _3337_ vssd1 vssd1 vccd1 vccd1 _3338_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6523_ _2857_ _2792_ _2829_ vssd1 vssd1 vccd1 vccd1 _2858_ sky130_fd_sc_hd__nand3_1
X_3735_ _3262_ _3264_ _3266_ _3268_ vssd1 vssd1 vccd1 vccd1 _3269_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6454_ _2792_ _2794_ _2764_ vssd1 vssd1 vccd1 vccd1 _2795_ sky130_fd_sc_hd__nand3_1
X_3666_ _3199_ vssd1 vssd1 vccd1 vccd1 _3200_ sky130_fd_sc_hd__buf_1
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5405_ _0890_ _0545_ _1878_ _1879_ _1880_ vssd1 vssd1 vccd1 vccd1 _1881_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6385_ _2669_ _2700_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1
+ vssd1 vccd1 vccd1 _2728_ sky130_fd_sc_hd__o21ai_1
X_3597_ _3059_ egd_top.BitStream_buffer.pc\[2\] _3096_ vssd1 vssd1 vccd1 vccd1 _3131_
+ sky130_fd_sc_hd__and3_4
X_5336_ _0671_ _3289_ _3336_ _3293_ vssd1 vssd1 vccd1 vccd1 _1812_ sky130_fd_sc_hd__o22ai_1
X_5267_ _1743_ vssd1 vssd1 vccd1 vccd1 _1744_ sky130_fd_sc_hd__inv_2
X_4218_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _0703_ sky130_fd_sc_hd__clkbuf_4
X_5198_ _1047_ _3204_ _1674_ vssd1 vssd1 vccd1 vccd1 _1675_ sky130_fd_sc_hd__o21ai_1
X_4149_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _0634_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2918_ _2918_ vssd1 vssd1 vccd1 vccd1 clknet_0__2918_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3520_ _3054_ _3042_ vssd1 vssd1 vccd1 vccd1 _3055_ sky130_fd_sc_hd__and2_1
X_3451_ _2940_ _2930_ vssd1 vssd1 vccd1 vccd1 _3001_ sky130_fd_sc_hd__nand2_1
X_6170_ net7 _3318_ _2557_ vssd1 vssd1 vccd1 vccd1 _2558_ sky130_fd_sc_hd__mux2_1
X_3382_ _2935_ _2936_ _2938_ vssd1 vssd1 vccd1 vccd1 _0320_ sky130_fd_sc_hd__a21oi_1
X_5121_ _0388_ _0400_ vssd1 vssd1 vccd1 vccd1 _1599_ sky130_fd_sc_hd__nand2_1
X_5052_ _1530_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1531_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4003_ egd_top.BitStream_buffer.BS_buffer\[17\] vssd1 vssd1 vccd1 vccd1 _0489_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5954_ _2408_ _2396_ vssd1 vssd1 vccd1 vccd1 _2409_ sky130_fd_sc_hd__and2_1
X_4905_ _0530_ _0372_ vssd1 vssd1 vccd1 vccd1 _1385_ sky130_fd_sc_hd__nand2_1
X_5885_ _0728_ _0544_ _2354_ _2355_ _2356_ vssd1 vssd1 vccd1 vccd1 _2357_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_47_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4836_ _1312_ _1313_ _1314_ _1315_ vssd1 vssd1 vccd1 vccd1 _1316_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6653__141 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__inv_2
X_4767_ _1232_ _1247_ vssd1 vssd1 vccd1 vccd1 _1248_ sky130_fd_sc_hd__and2_1
X_6506_ _2840_ _2841_ vssd1 vssd1 vccd1 vccd1 _2842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3718_ _3250_ _3251_ vssd1 vssd1 vccd1 vccd1 _3252_ sky130_fd_sc_hd__nand2_1
X_4698_ _3047_ _3184_ _3050_ _3187_ _1178_ vssd1 vssd1 vccd1 vccd1 _1179_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6437_ _1406_ _2744_ vssd1 vssd1 vccd1 vccd1 _2779_ sky130_fd_sc_hd__nor2_1
X_3649_ _3182_ vssd1 vssd1 vccd1 vccd1 _3183_ sky130_fd_sc_hd__buf_1
X_6368_ _2709_ _2710_ vssd1 vssd1 vccd1 vccd1 _2711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5319_ _0573_ _3184_ _0581_ _3187_ _1794_ vssd1 vssd1 vccd1 vccd1 _1795_ sky130_fd_sc_hd__a221oi_1
X_6299_ _2643_ vssd1 vssd1 vccd1 vccd1 _0162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5670_ _3154_ _3225_ vssd1 vssd1 vccd1 vccd1 _2143_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4621_ _0986_ _0386_ _1102_ vssd1 vssd1 vccd1 vccd1 _1103_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4552_ _3129_ vssd1 vssd1 vccd1 vccd1 _1034_ sky130_fd_sc_hd__inv_2
X_4483_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0966_ sky130_fd_sc_hd__inv_2
X_3503_ _2932_ vssd1 vssd1 vccd1 vccd1 _3042_ sky130_fd_sc_hd__buf_2
XFILLER_0_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6222_ _2960_ _2593_ _2592_ vssd1 vssd1 vccd1 vccd1 _2594_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3434_ _2986_ _2987_ vssd1 vssd1 vccd1 vccd1 _2988_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6153_ _2545_ _2529_ vssd1 vssd1 vccd1 vccd1 _2546_ sky130_fd_sc_hd__and2_1
X_6084_ _2498_ vssd1 vssd1 vccd1 vccd1 _0226_ sky130_fd_sc_hd__clkbuf_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _3361_ _3338_ _1579_ _1580_ _1581_ vssd1 vssd1 vccd1 vccd1 _1582_ sky130_fd_sc_hd__o2111a_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _0547_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1514_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5937_ _2397_ vssd1 vssd1 vccd1 vccd1 _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _2339_ vssd1 vssd1 vccd1 vccd1 _2340_ sky130_fd_sc_hd__inv_2
X_4819_ _1174_ _3176_ _3188_ _3179_ vssd1 vssd1 vccd1 vccd1 _1299_ sky130_fd_sc_hd__o22ai_1
X_5799_ _0548_ _3183_ egd_top.BitStream_buffer.BS_buffer\[7\] _3186_ _2270_ vssd1
+ vssd1 vccd1 vccd1 _2271_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6704__32 clknet_1_1__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__inv_2
XFILLER_0_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[4] sky130_fd_sc_hd__buf_12
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6753__1 clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__inv_2
X_6840_ net194 _0243_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[36\]
+ sky130_fd_sc_hd__dfxtp_1
X_6771_ net125 _0174_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[82\]
+ sky130_fd_sc_hd__dfxtp_1
X_5722_ _2193_ _2194_ vssd1 vssd1 vccd1 vccd1 _2195_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3983_ _2965_ _3063_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _0469_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5653_ _0479_ _0588_ _0482_ _0591_ _2126_ vssd1 vssd1 vccd1 vccd1 _2127_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4604_ _3365_ _3013_ vssd1 vssd1 vccd1 vccd1 _1086_ sky130_fd_sc_hd__nand2_1
X_5584_ _3329_ _0674_ vssd1 vssd1 vccd1 vccd1 _2058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4535_ _0593_ _0570_ vssd1 vssd1 vccd1 vccd1 _1018_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4466_ _3330_ _3347_ vssd1 vssd1 vccd1 vccd1 _0949_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6205_ _2580_ _2581_ vssd1 vssd1 vccd1 vccd1 _2582_ sky130_fd_sc_hd__and2_1
X_3417_ net198 vssd1 vssd1 vccd1 vccd1 _2971_ sky130_fd_sc_hd__inv_2
X_4397_ _0551_ _0548_ vssd1 vssd1 vccd1 vccd1 _0881_ sky130_fd_sc_hd__nand2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ _2534_ vssd1 vssd1 vccd1 vccd1 _0210_ sky130_fd_sc_hd__clkbuf_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ net7 _0437_ _2486_ vssd1 vssd1 vccd1 vccd1 _2487_ sky130_fd_sc_hd__mux2_1
X_5018_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _1497_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4320_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _0804_ sky130_fd_sc_hd__buf_4
X_4251_ _0468_ _0506_ _0732_ _0733_ _0735_ vssd1 vssd1 vccd1 vccd1 _0736_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_10_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4182_ _3322_ _3321_ _3331_ _3324_ _0666_ vssd1 vssd1 vccd1 vccd1 _0667_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6823_ net177 _0226_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[53\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3966_ _3153_ _2966_ vssd1 vssd1 vccd1 vccd1 _0452_ sky130_fd_sc_hd__and2_1
X_5705_ _2176_ _2177_ vssd1 vssd1 vccd1 vccd1 _2178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5636_ _0690_ _0505_ _2107_ _2108_ _2109_ vssd1 vssd1 vccd1 vccd1 _2110_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3897_ _0382_ vssd1 vssd1 vccd1 vccd1 _0383_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5567_ _3345_ _3230_ _3335_ _3234_ _2040_ vssd1 vssd1 vccd1 vccd1 _2041_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_79_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5498_ _0442_ _0447_ vssd1 vssd1 vccd1 vccd1 _1973_ sky130_fd_sc_hd__nand2_1
X_4518_ _0516_ _0496_ _1000_ vssd1 vssd1 vccd1 vccd1 _1001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4449_ _3246_ _0646_ vssd1 vssd1 vccd1 vccd1 _0932_ sky130_fd_sc_hd__nand2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _2522_ _2502_ vssd1 vssd1 vccd1 vccd1 _2523_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__2915_ clknet_0__2915_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2915_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3158_ _3299_ vssd1 vssd1 vccd1 vccd1 _3354_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3751_ _3284_ vssd1 vssd1 vccd1 vccd1 _3285_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6470_ _2800_ _2810_ _2716_ vssd1 vssd1 vccd1 vccd1 _2811_ sky130_fd_sc_hd__a21oi_1
X_3682_ _3044_ vssd1 vssd1 vccd1 vccd1 _3216_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5421_ _1776_ _3084_ _3262_ _3092_ vssd1 vssd1 vccd1 vccd1 _1896_ sky130_fd_sc_hd__o22ai_1
X_5352_ _1047_ _3363_ _1827_ vssd1 vssd1 vccd1 vccd1 _1828_ sky130_fd_sc_hd__o21ai_1
X_4303_ _3206_ _3016_ vssd1 vssd1 vccd1 vccd1 _0787_ sky130_fd_sc_hd__nand2_1
X_5283_ _1022_ _0556_ vssd1 vssd1 vccd1 vccd1 _1760_ sky130_fd_sc_hd__or2_1
X_4234_ _3108_ _0458_ _0718_ vssd1 vssd1 vccd1 vccd1 _0719_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _0645_ _0647_ _0648_ _0649_ vssd1 vssd1 vccd1 vccd1 _0650_ sky130_fd_sc_hd__and4_1
X_4096_ _0581_ vssd1 vssd1 vccd1 vccd1 _0582_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6806_ net160 _0209_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[70\]
+ sky130_fd_sc_hd__dfxtp_1
X_4998_ _0388_ _0703_ vssd1 vssd1 vccd1 vccd1 _1477_ sky130_fd_sc_hd__nand2_1
X_3949_ _0434_ vssd1 vssd1 vccd1 vccd1 _0435_ sky130_fd_sc_hd__buf_1
X_6746__71 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__inv_2
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5619_ _0708_ _0439_ _2092_ vssd1 vssd1 vccd1 vccd1 _2093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6595__88 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__inv_2
XFILLER_0_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5970_ net5 _0493_ _2415_ vssd1 vssd1 vccd1 vccd1 _2420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4921_ _0513_ _0589_ _0515_ _0592_ _1400_ vssd1 vssd1 vccd1 vccd1 _1401_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4852_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _1332_ sky130_fd_sc_hd__inv_2
X_3803_ _3122_ _3300_ vssd1 vssd1 vccd1 vccd1 _3337_ sky130_fd_sc_hd__nand2_1
X_4783_ _0372_ _0524_ _0691_ _0528_ _1263_ vssd1 vssd1 vccd1 vccd1 _1264_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6522_ _2768_ _2794_ vssd1 vssd1 vccd1 vccd1 _2857_ sky130_fd_sc_hd__nor2_1
X_3734_ _3267_ vssd1 vssd1 vccd1 vccd1 _3268_ sky130_fd_sc_hd__clkbuf_4
X_6453_ _1774_ _2707_ _2793_ vssd1 vssd1 vccd1 vccd1 _2794_ sky130_fd_sc_hd__o21ai_1
X_3665_ _3103_ _3167_ vssd1 vssd1 vccd1 vccd1 _3199_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5404_ _1150_ _0556_ vssd1 vssd1 vccd1 vccd1 _1880_ sky130_fd_sc_hd__or2_1
X_6384_ _2723_ _2726_ vssd1 vssd1 vccd1 vccd1 _2727_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3596_ _3128_ _3129_ vssd1 vssd1 vccd1 vccd1 _3130_ sky130_fd_sc_hd__nand2_1
X_5335_ _1809_ _1810_ vssd1 vssd1 vccd1 vccd1 _1811_ sky130_fd_sc_hd__nor2_1
X_5266_ _0478_ _0372_ _0481_ _0691_ vssd1 vssd1 vccd1 vccd1 _1743_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4217_ _0399_ _0701_ vssd1 vssd1 vccd1 vccd1 _0702_ sky130_fd_sc_hd__nand2_1
X_5197_ _3206_ _3037_ vssd1 vssd1 vccd1 vccd1 _1674_ sky130_fd_sc_hd__nand2_1
X_4148_ _3034_ _3184_ _3037_ _3187_ _0632_ vssd1 vssd1 vccd1 vccd1 _0633_ sky130_fd_sc_hd__a221oi_1
X_4079_ _3082_ _0543_ vssd1 vssd1 vccd1 vccd1 _0565_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0__2917_ _2917_ vssd1 vssd1 vccd1 vccd1 clknet_0__2917_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6630__120 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__inv_2
XFILLER_0_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6725__52 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__inv_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3450_ net30 net29 vssd1 vssd1 vccd1 vccd1 _3000_ sky130_fd_sc_hd__nand2_1
X_3381_ _2937_ vssd1 vssd1 vccd1 vccd1 _2938_ sky130_fd_sc_hd__clkbuf_4
X_5120_ _0339_ _0362_ _0335_ _0366_ _1597_ vssd1 vssd1 vccd1 vccd1 _1598_ sky130_fd_sc_hd__a221oi_1
X_5051_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] vssd1 vssd1 vccd1 vccd1
+ _1530_ sky130_fd_sc_hd__inv_2
X_4002_ _0487_ vssd1 vssd1 vccd1 vccd1 _0488_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5953_ net9 egd_top.BitStream_buffer.BS_buffer\[13\] _2379_ vssd1 vssd1 vccd1 vccd1
+ _2408_ sky130_fd_sc_hd__mux2_1
X_4904_ _1249_ _0506_ _1381_ _1382_ _1383_ vssd1 vssd1 vccd1 vccd1 _1384_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5884_ _0516_ _0555_ vssd1 vssd1 vccd1 vccd1 _2356_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4835_ _3258_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _1315_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _1236_ _1240_ _1243_ _1246_ vssd1 vssd1 vccd1 vccd1 _1247_ sky130_fd_sc_hd__and4_1
X_6505_ _2788_ _2811_ vssd1 vssd1 vccd1 vccd1 _2841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3717_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _3251_ sky130_fd_sc_hd__buf_4
XFILLER_0_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4697_ _0926_ _3190_ _1177_ vssd1 vssd1 vccd1 vccd1 _1178_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6436_ _2654_ _2777_ vssd1 vssd1 vccd1 vccd1 _2778_ sky130_fd_sc_hd__nor2_1
X_3648_ _3082_ _3166_ vssd1 vssd1 vccd1 vccd1 _3182_ sky130_fd_sc_hd__and2_1
X_6367_ _2685_ _2669_ vssd1 vssd1 vccd1 vccd1 _2710_ sky130_fd_sc_hd__nor2_2
X_3579_ _3112_ _3065_ vssd1 vssd1 vccd1 vccd1 _3113_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5318_ _0541_ _3190_ _1793_ vssd1 vssd1 vccd1 vccd1 _1794_ sky130_fd_sc_hd__o21ai_1
X_6298_ _2642_ _2372_ vssd1 vssd1 vccd1 vccd1 _2643_ sky130_fd_sc_hd__and2_1
X_5249_ _0403_ _0451_ vssd1 vssd1 vccd1 vccd1 _1726_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4620_ _0388_ _0429_ vssd1 vssd1 vccd1 vccd1 _1102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6637__126 clknet_1_0__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__inv_2
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4551_ _3144_ _3068_ _3149_ _3075_ _1032_ vssd1 vssd1 vccd1 vccd1 _1033_ sky130_fd_sc_hd__a221oi_1
X_4482_ _0380_ _0328_ _0389_ _0332_ _0964_ vssd1 vssd1 vccd1 vccd1 _0965_ sky130_fd_sc_hd__a221oi_1
X_3502_ net11 _3040_ _3006_ vssd1 vssd1 vccd1 vccd1 _3041_ sky130_fd_sc_hd__mux2_1
X_6221_ _2591_ _2592_ vssd1 vssd1 vccd1 vccd1 _2593_ sky130_fd_sc_hd__nand2_2
X_3433_ _2928_ _2939_ net34 net32 vssd1 vssd1 vccd1 vccd1 _2987_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ net11 _3069_ _2521_ vssd1 vssd1 vccd1 vccd1 _2545_ sky130_fd_sc_hd__mux2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _1332_ _3350_ vssd1 vssd1 vccd1 vccd1 _1581_ sky130_fd_sc_hd__or2_1
X_6083_ _2497_ _2475_ vssd1 vssd1 vccd1 vccd1 _2498_ sky130_fd_sc_hd__and2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _1501_ _1504_ _1508_ _1512_ vssd1 vssd1 vccd1 vccd1 _1513_ sky130_fd_sc_hd__and4_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5936_ _2395_ _2396_ vssd1 vssd1 vccd1 vccd1 _2397_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5867_ _0477_ egd_top.BitStream_buffer.BS_buffer\[40\] _0480_ egd_top.BitStream_buffer.BS_buffer\[41\]
+ vssd1 vssd1 vccd1 vccd1 _2339_ sky130_fd_sc_hd__a22o_1
X_4818_ _1286_ _1289_ _1293_ _1297_ vssd1 vssd1 vccd1 vccd1 _1298_ sky130_fd_sc_hd__and4_1
X_5798_ _0568_ _3189_ _2269_ vssd1 vssd1 vccd1 vccd1 _2270_ sky130_fd_sc_hd__o21ai_1
X_4749_ _1114_ _0386_ _1229_ vssd1 vssd1 vccd1 vccd1 _1230_ sky130_fd_sc_hd__o21ai_1
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[5] sky130_fd_sc_hd__buf_12
X_6419_ _2709_ _2726_ vssd1 vssd1 vccd1 vccd1 _2761_ sky130_fd_sc_hd__nand2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3982_ _0467_ vssd1 vssd1 vccd1 vccd1 _0468_ sky130_fd_sc_hd__inv_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6770_ net124 _0173_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[83\]
+ sky130_fd_sc_hd__dfxtp_1
X_5721_ _0351_ egd_top.BitStream_buffer.BS_buffer\[51\] _0354_ egd_top.BitStream_buffer.BS_buffer\[52\]
+ vssd1 vssd1 vccd1 vccd1 _2194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5652_ _0468_ _0594_ _0723_ _0597_ vssd1 vssd1 vccd1 vccd1 _2126_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603_ _1081_ _3338_ _1082_ _1083_ _1084_ vssd1 vssd1 vccd1 vccd1 _1085_ sky130_fd_sc_hd__o2111a_1
X_5583_ _3325_ _0675_ vssd1 vssd1 vccd1 vccd1 _2057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4534_ _0566_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _1017_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4465_ _3326_ _3345_ vssd1 vssd1 vccd1 vccd1 _0948_ sky130_fd_sc_hd__nand2_1
X_3416_ net30 _2969_ vssd1 vssd1 vccd1 vccd1 _2970_ sky130_fd_sc_hd__nor2_1
X_6204_ _2932_ vssd1 vssd1 vccd1 vccd1 _2581_ sky130_fd_sc_hd__clkbuf_4
X_4396_ _0547_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0880_
+ sky130_fd_sc_hd__nand2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6135_ _2533_ _2529_ vssd1 vssd1 vccd1 vccd1 _2534_ sky130_fd_sc_hd__and2_1
X_6066_ _2485_ vssd1 vssd1 vccd1 vccd1 _2486_ sky130_fd_sc_hd__buf_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5017_ _1480_ _1495_ vssd1 vssd1 vccd1 vccd1 _1496_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6899_ net97 _0302_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[123\]
+ sky130_fd_sc_hd__dfxtp_1
X_5919_ net5 _0573_ _2380_ vssd1 vssd1 vccd1 vccd1 _2385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6695__24 clknet_1_1__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__inv_2
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4250_ _0734_ _0518_ vssd1 vssd1 vccd1 vccd1 _0735_ sky130_fd_sc_hd__or2_1
X_4181_ _0664_ _0665_ vssd1 vssd1 vccd1 vccd1 _0666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6822_ net176 _0225_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[54\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3965_ egd_top.BitStream_buffer.BS_buffer\[61\] vssd1 vssd1 vccd1 vccd1 _0451_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3896_ _0381_ vssd1 vssd1 vccd1 vccd1 _0382_ sky130_fd_sc_hd__buf_1
XFILLER_0_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5704_ _3329_ _0675_ vssd1 vssd1 vccd1 vccd1 _2177_ sky130_fd_sc_hd__nand2_1
X_5635_ _1741_ _0517_ vssd1 vssd1 vccd1 vccd1 _2109_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5566_ _1444_ _3237_ _3348_ _3240_ vssd1 vssd1 vccd1 vccd1 _2040_ sky130_fd_sc_hd__o22ai_1
X_4517_ _0498_ _0509_ vssd1 vssd1 vccd1 vccd1 _1000_ sky130_fd_sc_hd__nand2_1
X_5497_ _0620_ _0414_ _1969_ _1970_ _1971_ vssd1 vssd1 vccd1 vccd1 _1972_ sky130_fd_sc_hd__o2111a_1
X_4448_ _3290_ _3231_ _3278_ _3235_ _0930_ vssd1 vssd1 vccd1 vccd1 _0931_ sky130_fd_sc_hd__a221oi_1
X_4379_ _0474_ _0482_ vssd1 vssd1 vccd1 vccd1 _0863_ sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ net7 _3107_ _2521_ vssd1 vssd1 vccd1 vccd1 _2522_ sky130_fd_sc_hd__mux2_1
X_6049_ net11 _0329_ _2451_ vssd1 vssd1 vccd1 vccd1 _2474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2914_ clknet_0__2914_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2914_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3750_ _3283_ vssd1 vssd1 vccd1 vccd1 _3284_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3681_ _3214_ vssd1 vssd1 vccd1 vccd1 _3215_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5420_ _3056_ _1893_ _1895_ vssd1 vssd1 vccd1 vccd1 _0287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5351_ _3365_ _3031_ vssd1 vssd1 vccd1 vccd1 _1827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4302_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _0786_ sky130_fd_sc_hd__inv_2
X_5282_ _0551_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1759_
+ sky130_fd_sc_hd__nand2_1
X_4233_ _0460_ _0455_ vssd1 vssd1 vccd1 vccd1 _0718_ sky130_fd_sc_hd__nand2_1
X_4164_ _3258_ _3251_ vssd1 vssd1 vccd1 vccd1 _0649_ sky130_fd_sc_hd__nand2_1
X_4095_ egd_top.BitStream_buffer.BS_buffer\[3\] vssd1 vssd1 vccd1 vccd1 _0581_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6805_ net159 _0208_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[71\]
+ sky130_fd_sc_hd__dfxtp_1
X_4997_ _0356_ _0362_ _0339_ _0366_ _1475_ vssd1 vssd1 vccd1 vccd1 _1476_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3948_ _3103_ _0395_ vssd1 vssd1 vccd1 vccd1 _0434_ sky130_fd_sc_hd__and2_1
X_3879_ _0364_ vssd1 vssd1 vccd1 vccd1 _0365_ sky130_fd_sc_hd__buf_1
X_5618_ _0441_ _0451_ vssd1 vssd1 vccd1 vccd1 _2092_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5549_ _1776_ _3123_ _2020_ _2021_ _2022_ vssd1 vssd1 vccd1 vccd1 _2023_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4920_ _0494_ _0595_ _0728_ _0598_ vssd1 vssd1 vccd1 vccd1 _1400_ sky130_fd_sc_hd__o22ai_1
X_4851_ _3345_ _3321_ _3335_ _3324_ _1330_ vssd1 vssd1 vccd1 vccd1 _1331_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3802_ _3335_ vssd1 vssd1 vccd1 vccd1 _3336_ sky130_fd_sc_hd__inv_2
X_4782_ _1261_ _1262_ vssd1 vssd1 vccd1 vccd1 _1263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6521_ _2854_ _2855_ vssd1 vssd1 vccd1 vccd1 _2856_ sky130_fd_sc_hd__nand2_1
X_3733_ _3139_ _3228_ vssd1 vssd1 vccd1 vccd1 _3267_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6452_ _2707_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1
+ vccd1 _2793_ sky130_fd_sc_hd__nand2_1
X_3664_ _3197_ vssd1 vssd1 vccd1 vccd1 _3198_ sky130_fd_sc_hd__buf_4
X_5403_ _0551_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1879_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6383_ _2724_ _2725_ vssd1 vssd1 vccd1 vccd1 _2726_ sky130_fd_sc_hd__nand2_1
X_3595_ egd_top.BitStream_buffer.BS_buffer\[68\] vssd1 vssd1 vccd1 vccd1 _3129_ sky130_fd_sc_hd__clkbuf_4
X_5334_ _3271_ _3318_ _3274_ _3322_ vssd1 vssd1 vccd1 vccd1 _1810_ sky130_fd_sc_hd__a22o_1
X_5265_ _0474_ _0689_ vssd1 vssd1 vccd1 vccd1 _1742_ sky130_fd_sc_hd__nand2_1
X_4216_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0701_ sky130_fd_sc_hd__clkbuf_4
X_5196_ _0577_ _3184_ _0573_ _3187_ _1672_ vssd1 vssd1 vccd1 vccd1 _1673_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4147_ _3216_ _3190_ _0631_ vssd1 vssd1 vccd1 vccd1 _0632_ sky130_fd_sc_hd__o21ai_1
X_4078_ _0563_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0564_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2916_ _2916_ vssd1 vssd1 vccd1 vccd1 clknet_0__2916_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3380_ _2932_ vssd1 vssd1 vccd1 vccd1 _2937_ sky130_fd_sc_hd__inv_2
X_5050_ _1465_ _1527_ _1528_ vssd1 vssd1 vccd1 vccd1 _1529_ sky130_fd_sc_hd__nand3_1
X_4001_ _0486_ vssd1 vssd1 vccd1 vccd1 _0487_ sky130_fd_sc_hd__buf_1
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5952_ _2407_ vssd1 vssd1 vccd1 vccd1 _0267_ sky130_fd_sc_hd__clkbuf_1
X_4903_ _0995_ _0518_ vssd1 vssd1 vccd1 vccd1 _1383_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5883_ _0550_ _0493_ vssd1 vssd1 vccd1 vccd1 _2355_ sky130_fd_sc_hd__nand2_1
X_4834_ _3254_ _3272_ vssd1 vssd1 vccd1 vccd1 _1314_ sky130_fd_sc_hd__nand2_1
X_4765_ _3115_ _0450_ _3095_ _0454_ _1245_ vssd1 vssd1 vccd1 vccd1 _1246_ sky130_fd_sc_hd__a221oi_1
X_6504_ _2839_ _2959_ vssd1 vssd1 vccd1 vccd1 _2840_ sky130_fd_sc_hd__nand2_2
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3716_ _3249_ vssd1 vssd1 vccd1 vccd1 _3250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6614__105 clknet_1_0__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__inv_2
X_4696_ _3192_ _3053_ vssd1 vssd1 vccd1 vccd1 _1177_ sky130_fd_sc_hd__nand2_1
X_3647_ _3025_ _3170_ _3028_ _3173_ _3180_ vssd1 vssd1 vccd1 vccd1 _3181_ sky130_fd_sc_hd__a221oi_1
X_6435_ _2653_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1
+ vccd1 vccd1 _2777_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6366_ _2706_ _2708_ vssd1 vssd1 vccd1 vccd1 _2709_ sky130_fd_sc_hd__nand2_2
X_3578_ _3097_ _3087_ vssd1 vssd1 vccd1 vccd1 _3112_ sky130_fd_sc_hd__nor2_2
X_5317_ _3192_ _0552_ vssd1 vssd1 vccd1 vccd1 _1793_ sky130_fd_sc_hd__nand2_1
X_6297_ net8 _3278_ net199 vssd1 vssd1 vccd1 vccd1 _2642_ sky130_fd_sc_hd__mux2_1
X_5248_ _0399_ _0455_ vssd1 vssd1 vccd1 vccd1 _1725_ sky130_fd_sc_hd__nand2_1
X_5179_ _3251_ _3068_ _0646_ _3075_ _1655_ vssd1 vssd1 vccd1 vccd1 _1656_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_66_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4550_ _0900_ _3084_ _1031_ _3092_ vssd1 vssd1 vccd1 vccd1 _1032_ sky130_fd_sc_hd__o22ai_1
X_4481_ _0962_ _0963_ vssd1 vssd1 vccd1 vccd1 _0964_ sky130_fd_sc_hd__nand2_1
X_3501_ egd_top.BitStream_buffer.BS_buffer\[123\] vssd1 vssd1 vccd1 vccd1 _3040_ sky130_fd_sc_hd__clkbuf_4
X_6220_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2592_ sky130_fd_sc_hd__nand2_2
X_3432_ net30 _2953_ net28 _2977_ _2985_ vssd1 vssd1 vccd1 vccd1 _2986_ sky130_fd_sc_hd__a311o_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _2544_ vssd1 vssd1 vccd1 vccd1 _0205_ sky130_fd_sc_hd__clkbuf_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _3344_ _0674_ vssd1 vssd1 vccd1 vccd1 _1580_ sky130_fd_sc_hd__nand2_1
X_6082_ net2 _0703_ _2486_ vssd1 vssd1 vccd1 vccd1 _2497_ sky130_fd_sc_hd__mux2_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _0346_ _0524_ _0353_ _0528_ _1511_ vssd1 vssd1 vccd1 vccd1 _1512_ sky130_fd_sc_hd__a221oi_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5935_ _2932_ vssd1 vssd1 vccd1 vccd1 _2396_ sky130_fd_sc_hd__buf_2
X_5866_ _0473_ _0356_ vssd1 vssd1 vccd1 vccd1 _2338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4817_ _0646_ _3148_ _3265_ _3152_ _1296_ vssd1 vssd1 vccd1 vccd1 _1297_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5797_ _3191_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _2269_
+ sky130_fd_sc_hd__nand2_1
X_4748_ _0388_ _0433_ vssd1 vssd1 vccd1 vccd1 _1229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4679_ _1031_ _3084_ _1159_ _3092_ vssd1 vssd1 vccd1 vccd1 _1160_ sky130_fd_sc_hd__o22ai_1
X_6418_ _2648_ net18 _2649_ _2956_ vssd1 vssd1 vccd1 vccd1 _2760_ sky130_fd_sc_hd__a31o_1
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[6] sky130_fd_sc_hd__buf_12
X_6349_ _2691_ _2669_ vssd1 vssd1 vccd1 vccd1 _2692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3981_ egd_top.BitStream_buffer.BS_buffer\[24\] vssd1 vssd1 vccd1 vccd1 _0467_ sky130_fd_sc_hd__clkbuf_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5720_ _0714_ _0344_ _0853_ _0348_ vssd1 vssd1 vccd1 vccd1 _2193_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _0756_ _0575_ _0596_ _0579_ _2124_ vssd1 vssd1 vccd1 vccd1 _2125_ sky130_fd_sc_hd__o221a_1
X_4602_ _0819_ _3350_ vssd1 vssd1 vccd1 vccd1 _1084_ sky130_fd_sc_hd__or2_1
X_5582_ _3025_ _3302_ _3028_ _3306_ _2055_ vssd1 vssd1 vccd1 vccd1 _2056_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_25_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4533_ _0563_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1016_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4464_ _3357_ _3303_ _0674_ _3307_ _0946_ vssd1 vssd1 vccd1 vccd1 _0947_ sky130_fd_sc_hd__a221oi_1
X_6203_ net11 _3304_ _2557_ vssd1 vssd1 vccd1 vccd1 _2580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4395_ _0866_ _0870_ _0874_ _0878_ vssd1 vssd1 vccd1 vccd1 _0879_ sky130_fd_sc_hd__and4_1
X_3415_ _2949_ vssd1 vssd1 vccd1 vccd1 _2969_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ net2 _3136_ _2521_ vssd1 vssd1 vccd1 vccd1 _2533_ sky130_fd_sc_hd__mux2_1
X_6065_ net200 _3004_ vssd1 vssd1 vccd1 vccd1 _2485_ sky130_fd_sc_hd__or2_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _1484_ _1488_ _1491_ _1494_ vssd1 vssd1 vccd1 vccd1 _1495_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5918_ _2384_ vssd1 vssd1 vccd1 vccd1 _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6898_ net96 _0301_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[124\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5849_ _2311_ _2314_ _2317_ _2320_ vssd1 vssd1 vccd1 vccd1 _2321_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6666__153 clknet_1_1__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__inv_2
XFILLER_0_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4180_ _3330_ _3327_ vssd1 vssd1 vccd1 vccd1 _0665_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6821_ net175 _0224_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[55\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3964_ _0449_ vssd1 vssd1 vccd1 vccd1 _0450_ sky130_fd_sc_hd__clkbuf_4
X_3895_ _3153_ _0324_ vssd1 vssd1 vccd1 vccd1 _0381_ sky130_fd_sc_hd__and2_1
X_5703_ _3325_ _2998_ vssd1 vssd1 vccd1 vccd1 _2176_ sky130_fd_sc_hd__nand2_1
X_5634_ _0511_ _0359_ vssd1 vssd1 vccd1 vccd1 _2108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ _2030_ _2033_ _2036_ _2038_ vssd1 vssd1 vccd1 vccd1 _2039_ sky130_fd_sc_hd__and4_1
X_4516_ _0995_ _0472_ _0996_ _0998_ vssd1 vssd1 vccd1 vccd1 _0999_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5496_ _1034_ _0426_ vssd1 vssd1 vccd1 vccd1 _1971_ sky130_fd_sc_hd__or2_1
X_4447_ _0794_ _3238_ _3287_ _3241_ vssd1 vssd1 vccd1 vccd1 _0930_ sky130_fd_sc_hd__o22ai_1
X_4378_ _0479_ vssd1 vssd1 vccd1 vccd1 _0862_ sky130_fd_sc_hd__inv_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _2520_ vssd1 vssd1 vccd1 vccd1 _2521_ sky130_fd_sc_hd__buf_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ _2473_ vssd1 vssd1 vccd1 vccd1 _0237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2913_ clknet_0__2913_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2913_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3680_ _3213_ vssd1 vssd1 vccd1 vccd1 _3214_ sky130_fd_sc_hd__buf_1
X_5350_ _0634_ _3338_ _1823_ _1824_ _1825_ vssd1 vssd1 vccd1 vccd1 _1826_ sky130_fd_sc_hd__o2111a_1
X_4301_ _3037_ _3184_ _3040_ _3187_ _0784_ vssd1 vssd1 vccd1 vccd1 _0785_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5281_ _0547_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1758_
+ sky130_fd_sc_hd__nand2_1
X_4232_ _0433_ _0432_ _0404_ _0436_ _0716_ vssd1 vssd1 vccd1 vccd1 _0717_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4163_ _3254_ _3247_ vssd1 vssd1 vccd1 vccd1 _0648_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4094_ _0579_ vssd1 vssd1 vccd1 vccd1 _0580_ sky130_fd_sc_hd__clkbuf_4
X_4996_ _1095_ _0369_ _1474_ vssd1 vssd1 vccd1 vccd1 _1475_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6804_ net158 _0207_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[72\]
+ sky130_fd_sc_hd__dfxtp_1
X_3947_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _0433_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3878_ _3112_ _0324_ vssd1 vssd1 vccd1 vccd1 _0364_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6597_ clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2916_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5617_ _3120_ _0413_ _2088_ _2089_ _2090_ vssd1 vssd1 vccd1 vccd1 _2091_ sky130_fd_sc_hd__o2111a_1
X_5548_ _1532_ _3140_ vssd1 vssd1 vccd1 vccd1 _2022_ sky130_fd_sc_hd__or2_1
X_5479_ _0703_ _0328_ _0400_ _0332_ _1953_ vssd1 vssd1 vccd1 vccd1 _1954_ sky130_fd_sc_hd__a221oi_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4850_ _1328_ _1329_ vssd1 vssd1 vccd1 vccd1 _1330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3801_ egd_top.BitStream_buffer.BS_buffer\[103\] vssd1 vssd1 vccd1 vccd1 _3335_ sky130_fd_sc_hd__buf_4
X_6586__79 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__inv_2
X_4781_ _0534_ _0363_ vssd1 vssd1 vccd1 vccd1 _1262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6520_ _2840_ _2847_ _2714_ vssd1 vssd1 vccd1 vccd1 _2855_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3732_ _3265_ vssd1 vssd1 vccd1 vccd1 _3266_ sky130_fd_sc_hd__inv_2
X_6451_ _2730_ _2723_ vssd1 vssd1 vccd1 vccd1 _2792_ sky130_fd_sc_hd__nor2_1
X_3663_ _3196_ vssd1 vssd1 vccd1 vccd1 _3197_ sky130_fd_sc_hd__buf_1
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6382_ _2701_ _2251_ _2668_ vssd1 vssd1 vccd1 vccd1 _2725_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5402_ _0547_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1878_
+ sky130_fd_sc_hd__nand2_1
X_5333_ _0656_ _3264_ _0807_ _3268_ vssd1 vssd1 vccd1 vccd1 _1809_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3594_ _3127_ vssd1 vssd1 vccd1 vccd1 _3128_ sky130_fd_sc_hd__clkbuf_4
X_5264_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _1741_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4215_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0700_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5195_ _0753_ _3190_ _1671_ vssd1 vssd1 vccd1 vccd1 _1672_ sky130_fd_sc_hd__o21ai_1
X_4146_ _3192_ _3040_ vssd1 vssd1 vccd1 vccd1 _0631_ sky130_fd_sc_hd__nand2_1
X_4077_ _0562_ vssd1 vssd1 vccd1 vccd1 _0563_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__2915_ _2915_ vssd1 vssd1 vccd1 vccd1 clknet_0__2915_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4979_ _3344_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _1458_
+ sky130_fd_sc_hd__nand2_1
X_6649_ clknet_1_1__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2920_ sky130_fd_sc_hd__buf_1
XFILLER_0_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4000_ _3109_ _0470_ vssd1 vssd1 vccd1 vccd1 _0486_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5951_ _2406_ _2396_ vssd1 vssd1 vccd1 vccd1 _2407_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _0512_ _0479_ vssd1 vssd1 vccd1 vccd1 _1382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ _0546_ _0513_ vssd1 vssd1 vccd1 vccd1 _2354_ sky130_fd_sc_hd__nand2_1
X_4833_ _3250_ _0804_ vssd1 vssd1 vccd1 vccd1 _1313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4764_ _1034_ _0458_ _1244_ vssd1 vssd1 vccd1 vccd1 _1245_ sky130_fd_sc_hd__o21ai_1
X_6503_ _2833_ _2838_ vssd1 vssd1 vccd1 vccd1 _2839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3715_ _3103_ _3228_ vssd1 vssd1 vccd1 vccd1 _3249_ sky130_fd_sc_hd__and2_1
X_6716__43 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__inv_2
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4695_ _3040_ _3170_ _3044_ _3173_ _1175_ vssd1 vssd1 vccd1 vccd1 _1176_ sky130_fd_sc_hd__a221oi_1
X_6434_ _2773_ _2775_ vssd1 vssd1 vccd1 vccd1 _2776_ sky130_fd_sc_hd__nand2_1
X_3646_ _3174_ _3176_ _3177_ _3179_ vssd1 vssd1 vccd1 vccd1 _3180_ sky130_fd_sc_hd__o22ai_1
X_6731__57 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__inv_2
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6365_ _2707_ _2370_ vssd1 vssd1 vccd1 vccd1 _2708_ sky130_fd_sc_hd__nand2_1
X_3577_ _3110_ vssd1 vssd1 vccd1 vccd1 _3111_ sky130_fd_sc_hd__clkbuf_4
X_6296_ _2641_ vssd1 vssd1 vccd1 vccd1 _0163_ sky130_fd_sc_hd__clkbuf_1
X_5316_ _0607_ _3170_ _0577_ _3173_ _1791_ vssd1 vssd1 vccd1 vccd1 _1792_ sky130_fd_sc_hd__a221oi_1
X_5247_ _1713_ _1717_ _1720_ _1723_ vssd1 vssd1 vccd1 vccd1 _1724_ sky130_fd_sc_hd__and4_1
X_5178_ _1532_ _3084_ _1654_ _3092_ vssd1 vssd1 vccd1 vccd1 _1655_ sky130_fd_sc_hd__o22ai_1
X_4129_ _3115_ vssd1 vssd1 vccd1 vccd1 _0614_ sky130_fd_sc_hd__inv_2
X_6660__148 clknet_1_1__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__inv_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3500_ _3039_ vssd1 vssd1 vccd1 vccd1 _0303_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4480_ _0338_ _0329_ vssd1 vssd1 vccd1 vccd1 _0963_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3431_ egd_top.BitStream_buffer.pc\[6\] _2970_ _2979_ _2984_ vssd1 vssd1 vccd1 vccd1
+ _2985_ sky130_fd_sc_hd__a31o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6150_ _2543_ _2529_ vssd1 vssd1 vccd1 vccd1 _2544_ sky130_fd_sc_hd__and2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _3340_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1579_
+ sky130_fd_sc_hd__nand2_1
X_6081_ _2496_ vssd1 vssd1 vccd1 vccd1 _0227_ sky130_fd_sc_hd__clkbuf_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _1509_ _1510_ vssd1 vssd1 vccd1 vccd1 _1511_ sky130_fd_sc_hd__nand2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5934_ net15 egd_top.BitStream_buffer.BS_buffer\[7\] _2380_ vssd1 vssd1 vccd1 vccd1
+ _2395_ sky130_fd_sc_hd__mux2_1
X_5865_ _2321_ _2336_ vssd1 vssd1 vccd1 vccd1 _2337_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4816_ _1294_ _1295_ vssd1 vssd1 vccd1 vccd1 _1296_ sky130_fd_sc_hd__nand2_1
X_5796_ _0552_ _3169_ _0540_ _3172_ _2267_ vssd1 vssd1 vccd1 vccd1 _2268_ sky130_fd_sc_hd__a221oi_1
X_4747_ _0346_ _0362_ _0353_ _0366_ _1227_ vssd1 vssd1 vccd1 vccd1 _1228_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4678_ _3144_ vssd1 vssd1 vccd1 vccd1 _1159_ sky130_fd_sc_hd__inv_2
X_6417_ _2647_ _2715_ _2718_ _2757_ _2759_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__a32o_2
X_3629_ _3157_ _3162_ vssd1 vssd1 vccd1 vccd1 _3163_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 la_data_out_23_16[7] sky130_fd_sc_hd__buf_12
X_6348_ _2685_ vssd1 vssd1 vccd1 vccd1 _2691_ sky130_fd_sc_hd__inv_4
X_6279_ net14 _0653_ _2613_ vssd1 vssd1 vccd1 vccd1 _2630_ sky130_fd_sc_hd__mux2_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_314 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6710__38 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__inv_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6643__132 clknet_1_1__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__inv_2
X_3980_ _0393_ _0465_ vssd1 vssd1 vccd1 vccd1 _0466_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5650_ _0890_ _0583_ vssd1 vssd1 vccd1 vccd1 _2124_ sky130_fd_sc_hd__or2_1
X_4601_ _3344_ _3297_ vssd1 vssd1 vccd1 vccd1 _1083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5581_ _2053_ _2054_ vssd1 vssd1 vccd1 vccd1 _2055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4532_ _0745_ _0545_ _1012_ _1013_ _1014_ vssd1 vssd1 vccd1 vccd1 _1015_ sky130_fd_sc_hd__o2111a_1
X_4463_ _0944_ _0945_ vssd1 vssd1 vccd1 vccd1 _0946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6202_ _2579_ vssd1 vssd1 vccd1 vccd1 _0189_ sky130_fd_sc_hd__clkbuf_1
X_3414_ egd_top.BitStream_buffer.pc\[6\] _2967_ vssd1 vssd1 vccd1 vccd1 _2968_ sky130_fd_sc_hd__nor2_1
X_4394_ _0359_ _0524_ _0363_ _0528_ _0877_ vssd1 vssd1 vccd1 vccd1 _0878_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ _2532_ vssd1 vssd1 vccd1 vccd1 _0211_ sky130_fd_sc_hd__clkbuf_1
X_6064_ _2484_ vssd1 vssd1 vccd1 vccd1 _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _3102_ _0450_ _3129_ _0454_ _1493_ vssd1 vssd1 vccd1 vccd1 _1494_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5917_ _2383_ _3042_ vssd1 vssd1 vccd1 vccd1 _2384_ sky130_fd_sc_hd__and2_1
X_6897_ net95 _0300_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[125\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5848_ _0421_ _0378_ _0411_ _0382_ _2319_ vssd1 vssd1 vccd1 vccd1 _2320_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5779_ _2251_ _2996_ _2937_ vssd1 vssd1 vccd1 vccd1 _2252_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6820_ net174 _0223_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[56\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _0448_ vssd1 vssd1 vccd1 vccd1 _0449_ sky130_fd_sc_hd__buf_1
X_3894_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _0380_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5702_ _3028_ _3302_ _3031_ _3306_ _2174_ vssd1 vssd1 vccd1 vccd1 _2175_ sky130_fd_sc_hd__a221oi_1
X_5633_ _0507_ _0689_ vssd1 vssd1 vccd1 vccd1 _2107_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5564_ egd_top.BitStream_buffer.BS_buffer\[10\] _3211_ egd_top.BitStream_buffer.BS_buffer\[11\]
+ _3214_ _2037_ vssd1 vssd1 vccd1 vccd1 _2038_ sky130_fd_sc_hd__a221oi_1
X_4515_ _0997_ vssd1 vssd1 vccd1 vccd1 _0998_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5495_ _0420_ _3136_ vssd1 vssd1 vccd1 vccd1 _1970_ sky130_fd_sc_hd__nand2_1
X_4446_ _0918_ _0921_ _0925_ _0928_ vssd1 vssd1 vccd1 vccd1 _0929_ sky130_fd_sc_hd__and4_1
X_4377_ _0843_ _0860_ vssd1 vssd1 vccd1 vccd1 _0861_ sky130_fd_sc_hd__and2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _3002_ _2973_ vssd1 vssd1 vccd1 vccd1 _2520_ sky130_fd_sc_hd__nand2_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _2472_ _2448_ vssd1 vssd1 vccd1 vccd1 _2473_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5280_ _1745_ _1748_ _1752_ _1756_ vssd1 vssd1 vccd1 vccd1 _1757_ sky130_fd_sc_hd__and4_1
X_4300_ _3219_ _3190_ _0783_ vssd1 vssd1 vccd1 vccd1 _0784_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4231_ _0714_ _0440_ _0715_ vssd1 vssd1 vccd1 vccd1 _0716_ sky130_fd_sc_hd__o21ai_1
X_4162_ _3250_ _0646_ vssd1 vssd1 vccd1 vccd1 _0647_ sky130_fd_sc_hd__nand2_1
X_4093_ _3112_ _0543_ vssd1 vssd1 vccd1 vccd1 _0579_ sky130_fd_sc_hd__nand2_1
X_4995_ _0371_ _0323_ vssd1 vssd1 vccd1 vccd1 _1474_ sky130_fd_sc_hd__nand2_1
X_6803_ net157 _0206_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[73\]
+ sky130_fd_sc_hd__dfxtp_1
X_3946_ _0431_ vssd1 vssd1 vccd1 vccd1 _0432_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6600__92 clknet_1_1__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__inv_2
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3877_ egd_top.BitStream_buffer.BS_buffer\[33\] vssd1 vssd1 vccd1 vccd1 _0363_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5616_ _3137_ _0425_ vssd1 vssd1 vccd1 vccd1 _2090_ sky130_fd_sc_hd__or2_1
X_5547_ _3132_ _3259_ vssd1 vssd1 vccd1 vccd1 _2021_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5478_ _1951_ _1952_ vssd1 vssd1 vccd1 vccd1 _1953_ sky130_fd_sc_hd__nand2_1
X_4429_ _3160_ _3149_ vssd1 vssd1 vccd1 vccd1 _0912_ sky130_fd_sc_hd__nand2_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6737__63 clknet_1_0__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__inv_2
XFILLER_0_91_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6752__77 clknet_1_1__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__inv_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4780_ _0530_ _0689_ vssd1 vssd1 vccd1 vccd1 _1261_ sky130_fd_sc_hd__nand2_1
X_3800_ _3318_ _3321_ _3322_ _3324_ _3333_ vssd1 vssd1 vccd1 vccd1 _3334_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3731_ egd_top.BitStream_buffer.BS_buffer\[85\] vssd1 vssd1 vccd1 vccd1 _3265_ sky130_fd_sc_hd__buf_4
XFILLER_0_15_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6450_ _2790_ _2788_ vssd1 vssd1 vccd1 vccd1 _2791_ sky130_fd_sc_hd__nand2_1
X_3662_ _3098_ _3166_ vssd1 vssd1 vccd1 vccd1 _3196_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5401_ _1865_ _1868_ _1872_ _1876_ vssd1 vssd1 vccd1 vccd1 _1877_ sky130_fd_sc_hd__and4_1
X_6381_ _2669_ _2700_ _2013_ vssd1 vssd1 vccd1 vccd1 _2724_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3593_ _3126_ _3065_ vssd1 vssd1 vccd1 vccd1 _3127_ sky130_fd_sc_hd__and2_1
X_5332_ _1804_ _1805_ _1806_ _1807_ vssd1 vssd1 vccd1 vccd1 _1808_ sky130_fd_sc_hd__and4_1
X_5263_ _1724_ _1739_ vssd1 vssd1 vccd1 vccd1 _1740_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4214_ _0684_ _0688_ _0694_ _0698_ vssd1 vssd1 vccd1 vccd1 _0699_ sky130_fd_sc_hd__and4_1
X_5194_ _3192_ _0581_ vssd1 vssd1 vccd1 vccd1 _1671_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4145_ _3028_ _3170_ _3031_ _3173_ _0629_ vssd1 vssd1 vccd1 vccd1 _0630_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4076_ _3061_ _0543_ vssd1 vssd1 vccd1 vccd1 _0562_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_0__2914_ _2914_ vssd1 vssd1 vccd1 vccd1 clknet_0__2914_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4978_ _3340_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _1457_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3929_ _3082_ _0395_ vssd1 vssd1 vccd1 vccd1 _0415_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6579_ _2910_ _2911_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__nand2_1
XFILLER_0_56_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6756__4 clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__inv_2
X_5950_ net10 egd_top.BitStream_buffer.BS_buffer\[12\] _2379_ vssd1 vssd1 vccd1 vccd1
+ _2406_ sky130_fd_sc_hd__mux2_1
X_4901_ _0508_ _0535_ vssd1 vssd1 vccd1 vccd1 _1381_ sky130_fd_sc_hd__nand2_1
X_5881_ _2341_ _2344_ _2348_ _2352_ vssd1 vssd1 vccd1 vccd1 _2353_ sky130_fd_sc_hd__and4_1
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ _3246_ _3275_ vssd1 vssd1 vccd1 vccd1 _1312_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4763_ _0460_ _3102_ vssd1 vssd1 vccd1 vccd1 _1244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4694_ _1047_ _3176_ _1174_ _3179_ vssd1 vssd1 vccd1 vccd1 _1175_ sky130_fd_sc_hd__o22ai_1
X_3714_ _3246_ _3247_ vssd1 vssd1 vccd1 vccd1 _3248_ sky130_fd_sc_hd__nand2_1
X_6502_ _2834_ _2835_ _2689_ _2694_ _2837_ vssd1 vssd1 vccd1 vccd1 _2838_ sky130_fd_sc_hd__o32a_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6433_ _2662_ _2774_ _2688_ vssd1 vssd1 vccd1 vccd1 _2775_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3645_ _3178_ vssd1 vssd1 vccd1 vccd1 _3179_ sky130_fd_sc_hd__clkbuf_4
X_6364_ _2669_ _2700_ vssd1 vssd1 vccd1 vccd1 _2707_ sky130_fd_sc_hd__nor2_4
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3576_ _3109_ _3065_ vssd1 vssd1 vccd1 vccd1 _3110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6295_ _2640_ _2372_ vssd1 vssd1 vccd1 vccd1 _2641_ sky130_fd_sc_hd__and2_1
X_5315_ _0638_ _3176_ _0790_ _3179_ vssd1 vssd1 vccd1 vccd1 _1791_ sky130_fd_sc_hd__o22ai_1
X_5246_ _0703_ _0379_ _0400_ _0383_ _1722_ vssd1 vssd1 vccd1 vccd1 _1723_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5177_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _1654_ sky130_fd_sc_hd__inv_2
X_4128_ _3069_ _3068_ _3161_ _3075_ _0612_ vssd1 vssd1 vccd1 vccd1 _0613_ sky130_fd_sc_hd__a221oi_1
X_4059_ _0544_ vssd1 vssd1 vccd1 vccd1 _0545_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ _2982_ _2983_ _2970_ vssd1 vssd1 vccd1 vccd1 _2984_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6080_ _2495_ _2475_ vssd1 vssd1 vccd1 vccd1 _2496_ sky130_fd_sc_hd__and2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _3314_ _3321_ _3310_ _3324_ _1577_ vssd1 vssd1 vccd1 vccd1 _1578_ sky130_fd_sc_hd__a221oi_1
X_5031_ _0534_ _0372_ vssd1 vssd1 vccd1 vccd1 _1510_ sky130_fd_sc_hd__nand2_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6620__111 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__inv_2
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5933_ _2394_ vssd1 vssd1 vccd1 vccd1 _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5864_ _2325_ _2329_ _2332_ _2335_ vssd1 vssd1 vccd1 vccd1 _2336_ sky130_fd_sc_hd__and4_1
XFILLER_0_75_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4815_ _3160_ _3259_ vssd1 vssd1 vccd1 vccd1 _1295_ sky130_fd_sc_hd__nand2_1
X_5795_ _0574_ _3175_ _0582_ _3178_ vssd1 vssd1 vccd1 vccd1 _2267_ sky130_fd_sc_hd__o22ai_1
X_4746_ _0833_ _0369_ _1226_ vssd1 vssd1 vccd1 vccd1 _1227_ sky130_fd_sc_hd__o21ai_1
X_4677_ _3056_ _1156_ _1158_ vssd1 vssd1 vccd1 vccd1 _0293_ sky130_fd_sc_hd__o21a_1
X_6416_ _2758_ _2713_ vssd1 vssd1 vccd1 vccd1 _2759_ sky130_fd_sc_hd__nand2_1
X_3628_ _3160_ _3161_ vssd1 vssd1 vccd1 vccd1 _3162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 la_data_out_26_24[0] sky130_fd_sc_hd__buf_12
X_6347_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] _2689_ vssd1 vssd1 vccd1
+ vccd1 _2690_ sky130_fd_sc_hd__nor2_1
X_3559_ _3077_ _3084_ _3086_ _3092_ vssd1 vssd1 vccd1 vccd1 _3093_ sky130_fd_sc_hd__o22ai_1
X_6278_ _2629_ vssd1 vssd1 vccd1 vccd1 _0169_ sky130_fd_sc_hd__clkbuf_1
X_5229_ _0916_ _3363_ _1705_ vssd1 vssd1 vccd1 vccd1 _1706_ sky130_fd_sc_hd__o21ai_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4600_ _3340_ _3314_ vssd1 vssd1 vccd1 vccd1 _1082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5580_ _3312_ _3019_ vssd1 vssd1 vccd1 vccd1 _2054_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4531_ _0750_ _0556_ vssd1 vssd1 vccd1 vccd1 _1014_ sky130_fd_sc_hd__or2_1
X_4462_ _3313_ _3304_ vssd1 vssd1 vccd1 vccd1 _0945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6201_ _2578_ _2554_ vssd1 vssd1 vccd1 vccd1 _2579_ sky130_fd_sc_hd__and2_1
X_3413_ _2964_ _2966_ vssd1 vssd1 vccd1 vccd1 _2967_ sky130_fd_sc_hd__and2_1
X_4393_ _0875_ _0876_ vssd1 vssd1 vccd1 vccd1 _0877_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _2531_ _2529_ vssd1 vssd1 vccd1 vccd1 _2532_ sky130_fd_sc_hd__and2_1
X_6063_ _2483_ _2475_ vssd1 vssd1 vccd1 vccd1 _2484_ sky130_fd_sc_hd__and2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _0620_ _0458_ _1492_ vssd1 vssd1 vccd1 vccd1 _1493_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5916_ net6 _0577_ _2380_ vssd1 vssd1 vccd1 vccd1 _2383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6896_ net94 _0299_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[126\]
+ sky130_fd_sc_hd__dfxtp_1
X_5847_ _0848_ _0385_ _2318_ vssd1 vssd1 vccd1 vccd1 _2319_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5778_ egd_top.BitStream_buffer.BitStream_buffer_output\[2\] vssd1 vssd1 vccd1 vccd1
+ _2251_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4729_ _3344_ _3304_ vssd1 vssd1 vccd1 vccd1 _1210_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6627__117 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__inv_2
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5701_ _2172_ _2173_ vssd1 vssd1 vccd1 vccd1 _2174_ sky130_fd_sc_hd__nand2_1
X_3962_ _3158_ _2966_ vssd1 vssd1 vccd1 vccd1 _0448_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3893_ _0378_ vssd1 vssd1 vccd1 vccd1 _0379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5632_ _0535_ _0487_ _0531_ _0491_ _2105_ vssd1 vssd1 vccd1 vccd1 _2106_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5563_ _0745_ _3217_ _0568_ _3220_ vssd1 vssd1 vccd1 vccd1 _2037_ sky130_fd_sc_hd__o22ai_1
X_4514_ _0478_ _0531_ _0481_ _0521_ vssd1 vssd1 vccd1 vccd1 _0997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5494_ _0416_ _3102_ vssd1 vssd1 vccd1 vccd1 _1969_ sky130_fd_sc_hd__nand2_1
X_6686__16 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__inv_2
X_4445_ _0577_ _3212_ _0573_ _3215_ _0927_ vssd1 vssd1 vccd1 vccd1 _0928_ sky130_fd_sc_hd__a221oi_1
X_4376_ _0847_ _0852_ _0856_ _0859_ vssd1 vssd1 vccd1 vccd1 _0860_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6115_ _2519_ vssd1 vssd1 vccd1 vccd1 _0216_ sky130_fd_sc_hd__clkbuf_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ net12 _0323_ _2451_ vssd1 vssd1 vccd1 vccd1 _2472_ sky130_fd_sc_hd__mux2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6879_ net77 _0282_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4230_ _0442_ _0429_ vssd1 vssd1 vccd1 vccd1 _0715_ sky130_fd_sc_hd__nand2_1
X_4161_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _0646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4092_ _0577_ vssd1 vssd1 vccd1 vccd1 _0578_ sky130_fd_sc_hd__inv_2
X_6802_ net156 _0205_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[74\]
+ sky130_fd_sc_hd__dfxtp_1
X_4994_ _1471_ _1472_ vssd1 vssd1 vccd1 vccd1 _1473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3945_ _0430_ vssd1 vssd1 vccd1 vccd1 _0431_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3876_ _0361_ vssd1 vssd1 vccd1 vccd1 _0362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5615_ _0419_ _3134_ vssd1 vssd1 vccd1 vccd1 _2089_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5546_ _3127_ _3255_ vssd1 vssd1 vccd1 vccd1 _2020_ sky130_fd_sc_hd__nand2_1
X_5477_ _0338_ _0433_ vssd1 vssd1 vccd1 vccd1 _1952_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4428_ _3155_ _3255_ vssd1 vssd1 vccd1 vccd1 _0911_ sky130_fd_sc_hd__nand2_1
X_4359_ _0832_ _0836_ _0839_ _0842_ vssd1 vssd1 vccd1 vccd1 _0843_ sky130_fd_sc_hd__and4_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ _2460_ _2448_ vssd1 vssd1 vccd1 vccd1 _2461_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3730_ _3263_ vssd1 vssd1 vccd1 vccd1 _3264_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3661_ _3031_ _3184_ _3034_ _3187_ _3194_ vssd1 vssd1 vccd1 vccd1 _3195_ sky130_fd_sc_hd__a221oi_1
X_5400_ _0339_ _0524_ _0335_ _0528_ _1875_ vssd1 vssd1 vccd1 vccd1 _1876_ sky130_fd_sc_hd__a221oi_1
X_6380_ _2721_ _2722_ vssd1 vssd1 vccd1 vccd1 _2723_ sky130_fd_sc_hd__nand2_1
X_3592_ _3125_ vssd1 vssd1 vccd1 vccd1 _3126_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5331_ _3258_ _3286_ vssd1 vssd1 vccd1 vccd1 _1807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5262_ _1728_ _1732_ _1735_ _1738_ vssd1 vssd1 vccd1 vccd1 _1739_ sky130_fd_sc_hd__and4_1
XFILLER_0_76_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4213_ _0380_ _0379_ _0389_ _0383_ _0697_ vssd1 vssd1 vccd1 vccd1 _0698_ sky130_fd_sc_hd__a221oi_1
X_5193_ _3053_ _3170_ _0607_ _3173_ _1669_ vssd1 vssd1 vccd1 vccd1 _1670_ sky130_fd_sc_hd__a221oi_1
X_4144_ _3177_ _3176_ _0628_ _3179_ vssd1 vssd1 vccd1 vccd1 _0629_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _0560_ vssd1 vssd1 vccd1 vccd1 _0561_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2913_ _2913_ vssd1 vssd1 vccd1 vccd1 clknet_0__2913_ sky130_fd_sc_hd__clkbuf_16
X_4977_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _1456_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3928_ _0413_ vssd1 vssd1 vccd1 vccd1 _0414_ sky130_fd_sc_hd__clkbuf_4
X_3859_ _0344_ vssd1 vssd1 vccd1 vccd1 _0345_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6578_ net18 _2650_ _2956_ _2883_ vssd1 vssd1 vccd1 vccd1 _2911_ sky130_fd_sc_hd__a211o_1
X_5529_ _0734_ _0561_ _2001_ _2002_ _2003_ vssd1 vssd1 vccd1 vccd1 _2004_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6591__84 clknet_1_1__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__inv_2
XFILLER_0_52_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5880_ _0376_ _0523_ _0380_ _0527_ _2351_ vssd1 vssd1 vccd1 vccd1 _2352_ sky130_fd_sc_hd__a221oi_1
X_4900_ _0509_ _0488_ _0503_ _0492_ _1379_ vssd1 vssd1 vccd1 vccd1 _1380_ sky130_fd_sc_hd__a221oi_1
X_4831_ _3318_ _3231_ _3322_ _3235_ _1310_ vssd1 vssd1 vccd1 vccd1 _1311_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4762_ _0701_ _0432_ _0417_ _0436_ _1242_ vssd1 vssd1 vccd1 vccd1 _1243_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4693_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _1174_ sky130_fd_sc_hd__inv_2
X_3713_ egd_top.BitStream_buffer.BS_buffer\[81\] vssd1 vssd1 vccd1 vccd1 _3247_ sky130_fd_sc_hd__clkbuf_4
X_6501_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2836_ vssd1 vssd1
+ vccd1 vccd1 _2837_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6432_ _1652_ _2660_ vssd1 vssd1 vccd1 vccd1 _2774_ sky130_fd_sc_hd__nor2_1
X_3644_ _3139_ _3167_ vssd1 vssd1 vccd1 vccd1 _3178_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6363_ _2669_ _2700_ _2132_ vssd1 vssd1 vccd1 vccd1 _2706_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3575_ _3097_ _3079_ vssd1 vssd1 vccd1 vccd1 _3109_ sky130_fd_sc_hd__nor2_4
X_6294_ net9 _3290_ net199 vssd1 vssd1 vccd1 vccd1 _2640_ sky130_fd_sc_hd__mux2_1
X_5314_ _1778_ _1781_ _1785_ _1789_ vssd1 vssd1 vccd1 vccd1 _1790_ sky130_fd_sc_hd__and4_1
X_5245_ _0705_ _0386_ _1721_ vssd1 vssd1 vccd1 vccd1 _1722_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5176_ _3056_ _1651_ _1653_ vssd1 vssd1 vccd1 vccd1 _0289_ sky130_fd_sc_hd__o21a_1
X_4127_ _3086_ _3084_ _0611_ _3092_ vssd1 vssd1 vccd1 vccd1 _0612_ sky130_fd_sc_hd__o22ai_1
X_4058_ _3139_ _0543_ vssd1 vssd1 vccd1 vccd1 _0544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _0530_ _0691_ vssd1 vssd1 vccd1 vccd1 _1509_ sky130_fd_sc_hd__nand2_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5932_ _2393_ _3042_ vssd1 vssd1 vccd1 vccd1 _2394_ sky130_fd_sc_hd__and2_1
X_5863_ _3057_ _0449_ _3069_ _0453_ _2334_ vssd1 vssd1 vccd1 vccd1 _2335_ sky130_fd_sc_hd__a221oi_1
X_5794_ _2254_ _2257_ _2261_ _2265_ vssd1 vssd1 vccd1 vccd1 _2266_ sky130_fd_sc_hd__and4_1
X_4814_ _3155_ _3251_ vssd1 vssd1 vccd1 vccd1 _1294_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4745_ _0371_ _0339_ vssd1 vssd1 vccd1 vccd1 _1226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4676_ _1157_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1158_ sky130_fd_sc_hd__a21oi_1
X_6415_ _2754_ _2959_ vssd1 vssd1 vccd1 vccd1 _2758_ sky130_fd_sc_hd__nand2_2
X_3627_ egd_top.BitStream_buffer.BS_buffer\[76\] vssd1 vssd1 vccd1 vccd1 _3161_ sky130_fd_sc_hd__clkbuf_4
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 la_data_out_26_24[1] sky130_fd_sc_hd__buf_12
X_6346_ _2688_ vssd1 vssd1 vccd1 vccd1 _2689_ sky130_fd_sc_hd__clkinvlp_2
X_3558_ _3091_ vssd1 vssd1 vccd1 vccd1 _3092_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3489_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _3031_ sky130_fd_sc_hd__clkbuf_4
X_6277_ _2628_ _2372_ vssd1 vssd1 vccd1 vccd1 _2629_ sky130_fd_sc_hd__and2_1
X_5228_ _3365_ _3028_ vssd1 vssd1 vccd1 vccd1 _1705_ sky130_fd_sc_hd__nand2_1
X_5159_ _0551_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1637_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _0551_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _1013_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6650__138 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__inv_2
X_4461_ _3309_ _3353_ vssd1 vssd1 vccd1 vccd1 _0944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6200_ net12 _3297_ _2557_ vssd1 vssd1 vccd1 vccd1 _2578_ sky130_fd_sc_hd__mux2_1
X_3412_ _2965_ egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\] vssd1
+ vssd1 vccd1 vccd1 _2966_ sky130_fd_sc_hd__and3_1
X_4392_ _0534_ _0521_ vssd1 vssd1 vccd1 vccd1 _0876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ net3 _3129_ _2521_ vssd1 vssd1 vccd1 vccd1 _2531_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ net1 _0695_ _2450_ vssd1 vssd1 vccd1 vccd1 _2483_ sky130_fd_sc_hd__mux2_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _0460_ _3136_ vssd1 vssd1 vccd1 vccd1 _1492_ sky130_fd_sc_hd__nand2_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6607__99 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2919_ clknet_0__2919_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2919_
+ sky130_fd_sc_hd__clkbuf_16
X_6895_ net93 _0298_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[127\]
+ sky130_fd_sc_hd__dfxtp_1
X_5915_ _2382_ vssd1 vssd1 vccd1 vccd1 _0279_ sky130_fd_sc_hd__clkbuf_1
X_5846_ _0387_ _0447_ vssd1 vssd1 vccd1 vccd1 _2318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5777_ _2188_ _2248_ _2249_ vssd1 vssd1 vccd1 vccd1 _2250_ sky130_fd_sc_hd__nand3_2
X_4728_ _3340_ _3310_ vssd1 vssd1 vccd1 vccd1 _1209_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4659_ _0551_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _1141_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6329_ _2671_ _2013_ vssd1 vssd1 vccd1 vccd1 _2672_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3961_ egd_top.BitStream_buffer.BS_buffer\[60\] vssd1 vssd1 vccd1 vccd1 _0447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5700_ _3312_ _3022_ vssd1 vssd1 vccd1 vccd1 _2173_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3892_ _0377_ vssd1 vssd1 vccd1 vccd1 _0378_ sky130_fd_sc_hd__buf_1
X_5631_ _1373_ _0495_ _2104_ vssd1 vssd1 vccd1 vccd1 _2105_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5562_ _3050_ _3197_ _3053_ _3200_ _2035_ vssd1 vssd1 vccd1 vccd1 _2036_ sky130_fd_sc_hd__a221oi_1
X_4513_ _0474_ _0535_ vssd1 vssd1 vccd1 vccd1 _0996_ sky130_fd_sc_hd__nand2_1
X_5493_ _3108_ _0397_ _1965_ _1966_ _1967_ vssd1 vssd1 vccd1 vccd1 _1968_ sky130_fd_sc_hd__o2111a_1
X_4444_ _0790_ _3218_ _0926_ _3221_ vssd1 vssd1 vccd1 vccd1 _0927_ sky130_fd_sc_hd__o22ai_1
X_4375_ _0461_ _0450_ _0455_ _0454_ _0858_ vssd1 vssd1 vccd1 vccd1 _0859_ sky130_fd_sc_hd__a221oi_1
X_6114_ _2518_ _2502_ vssd1 vssd1 vccd1 vccd1 _2519_ sky130_fd_sc_hd__and2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _2471_ vssd1 vssd1 vccd1 vccd1 _0238_ sky130_fd_sc_hd__clkbuf_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6878_ net76 _0281_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5829_ _0922_ _3349_ vssd1 vssd1 vccd1 vccd1 _2301_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4160_ _3246_ _3259_ vssd1 vssd1 vccd1 vccd1 _0645_ sky130_fd_sc_hd__nand2_1
X_6691__20 clknet_1_1__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__inv_2
XFILLER_0_4_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ egd_top.BitStream_buffer.BS_buffer\[1\] vssd1 vssd1 vccd1 vccd1 _0577_ sky130_fd_sc_hd__clkbuf_4
X_6801_ net155 _0204_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[75\]
+ sky130_fd_sc_hd__dfxtp_1
X_4993_ _0352_ egd_top.BitStream_buffer.BS_buffer\[45\] _0355_ _0389_ vssd1 vssd1
+ vccd1 vccd1 _1472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3944_ _3098_ _2966_ vssd1 vssd1 vccd1 vccd1 _0430_ sky130_fd_sc_hd__and2_1
X_6656__144 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__inv_2
XFILLER_0_73_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3875_ _0360_ vssd1 vssd1 vccd1 vccd1 _0361_ sky130_fd_sc_hd__buf_1
XFILLER_0_60_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5614_ _0415_ _3129_ vssd1 vssd1 vccd1 vccd1 _2088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5545_ _3144_ _3100_ _3149_ _3105_ _2018_ vssd1 vssd1 vccd1 vccd1 _2019_ sky130_fd_sc_hd__a221oi_1
X_5476_ _0334_ _0404_ vssd1 vssd1 vccd1 vccd1 _1951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4427_ _0611_ _3124_ _0907_ _0908_ _0909_ vssd1 vssd1 vccd1 vccd1 _0910_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_1_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4358_ _0389_ _0379_ _0695_ _0383_ _0841_ vssd1 vssd1 vccd1 vccd1 _0842_ sky130_fd_sc_hd__a221oi_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _3120_ _3141_ vssd1 vssd1 vccd1 vccd1 _0773_ sky130_fd_sc_hd__or2_1
X_6028_ net3 _0691_ _2451_ vssd1 vssd1 vccd1 vccd1 _2460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6728__54 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__inv_2
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3660_ _3188_ _3190_ _3193_ vssd1 vssd1 vccd1 vccd1 _3194_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6743__68 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__inv_2
X_3591_ _3080_ egd_top.BitStream_buffer.pc\[2\] _3096_ vssd1 vssd1 vccd1 vccd1 _3125_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5330_ _3254_ _3225_ vssd1 vssd1 vccd1 vccd1 _1806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5261_ _3136_ _0450_ _3134_ _0454_ _1737_ vssd1 vssd1 vccd1 vccd1 _1738_ sky130_fd_sc_hd__a221oi_1
X_4212_ _0438_ _0386_ _0696_ vssd1 vssd1 vccd1 vccd1 _0697_ sky130_fd_sc_hd__o21ai_1
X_5192_ _3219_ _3176_ _0638_ _3179_ vssd1 vssd1 vccd1 vccd1 _1669_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4143_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _0628_ sky130_fd_sc_hd__inv_2
X_4074_ _3072_ _0543_ vssd1 vssd1 vccd1 vccd1 _0560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4976_ _3335_ _3321_ _3314_ _3324_ _1454_ vssd1 vssd1 vccd1 vccd1 _1455_ sky130_fd_sc_hd__a221oi_1
X_3927_ _3072_ _0395_ vssd1 vssd1 vccd1 vccd1 _0413_ sky130_fd_sc_hd__nand2_1
X_3858_ _3126_ _0325_ vssd1 vssd1 vccd1 vccd1 _0344_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6577_ _2909_ _2756_ vssd1 vssd1 vccd1 vccd1 _2910_ sky130_fd_sc_hd__nand2_1
X_3789_ _3298_ _3244_ vssd1 vssd1 vccd1 vccd1 _3323_ sky130_fd_sc_hd__nor2_1
X_5528_ _0867_ _0570_ vssd1 vssd1 vccd1 vccd1 _2003_ sky130_fd_sc_hd__or2_1
X_5459_ _3309_ _3019_ vssd1 vssd1 vccd1 vccd1 _1934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4830_ _0656_ _3238_ _0807_ _3241_ vssd1 vssd1 vccd1 vccd1 _1310_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4761_ _0394_ _0440_ _1241_ vssd1 vssd1 vccd1 vccd1 _1242_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3712_ _3245_ vssd1 vssd1 vccd1 vccd1 _3246_ sky130_fd_sc_hd__clkbuf_4
X_4692_ _1161_ _1164_ _1168_ _1172_ vssd1 vssd1 vccd1 vccd1 _1173_ sky130_fd_sc_hd__and4_1
X_6500_ _2744_ _2734_ vssd1 vssd1 vccd1 vccd1 _2836_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3643_ _3022_ vssd1 vssd1 vccd1 vccd1 _3177_ sky130_fd_sc_hd__inv_2
X_6431_ _2771_ _2772_ _2733_ vssd1 vssd1 vccd1 vccd1 _2773_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6362_ _2702_ _2704_ vssd1 vssd1 vccd1 vccd1 _2705_ sky130_fd_sc_hd__nor2_1
X_5313_ _0653_ _3148_ _0804_ _3152_ _1788_ vssd1 vssd1 vccd1 vccd1 _1789_ sky130_fd_sc_hd__a221oi_1
X_3574_ _3107_ vssd1 vssd1 vccd1 vccd1 _3108_ sky130_fd_sc_hd__inv_2
X_6293_ _2639_ vssd1 vssd1 vccd1 vccd1 _0164_ sky130_fd_sc_hd__clkbuf_1
X_5244_ _0388_ _0701_ vssd1 vssd1 vccd1 vccd1 _1721_ sky130_fd_sc_hd__nand2_1
X_5175_ _1652_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1653_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4126_ _3057_ vssd1 vssd1 vccd1 vccd1 _0611_ sky130_fd_sc_hd__inv_2
X_4057_ _0542_ vssd1 vssd1 vccd1 vccd1 _0543_ sky130_fd_sc_hd__clkbuf_4
X_4959_ _3254_ _3275_ vssd1 vssd1 vccd1 vccd1 _1438_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6707__35 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__inv_2
XFILLER_0_61_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6722__49 clknet_1_0__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__inv_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5931_ net16 _0548_ _2380_ vssd1 vssd1 vccd1 vccd1 _2393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5862_ _1031_ _0457_ _2333_ vssd1 vssd1 vccd1 vccd1 _2334_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5793_ _3286_ _3147_ _3290_ _3151_ _2264_ vssd1 vssd1 vccd1 vccd1 _2265_ sky130_fd_sc_hd__a221oi_1
X_4813_ _1031_ _3124_ _1290_ _1291_ _1292_ vssd1 vssd1 vccd1 vccd1 _1293_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_90_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4744_ _1223_ _1224_ vssd1 vssd1 vccd1 vccd1 _1225_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] vssd1 vssd1 vccd1 vccd1
+ _1157_ sky130_fd_sc_hd__inv_4
X_6414_ _2714_ _2719_ _2755_ _2756_ vssd1 vssd1 vccd1 vccd1 _2757_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3626_ _3159_ vssd1 vssd1 vccd1 vccd1 _3160_ sky130_fd_sc_hd__clkbuf_4
X_3557_ _3090_ _3065_ vssd1 vssd1 vccd1 vccd1 _3091_ sky130_fd_sc_hd__nand2_1
X_6345_ _2669_ _2687_ vssd1 vssd1 vccd1 vccd1 _2688_ sky130_fd_sc_hd__nor2_2
X_6276_ net15 _3275_ _2613_ vssd1 vssd1 vccd1 vccd1 _2628_ sky130_fd_sc_hd__mux2_1
X_3488_ _3030_ vssd1 vssd1 vccd1 vccd1 _0306_ sky130_fd_sc_hd__clkbuf_1
X_5227_ _3202_ _3338_ _1701_ _1702_ _1703_ vssd1 vssd1 vccd1 vccd1 _1704_ sky130_fd_sc_hd__o2111a_1
X_5158_ _0547_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1636_
+ sky130_fd_sc_hd__nand2_1
X_4109_ _0594_ vssd1 vssd1 vccd1 vccd1 _0595_ sky130_fd_sc_hd__clkbuf_4
X_5089_ _1565_ _1566_ vssd1 vssd1 vccd1 vccd1 _1567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4460_ _0931_ _0936_ _0939_ _0942_ vssd1 vssd1 vccd1 vccd1 _0943_ sky130_fd_sc_hd__and4_1
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4391_ _0530_ _0525_ vssd1 vssd1 vccd1 vccd1 _0875_ sky130_fd_sc_hd__nand2_1
X_3411_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2965_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6130_ _2530_ vssd1 vssd1 vccd1 vccd1 _0212_ sky130_fd_sc_hd__clkbuf_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _2482_ vssd1 vssd1 vccd1 vccd1 _0233_ sky130_fd_sc_hd__clkbuf_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _0423_ _0432_ _0421_ _0436_ _1490_ vssd1 vssd1 vccd1 vccd1 _1491_ sky130_fd_sc_hd__a221oi_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__2918_ clknet_0__2918_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2918_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6894_ net92 _0297_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[15\]
+ sky130_fd_sc_hd__dfxtp_1
X_5914_ _2381_ _3042_ vssd1 vssd1 vccd1 vccd1 _2382_ sky130_fd_sc_hd__and2_1
X_5845_ _0389_ _0361_ _0695_ _0365_ _2316_ vssd1 vssd1 vccd1 vccd1 _2317_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5776_ _0605_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _2249_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4727_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _1208_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4658_ _0547_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _1140_
+ sky130_fd_sc_hd__nand2_1
X_3609_ _3120_ _3124_ _3130_ _3135_ _3142_ vssd1 vssd1 vccd1 vccd1 _3143_ sky130_fd_sc_hd__o2111a_1
X_4589_ _3331_ _3281_ _3327_ _3285_ _1070_ vssd1 vssd1 vccd1 vccd1 _1071_ sky130_fd_sc_hd__a221oi_1
X_6328_ _2670_ _2132_ vssd1 vssd1 vccd1 vccd1 _2671_ sky130_fd_sc_hd__nand2_1
X_6259_ _2616_ _2581_ vssd1 vssd1 vccd1 vccd1 _2617_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3960_ _0429_ _0432_ _0433_ _0436_ _0445_ vssd1 vssd1 vccd1 vccd1 _0446_ sky130_fd_sc_hd__a221oi_1
X_3891_ _3158_ _0324_ vssd1 vssd1 vccd1 vccd1 _0377_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5630_ _0497_ _0525_ vssd1 vssd1 vccd1 vccd1 _2104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5561_ _3216_ _3203_ _2034_ vssd1 vssd1 vccd1 vccd1 _2035_ sky130_fd_sc_hd__o21ai_1
X_4512_ _0482_ vssd1 vssd1 vccd1 vccd1 _0995_ sky130_fd_sc_hd__inv_2
X_5492_ _0767_ _0408_ vssd1 vssd1 vccd1 vccd1 _1967_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ _0607_ vssd1 vssd1 vccd1 vccd1 _0926_ sky130_fd_sc_hd__inv_2
X_4374_ _0614_ _0458_ _0857_ vssd1 vssd1 vccd1 vccd1 _0858_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6113_ net1 _0455_ _2485_ vssd1 vssd1 vccd1 vccd1 _2518_ sky130_fd_sc_hd__mux2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _2470_ _2448_ vssd1 vssd1 vccd1 vccd1 _2471_ sky130_fd_sc_hd__and2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6749__74 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__inv_2
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6877_ net75 _0280_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.buffer_index\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5828_ _3343_ _3019_ vssd1 vssd1 vccd1 vccd1 _2300_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5759_ _2230_ _2231_ vssd1 vssd1 vccd1 vccd1 _2232_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6633__123 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__inv_2
XFILLER_0_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4090_ _0575_ vssd1 vssd1 vccd1 vccd1 _0576_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6800_ net154 _0203_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[76\]
+ sky130_fd_sc_hd__dfxtp_1
X_4992_ _1346_ _0345_ _1470_ _0349_ vssd1 vssd1 vccd1 vccd1 _1471_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3943_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _0429_ sky130_fd_sc_hd__clkbuf_4
X_6662_ clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2921_ sky130_fd_sc_hd__buf_1
X_3874_ _3109_ _0324_ vssd1 vssd1 vccd1 vccd1 _0360_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5613_ _0614_ _0396_ _2084_ _2085_ _2086_ vssd1 vssd1 vccd1 vccd1 _2087_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5544_ _0900_ _3110_ _2017_ vssd1 vssd1 vccd1 vccd1 _2018_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5475_ _1909_ _1920_ _1933_ _1949_ vssd1 vssd1 vccd1 vccd1 _1950_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4426_ _3077_ _3141_ vssd1 vssd1 vccd1 vccd1 _0909_ sky130_fd_sc_hd__or2_1
X_4357_ _0714_ _0386_ _0840_ vssd1 vssd1 vccd1 vccd1 _0841_ sky130_fd_sc_hd__o21ai_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _3133_ _3076_ vssd1 vssd1 vccd1 vccd1 _0772_ sky130_fd_sc_hd__nand2_1
X_6027_ _2459_ vssd1 vssd1 vccd1 vccd1 _0244_ sky130_fd_sc_hd__clkbuf_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _3123_ vssd1 vssd1 vccd1 vccd1 _3124_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_526 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5260_ _3077_ _0458_ _1736_ vssd1 vssd1 vccd1 vccd1 _1737_ sky130_fd_sc_hd__o21ai_1
X_4211_ _0388_ _0695_ vssd1 vssd1 vccd1 vccd1 _0696_ sky130_fd_sc_hd__nand2_1
X_5191_ _1656_ _1659_ _1663_ _1667_ vssd1 vssd1 vccd1 vccd1 _1668_ sky130_fd_sc_hd__and4_1
X_4142_ _0613_ _0617_ _0622_ _0626_ vssd1 vssd1 vccd1 vccd1 _0627_ sky130_fd_sc_hd__and4_1
X_4073_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0559_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4975_ _1452_ _1453_ vssd1 vssd1 vccd1 vccd1 _1454_ sky130_fd_sc_hd__nand2_1
X_3926_ _0411_ vssd1 vssd1 vccd1 vccd1 _0412_ sky130_fd_sc_hd__inv_2
X_6714_ clknet_1_0__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2925_ sky130_fd_sc_hd__buf_1
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3857_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _0343_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6576_ _2904_ _2908_ vssd1 vssd1 vccd1 vccd1 _2909_ sky130_fd_sc_hd__nand2_1
X_3788_ egd_top.BitStream_buffer.BS_buffer\[97\] vssd1 vssd1 vccd1 vccd1 _3322_ sky130_fd_sc_hd__buf_4
X_5527_ _0566_ _0499_ vssd1 vssd1 vccd1 vccd1 _2002_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5458_ _1922_ _1927_ _1930_ _1932_ vssd1 vssd1 vccd1 vccd1 _1933_ sky130_fd_sc_hd__and4_1
X_5389_ _0367_ _0472_ _1862_ _1864_ vssd1 vssd1 vccd1 vccd1 _1865_ sky130_fd_sc_hd__o211a_1
X_4409_ _0883_ _0887_ _0889_ _0892_ vssd1 vssd1 vccd1 vccd1 _0893_ sky130_fd_sc_hd__and4_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4760_ _0442_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _1241_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3711_ _3226_ _3244_ vssd1 vssd1 vccd1 vccd1 _3245_ sky130_fd_sc_hd__nor2_1
X_4691_ _3251_ _3148_ _0646_ _3152_ _1171_ vssd1 vssd1 vccd1 vccd1 _1172_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3642_ _3175_ vssd1 vssd1 vccd1 vccd1 _3176_ sky130_fd_sc_hd__clkbuf_4
X_6430_ _1157_ _2734_ vssd1 vssd1 vccd1 vccd1 _2772_ sky130_fd_sc_hd__nor2_1
X_6361_ _2703_ _0897_ _2666_ vssd1 vssd1 vccd1 vccd1 _2704_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3573_ egd_top.BitStream_buffer.BS_buffer\[64\] vssd1 vssd1 vccd1 vccd1 _3107_ sky130_fd_sc_hd__clkbuf_4
X_5312_ _1786_ _1787_ vssd1 vssd1 vccd1 vccd1 _1788_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6292_ _2638_ _2372_ vssd1 vssd1 vccd1 vccd1 _2639_ sky130_fd_sc_hd__and2_1
X_5243_ _0335_ _0362_ _0323_ _0366_ _1719_ vssd1 vssd1 vccd1 vccd1 _1720_ sky130_fd_sc_hd__a221oi_1
X_5174_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] vssd1 vssd1 vccd1 vccd1
+ _1652_ sky130_fd_sc_hd__inv_2
X_4125_ _3056_ _0609_ _0610_ vssd1 vssd1 vccd1 vccd1 _0297_ sky130_fd_sc_hd__o21a_1
X_4056_ _2965_ _3062_ _3063_ vssd1 vssd1 vccd1 vccd1 _0542_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4958_ _3250_ _3225_ vssd1 vssd1 vccd1 vccd1 _1437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3909_ _2966_ vssd1 vssd1 vccd1 vccd1 _0395_ sky130_fd_sc_hd__buf_2
X_4889_ _3137_ _0458_ _1368_ vssd1 vssd1 vccd1 vccd1 _1369_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6559_ _2844_ _2892_ vssd1 vssd1 vccd1 vccd1 _2893_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5930_ _2392_ vssd1 vssd1 vccd1 vccd1 _0274_ sky130_fd_sc_hd__clkbuf_1
X_5861_ _0459_ _3161_ vssd1 vssd1 vccd1 vccd1 _2333_ sky130_fd_sc_hd__nand2_1
X_5792_ _2262_ _2263_ vssd1 vssd1 vccd1 vccd1 _2264_ sky130_fd_sc_hd__nand2_1
X_4812_ _0764_ _3141_ vssd1 vssd1 vccd1 vccd1 _1292_ sky130_fd_sc_hd__or2_1
X_4743_ _0352_ egd_top.BitStream_buffer.BS_buffer\[43\] _0355_ _0376_ vssd1 vssd1
+ vccd1 vccd1 _1224_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6413_ net17 _2955_ vssd1 vssd1 vccd1 vccd1 _2756_ sky130_fd_sc_hd__nor2_2
X_4674_ _1090_ _1154_ _1155_ vssd1 vssd1 vccd1 vccd1 _1156_ sky130_fd_sc_hd__nand3_1
X_3625_ _3158_ _3065_ vssd1 vssd1 vccd1 vccd1 _3159_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6344_ _2681_ _2685_ _2686_ vssd1 vssd1 vccd1 vccd1 _2687_ sky130_fd_sc_hd__nand3_1
X_3556_ _3089_ vssd1 vssd1 vccd1 vccd1 _3090_ sky130_fd_sc_hd__clkbuf_4
X_6275_ _2627_ vssd1 vssd1 vccd1 vccd1 _0170_ sky130_fd_sc_hd__clkbuf_1
X_3487_ _3029_ _2933_ vssd1 vssd1 vccd1 vccd1 _3030_ sky130_fd_sc_hd__and2_1
X_5226_ _1456_ _3350_ vssd1 vssd1 vccd1 vccd1 _1703_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5157_ _1623_ _1626_ _1630_ _1634_ vssd1 vssd1 vccd1 vccd1 _1635_ sky130_fd_sc_hd__and4_1
X_4108_ _3158_ _0543_ vssd1 vssd1 vccd1 vccd1 _0594_ sky130_fd_sc_hd__nand2_1
X_5088_ _3271_ _3278_ _3274_ _3282_ vssd1 vssd1 vccd1 vccd1 _1566_ sky130_fd_sc_hd__a22o_1
X_4039_ egd_top.BitStream_buffer.BS_buffer\[31\] vssd1 vssd1 vccd1 vccd1 _0525_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6698__27 clknet_1_0__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__inv_2
X_4390_ _0723_ _0506_ _0871_ _0872_ _0873_ vssd1 vssd1 vccd1 vccd1 _0874_ sky130_fd_sc_hd__o2111a_1
X_3410_ _2954_ _2963_ vssd1 vssd1 vccd1 vccd1 _2964_ sky130_fd_sc_hd__nor2_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ _2481_ _2475_ vssd1 vssd1 vccd1 vccd1 _2482_ sky130_fd_sc_hd__and2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _0406_ _0440_ _1489_ vssd1 vssd1 vccd1 vccd1 _1490_ sky130_fd_sc_hd__o21ai_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2917_ clknet_0__2917_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2917_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_451 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6893_ net91 _0296_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ sky130_fd_sc_hd__dfxtp_1
X_5913_ net7 _0607_ _2380_ vssd1 vssd1 vccd1 vccd1 _2381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5844_ _0438_ _0368_ _2315_ vssd1 vssd1 vccd1 vccd1 _2316_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5775_ _2218_ _2234_ _2247_ vssd1 vssd1 vccd1 vccd1 _2248_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4726_ _3347_ _3321_ _3345_ _3324_ _1206_ vssd1 vssd1 vccd1 vccd1 _1207_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4657_ _1127_ _1130_ _1134_ _1138_ vssd1 vssd1 vccd1 vccd1 _1139_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3608_ _3137_ _3141_ vssd1 vssd1 vccd1 vccd1 _3142_ sky130_fd_sc_hd__or2_1
X_6327_ _2251_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2670_ sky130_fd_sc_hd__nand2_1
X_4588_ _0940_ _3289_ _1069_ _3293_ vssd1 vssd1 vccd1 vccd1 _1070_ sky130_fd_sc_hd__o22ai_1
X_3539_ _3072_ _3065_ vssd1 vssd1 vccd1 vccd1 _3073_ sky130_fd_sc_hd__and2_1
X_6258_ net6 _3247_ _2613_ vssd1 vssd1 vccd1 vccd1 _2616_ sky130_fd_sc_hd__mux2_1
X_6189_ _2570_ _2554_ vssd1 vssd1 vccd1 vccd1 _2571_ sky130_fd_sc_hd__and2_1
X_5209_ _1682_ _1683_ _1684_ _1685_ vssd1 vssd1 vccd1 vccd1 _1686_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3890_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _0376_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5560_ _3205_ _3047_ vssd1 vssd1 vccd1 vccd1 _2034_ sky130_fd_sc_hd__nand2_1
X_4511_ _0976_ _0993_ vssd1 vssd1 vccd1 vccd1 _0994_ sky130_fd_sc_hd__and2_1
X_5491_ _0403_ _0455_ vssd1 vssd1 vccd1 vccd1 _1966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4442_ _3022_ _3198_ _3025_ _3201_ _0924_ vssd1 vssd1 vccd1 vccd1 _0925_ sky130_fd_sc_hd__a221oi_1
X_4373_ _0460_ _3107_ vssd1 vssd1 vccd1 vccd1 _0857_ sky130_fd_sc_hd__nand2_1
X_6112_ _2517_ vssd1 vssd1 vccd1 vccd1 _0217_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ net13 _0335_ _2451_ vssd1 vssd1 vccd1 vccd1 _2470_ sky130_fd_sc_hd__mux2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6876_ net74 _0279_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5827_ _3339_ _3013_ vssd1 vssd1 vccd1 vccd1 _2299_ sky130_fd_sc_hd__nand2_1
X_5758_ _0533_ _0335_ vssd1 vssd1 vccd1 vccd1 _2231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4709_ _3254_ _3265_ vssd1 vssd1 vccd1 vccd1 _1190_ sky130_fd_sc_hd__nand2_1
X_5689_ _3249_ _3318_ vssd1 vssd1 vccd1 vccd1 _2162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4991_ egd_top.BitStream_buffer.BS_buffer\[44\] vssd1 vssd1 vccd1 vccd1 _1470_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3942_ _0412_ _0414_ _0418_ _0422_ _0427_ vssd1 vssd1 vccd1 vccd1 _0428_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3873_ egd_top.BitStream_buffer.BS_buffer\[32\] vssd1 vssd1 vccd1 vccd1 _0359_ sky130_fd_sc_hd__buf_4
XFILLER_0_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6617__108 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__inv_2
X_5612_ _0903_ _0407_ vssd1 vssd1 vccd1 vccd1 _2086_ sky130_fd_sc_hd__or2_1
X_5543_ _3113_ _3156_ vssd1 vssd1 vccd1 vccd1 _2017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5474_ _1937_ _1941_ _1945_ _1948_ vssd1 vssd1 vccd1 vccd1 _1949_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4425_ _3133_ _3085_ vssd1 vssd1 vccd1 vccd1 _0908_ sky130_fd_sc_hd__nand2_1
X_4356_ _0388_ _0437_ vssd1 vssd1 vccd1 vccd1 _0840_ sky130_fd_sc_hd__nand2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _3128_ _3134_ vssd1 vssd1 vccd1 vccd1 _0771_ sky130_fd_sc_hd__nand2_1
X_6026_ _2458_ _2448_ vssd1 vssd1 vccd1 vccd1 _2459_ sky130_fd_sc_hd__and2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6588__81 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__inv_2
XFILLER_0_9_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6859_ net57 _0262_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[17\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ egd_top.BitStream_buffer.BS_buffer\[47\] vssd1 vssd1 vccd1 vccd1 _0695_ sky130_fd_sc_hd__clkbuf_4
X_5190_ _3275_ _3148_ _0653_ _3152_ _1666_ vssd1 vssd1 vccd1 vccd1 _1667_ sky130_fd_sc_hd__a221oi_2
X_4141_ _3149_ _3148_ _3255_ _3152_ _0625_ vssd1 vssd1 vccd1 vccd1 _0626_ sky130_fd_sc_hd__a221oi_1
X_4072_ _0541_ _0545_ _0549_ _0553_ _0557_ vssd1 vssd1 vccd1 vccd1 _0558_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4974_ _3330_ _3310_ vssd1 vssd1 vccd1 vccd1 _1453_ sky130_fd_sc_hd__nand2_1
X_3925_ egd_top.BitStream_buffer.BS_buffer\[59\] vssd1 vssd1 vccd1 vccd1 _0411_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3856_ _0323_ _0328_ _0329_ _0332_ _0341_ vssd1 vssd1 vccd1 vccd1 _0342_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6575_ _2906_ _2907_ vssd1 vssd1 vccd1 vccd1 _2908_ sky130_fd_sc_hd__nand2_1
X_3787_ _3320_ vssd1 vssd1 vccd1 vccd1 _3321_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5526_ _0563_ _0515_ vssd1 vssd1 vccd1 vccd1 _2001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5457_ _3310_ _3281_ _3297_ _3285_ _1931_ vssd1 vssd1 vccd1 vccd1 _1932_ sky130_fd_sc_hd__a221oi_1
X_4408_ egd_top.BitStream_buffer.BS_buffer\[16\] _0589_ _0489_ _0592_ _0891_ vssd1
+ vssd1 vccd1 vccd1 _0892_ sky130_fd_sc_hd__a221oi_1
X_5388_ _1863_ vssd1 vssd1 vccd1 vccd1 _1864_ sky130_fd_sc_hd__inv_2
X_4339_ _0819_ _3338_ _0820_ _0821_ _0822_ vssd1 vssd1 vccd1 vccd1 _0823_ sky130_fd_sc_hd__o2111a_1
X_6009_ _2446_ vssd1 vssd1 vccd1 vccd1 _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3710_ _3112_ vssd1 vssd1 vccd1 vccd1 _3244_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4690_ _1169_ _1170_ vssd1 vssd1 vccd1 vccd1 _1171_ sky130_fd_sc_hd__nand2_1
X_3641_ _3126_ _3167_ vssd1 vssd1 vccd1 vccd1 _3175_ sky130_fd_sc_hd__nand2_1
X_6360_ _2687_ vssd1 vssd1 vccd1 vccd1 _2703_ sky130_fd_sc_hd__inv_2
X_3572_ _3105_ vssd1 vssd1 vccd1 vccd1 _3106_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5311_ _3160_ _3272_ vssd1 vssd1 vccd1 vccd1 _1787_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6291_ net10 _3286_ net199 vssd1 vssd1 vccd1 vccd1 _2638_ sky130_fd_sc_hd__mux2_1
X_5242_ _1346_ _0369_ _1718_ vssd1 vssd1 vccd1 vccd1 _1719_ sky130_fd_sc_hd__o21ai_1
X_5173_ _1587_ _1649_ _1650_ vssd1 vssd1 vccd1 vccd1 _1651_ sky130_fd_sc_hd__nand3_1
X_4124_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] _2997_ _2989_ vssd1
+ vssd1 vccd1 vccd1 _0610_ sky130_fd_sc_hd__o21a_1
Xinput1 la_data_in_58_43[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__clkbuf_8
X_4055_ _0540_ vssd1 vssd1 vccd1 vccd1 _0541_ sky130_fd_sc_hd__inv_2
X_4957_ _3246_ _0653_ vssd1 vssd1 vccd1 vccd1 _1436_ sky130_fd_sc_hd__nand2_1
X_3908_ egd_top.BitStream_buffer.BS_buffer\[53\] vssd1 vssd1 vccd1 vccd1 _0394_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4888_ _0460_ _3129_ vssd1 vssd1 vccd1 vccd1 _1368_ sky130_fd_sc_hd__nand2_1
X_3839_ _0324_ vssd1 vssd1 vccd1 vccd1 _0325_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6558_ _2866_ _2959_ _2884_ vssd1 vssd1 vccd1 vccd1 _2892_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5509_ _0690_ _0472_ _1981_ _1983_ vssd1 vssd1 vccd1 vccd1 _1984_ sky130_fd_sc_hd__o211a_1
X_6489_ _2817_ _2818_ vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__nand2_1
X_6669__156 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__inv_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5860_ _3107_ _0431_ _3115_ _0435_ _2331_ vssd1 vssd1 vccd1 vccd1 _2332_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_48_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _3133_ _3161_ vssd1 vssd1 vccd1 vccd1 _1291_ sky130_fd_sc_hd__nand2_1
X_5791_ _3159_ _3225_ vssd1 vssd1 vccd1 vccd1 _2263_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4742_ _1095_ _0345_ _1222_ _0349_ vssd1 vssd1 vccd1 vccd1 _1223_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4673_ _0606_ _0552_ vssd1 vssd1 vccd1 vccd1 _1155_ sky130_fd_sc_hd__nand2_1
X_6412_ _2754_ _2959_ _2712_ vssd1 vssd1 vccd1 vccd1 _2755_ sky130_fd_sc_hd__nand3_1
X_3624_ _2954_ _3079_ vssd1 vssd1 vccd1 vccd1 _3158_ sky130_fd_sc_hd__nor2_4
XFILLER_0_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6677__7 clknet_1_1__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__inv_2
XFILLER_0_11_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6343_ _2996_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] vssd1 vssd1
+ vccd1 vccd1 _2686_ sky130_fd_sc_hd__nor2_2
X_3555_ _3088_ _3060_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3089_
+ sky130_fd_sc_hd__and3_1
X_6712__40 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__inv_2
X_3486_ net15 _3028_ _3007_ vssd1 vssd1 vccd1 vccd1 _3029_ sky130_fd_sc_hd__mux2_1
X_6274_ _2626_ _2581_ vssd1 vssd1 vccd1 vccd1 _2627_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5225_ _3344_ _0675_ vssd1 vssd1 vccd1 vccd1 _1702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5156_ _0353_ _0524_ _0356_ _0528_ _1633_ vssd1 vssd1 vccd1 vccd1 _1634_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5087_ _3287_ _3264_ _3291_ _3268_ vssd1 vssd1 vccd1 vccd1 _1565_ sky130_fd_sc_hd__o22ai_1
X_4107_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0593_ sky130_fd_sc_hd__inv_2
X_4038_ _0523_ vssd1 vssd1 vccd1 vccd1 _0524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ net14 _0467_ _2415_ vssd1 vssd1 vccd1 vccd1 _2433_ sky130_fd_sc_hd__mux2_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _0442_ _0417_ vssd1 vssd1 vccd1 vccd1 _1489_ sky130_fd_sc_hd__nand2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2916_ clknet_0__2916_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2916_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6892_ net90 _0295_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_5912_ _2379_ vssd1 vssd1 vccd1 vccd1 _2380_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5843_ _0370_ _0443_ vssd1 vssd1 vccd1 vccd1 _2315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5774_ _2238_ _2242_ _2244_ _2246_ vssd1 vssd1 vccd1 vccd1 _2247_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4725_ _1204_ _1205_ vssd1 vssd1 vccd1 vccd1 _1206_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4656_ _0689_ _0524_ _0372_ _0528_ _1137_ vssd1 vssd1 vccd1 vccd1 _1138_ sky130_fd_sc_hd__a221oi_1
X_4587_ _3322_ vssd1 vssd1 vccd1 vccd1 _1069_ sky130_fd_sc_hd__inv_2
X_3607_ _3140_ vssd1 vssd1 vccd1 vccd1 _3141_ sky130_fd_sc_hd__buf_2
XFILLER_0_12_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6326_ _2668_ vssd1 vssd1 vccd1 vccd1 _2669_ sky130_fd_sc_hd__inv_6
X_3538_ _3071_ vssd1 vssd1 vccd1 vccd1 _3072_ sky130_fd_sc_hd__buf_2
X_3469_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _3016_ sky130_fd_sc_hd__clkbuf_4
X_6257_ _2615_ vssd1 vssd1 vccd1 vccd1 _0176_ sky130_fd_sc_hd__clkbuf_1
X_6188_ net16 _3345_ _2557_ vssd1 vssd1 vccd1 vccd1 _2570_ sky130_fd_sc_hd__mux2_1
X_5208_ _3258_ _3232_ vssd1 vssd1 vccd1 vccd1 _1685_ sky130_fd_sc_hd__nand2_1
X_5139_ _1606_ _1610_ _1613_ _1616_ vssd1 vssd1 vccd1 vccd1 _1617_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4510_ _0980_ _0985_ _0989_ _0992_ vssd1 vssd1 vccd1 vccd1 _0993_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5490_ _0399_ _3115_ vssd1 vssd1 vccd1 vccd1 _1965_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4441_ _0922_ _3204_ _0923_ vssd1 vssd1 vccd1 vccd1 _0924_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4372_ _0404_ _0432_ _0703_ _0436_ _0855_ vssd1 vssd1 vccd1 vccd1 _0856_ sky130_fd_sc_hd__a221oi_1
X_6111_ _2516_ _2502_ vssd1 vssd1 vccd1 vccd1 _2517_ sky130_fd_sc_hd__and2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _2469_ vssd1 vssd1 vccd1 vccd1 _0239_ sky130_fd_sc_hd__clkbuf_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6875_ net73 _0278_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5826_ _0674_ _3320_ _0675_ _3323_ _2297_ vssd1 vssd1 vccd1 vccd1 _2298_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5757_ _0529_ _0323_ vssd1 vssd1 vccd1 vccd1 _2230_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4708_ _3250_ _0653_ vssd1 vssd1 vccd1 vccd1 _1189_ sky130_fd_sc_hd__nand2_1
X_5688_ _3245_ _3278_ vssd1 vssd1 vccd1 vccd1 _2161_ sky130_fd_sc_hd__nand2_1
X_4639_ _1109_ _1113_ _1117_ _1120_ vssd1 vssd1 vccd1 vccd1 _1121_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6309_ _2651_ _2997_ vssd1 vssd1 vccd1 vccd1 _2652_ sky130_fd_sc_hd__nand2_1
X_6640__129 clknet_1_0__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__inv_2
XFILLER_0_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4990_ _0443_ _0328_ _0429_ _0332_ _1468_ vssd1 vssd1 vccd1 vccd1 _1469_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3941_ _0424_ _0426_ vssd1 vssd1 vccd1 vccd1 _0427_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3872_ _0350_ _0357_ vssd1 vssd1 vccd1 vccd1 _0358_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5611_ _0402_ _3107_ vssd1 vssd1 vccd1 vccd1 _2085_ sky130_fd_sc_hd__nand2_1
X_5542_ _3272_ _3067_ _3275_ _3074_ _2015_ vssd1 vssd1 vccd1 vccd1 _2016_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5473_ _3028_ _3356_ _3031_ _3360_ _1947_ vssd1 vssd1 vccd1 vccd1 _1948_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4424_ _3128_ _3119_ vssd1 vssd1 vccd1 vccd1 _0907_ sky130_fd_sc_hd__nand2_1
X_4355_ _0689_ _0362_ _0372_ _0366_ _0838_ vssd1 vssd1 vccd1 vccd1 _0839_ sky130_fd_sc_hd__a221oi_1
X_6682__12 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__inv_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _3129_ _3101_ _3136_ _3106_ _0769_ vssd1 vssd1 vccd1 vccd1 _0770_ sky130_fd_sc_hd__a221oi_1
X_6025_ net4 _0372_ _2451_ vssd1 vssd1 vccd1 vccd1 _2458_ sky130_fd_sc_hd__mux2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6858_ net56 _0261_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[18\]
+ sky130_fd_sc_hd__dfxtp_1
X_5809_ _3249_ _3322_ vssd1 vssd1 vccd1 vccd1 _2281_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6789_ net143 _0192_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[103\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4140_ _0623_ _0624_ vssd1 vssd1 vccd1 vccd1 _0625_ sky130_fd_sc_hd__nand2_1
X_4071_ _0554_ _0556_ vssd1 vssd1 vccd1 vccd1 _0557_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _3326_ _3297_ vssd1 vssd1 vccd1 vccd1 _1452_ sky130_fd_sc_hd__nand2_1
X_3924_ _0394_ _0397_ _0401_ _0405_ _0409_ vssd1 vssd1 vccd1 vccd1 _0410_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_18_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6719__46 clknet_1_0__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__inv_2
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3855_ _0336_ _0340_ vssd1 vssd1 vccd1 vccd1 _0341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6574_ _2717_ _2712_ vssd1 vssd1 vccd1 vccd1 _2907_ sky130_fd_sc_hd__nor2_1
X_3786_ _3319_ vssd1 vssd1 vccd1 vccd1 _3320_ sky130_fd_sc_hd__buf_1
XFILLER_0_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5525_ _1022_ _0545_ _1997_ _1998_ _1999_ vssd1 vssd1 vccd1 vccd1 _2000_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5456_ _3336_ _3289_ _0668_ _3293_ vssd1 vssd1 vccd1 vccd1 _1931_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4407_ _0756_ _0595_ _0890_ _0598_ vssd1 vssd1 vccd1 vccd1 _0891_ sky130_fd_sc_hd__o22ai_1
X_5387_ _0478_ _0691_ _0481_ _0346_ vssd1 vssd1 vccd1 vccd1 _1863_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4338_ _3336_ _3350_ vssd1 vssd1 vccd1 vccd1 _0822_ sky130_fd_sc_hd__or2_1
X_4269_ _0753_ _0584_ vssd1 vssd1 vccd1 vccd1 _0754_ sky130_fd_sc_hd__or2_1
X_6008_ _2445_ _2423_ vssd1 vssd1 vccd1 vccd1 _2446_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6646__135 clknet_1_1__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__inv_2
XFILLER_0_1_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3640_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _3174_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3571_ _3104_ vssd1 vssd1 vccd1 vccd1 _3105_ sky130_fd_sc_hd__buf_1
X_6290_ _2637_ vssd1 vssd1 vccd1 vccd1 _0165_ sky130_fd_sc_hd__clkbuf_1
X_5310_ _3155_ _3275_ vssd1 vssd1 vccd1 vccd1 _1786_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5241_ _0371_ _0376_ vssd1 vssd1 vccd1 vccd1 _1718_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5172_ _0606_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _1650_
+ sky130_fd_sc_hd__nand2_1
X_4123_ _0322_ _0602_ _0608_ vssd1 vssd1 vccd1 vccd1 _0609_ sky130_fd_sc_hd__nand3_1
Xinput2 la_data_in_58_43[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_8
X_4054_ egd_top.BitStream_buffer.BS_buffer\[5\] vssd1 vssd1 vccd1 vccd1 _0540_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _3322_ _3231_ _3331_ _3235_ _1434_ vssd1 vssd1 vccd1 vccd1 _1435_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3907_ _0342_ _0358_ _0375_ _0392_ vssd1 vssd1 vccd1 vccd1 _0393_ sky130_fd_sc_hd__and4_1
X_4887_ _0417_ _0432_ _0423_ _0436_ _1366_ vssd1 vssd1 vccd1 vccd1 _1367_ sky130_fd_sc_hd__a221oi_1
X_3838_ _2965_ _3062_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _0324_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6557_ _2890_ _2884_ vssd1 vssd1 vccd1 vccd1 _2891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5508_ _1982_ vssd1 vssd1 vccd1 vccd1 _1983_ sky130_fd_sc_hd__inv_2
X_3769_ _3302_ vssd1 vssd1 vccd1 vccd1 _3303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6488_ _2825_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ sky130_fd_sc_hd__inv_2
X_5439_ _0581_ _3184_ _0552_ _3187_ _1913_ vssd1 vssd1 vccd1 vccd1 _1914_ sky130_fd_sc_hd__a221oi_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4810_ _3128_ _3057_ vssd1 vssd1 vccd1 vccd1 _1290_ sky130_fd_sc_hd__nand2_1
X_5790_ _3154_ _3232_ vssd1 vssd1 vccd1 vccd1 _2262_ sky130_fd_sc_hd__nand2_1
X_4741_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _1222_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4672_ _1122_ _1139_ _1153_ vssd1 vssd1 vccd1 vccd1 _1154_ sky130_fd_sc_hd__and3_1
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6411_ _2732_ _2753_ vssd1 vssd1 vccd1 vccd1 _2754_ sky130_fd_sc_hd__nand2_1
X_3623_ _3155_ _3156_ vssd1 vssd1 vccd1 vccd1 _3157_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6342_ _2683_ _2658_ _2684_ vssd1 vssd1 vccd1 vccd1 _2685_ sky130_fd_sc_hd__o21bai_4
X_3554_ _3087_ vssd1 vssd1 vccd1 vccd1 _3088_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3485_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _3028_ sky130_fd_sc_hd__clkbuf_4
X_6273_ net16 _3272_ _2613_ vssd1 vssd1 vccd1 vccd1 _2626_ sky130_fd_sc_hd__mux2_1
X_5224_ _3340_ egd_top.BitStream_buffer.BS_buffer\[109\] vssd1 vssd1 vccd1 vccd1 _1701_
+ sky130_fd_sc_hd__nand2_1
X_5155_ _1631_ _1632_ vssd1 vssd1 vccd1 vccd1 _1633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4106_ _0591_ vssd1 vssd1 vccd1 vccd1 _0592_ sky130_fd_sc_hd__clkbuf_4
X_5086_ _1560_ _1561_ _1562_ _1563_ vssd1 vssd1 vccd1 vccd1 _1564_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4037_ _0522_ vssd1 vssd1 vccd1 vccd1 _0523_ sky130_fd_sc_hd__buf_1
XFILLER_0_63_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _2432_ vssd1 vssd1 vccd1 vccd1 _0256_ sky130_fd_sc_hd__clkbuf_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4939_ _3155_ _0646_ vssd1 vssd1 vccd1 vccd1 _1418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2915_ clknet_0__2915_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2915_
+ sky130_fd_sc_hd__clkbuf_16
X_5911_ _3002_ _2979_ vssd1 vssd1 vccd1 vccd1 _2379_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6891_ net89 _0294_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_5842_ _2312_ _2313_ vssd1 vssd1 vccd1 vccd1 _2314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5773_ _0482_ _0588_ _0535_ _0591_ _2245_ vssd1 vssd1 vccd1 vccd1 _2246_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4724_ _3330_ _3335_ vssd1 vssd1 vccd1 vccd1 _1205_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4655_ _1135_ _1136_ vssd1 vssd1 vccd1 vccd1 _1137_ sky130_fd_sc_hd__nand2_1
X_6689__18 clknet_1_1__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__inv_2
X_4586_ _1066_ _1067_ vssd1 vssd1 vccd1 vccd1 _1068_ sky130_fd_sc_hd__nor2_1
X_3606_ _3139_ _3064_ vssd1 vssd1 vccd1 vccd1 _3140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6325_ _2659_ _2667_ vssd1 vssd1 vccd1 vccd1 _2668_ sky130_fd_sc_hd__nor2_2
X_3537_ _3070_ _3060_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3071_
+ sky130_fd_sc_hd__and3_1
X_3468_ _3015_ vssd1 vssd1 vccd1 vccd1 _0311_ sky130_fd_sc_hd__clkbuf_1
X_6256_ _2614_ _2581_ vssd1 vssd1 vccd1 vccd1 _2615_ sky130_fd_sc_hd__and2_1
X_6187_ _2569_ vssd1 vssd1 vccd1 vccd1 _0194_ sky130_fd_sc_hd__clkbuf_1
X_3399_ net29 vssd1 vssd1 vccd1 vccd1 _2953_ sky130_fd_sc_hd__inv_2
X_5207_ _3254_ _0804_ vssd1 vssd1 vccd1 vccd1 _1684_ sky130_fd_sc_hd__nand2_1
X_5138_ _3129_ _0450_ _3136_ _0454_ _1615_ vssd1 vssd1 vccd1 vccd1 _1616_ sky130_fd_sc_hd__a221oi_1
X_5069_ _3216_ _3176_ _3219_ _3179_ vssd1 vssd1 vccd1 vccd1 _1547_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4440_ _3206_ _3019_ vssd1 vssd1 vccd1 vccd1 _0923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4371_ _0853_ _0440_ _0854_ vssd1 vssd1 vccd1 vccd1 _0855_ sky130_fd_sc_hd__o21ai_1
X_6110_ net8 _0461_ _2485_ vssd1 vssd1 vccd1 vccd1 _2516_ sky130_fd_sc_hd__mux2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _2468_ _2448_ vssd1 vssd1 vccd1 vccd1 _2469_ sky130_fd_sc_hd__and2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6874_ net72 _0277_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6603__95 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__inv_2
X_5825_ _2295_ _2296_ vssd1 vssd1 vccd1 vccd1 _2297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ _0343_ _0505_ _2226_ _2227_ _2228_ vssd1 vssd1 vccd1 vccd1 _2229_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5687_ _3335_ _3230_ _3314_ _3234_ _2159_ vssd1 vssd1 vccd1 vccd1 _2160_ sky130_fd_sc_hd__a221oi_1
X_4707_ _3246_ _3272_ vssd1 vssd1 vccd1 vccd1 _1188_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4638_ _3107_ _0450_ _3115_ _0454_ _1119_ vssd1 vssd1 vccd1 vccd1 _1120_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4569_ _0790_ _3190_ _1050_ vssd1 vssd1 vccd1 vccd1 _1051_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6308_ egd_top.BitStream_buffer.BitStream_buffer_output\[15\] egd_top.BitStream_buffer.BitStream_buffer_output\[14\]
+ vssd1 vssd1 vccd1 vccd1 _2651_ sky130_fd_sc_hd__nor2_1
X_6239_ _2605_ vssd1 vssd1 vccd1 vccd1 _0181_ sky130_fd_sc_hd__inv_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _0425_ vssd1 vssd1 vccd1 vccd1 _0426_ sky130_fd_sc_hd__buf_2
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3871_ _0352_ _0353_ _0355_ _0356_ vssd1 vssd1 vccd1 vccd1 _0357_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5610_ _0398_ _3095_ vssd1 vssd1 vccd1 vccd1 _2084_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5541_ _3262_ _3083_ _3266_ _3091_ vssd1 vssd1 vccd1 vccd1 _2015_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5472_ _1174_ _3363_ _1946_ vssd1 vssd1 vccd1 vccd1 _1947_ sky130_fd_sc_hd__o21ai_1
X_4423_ _3136_ _3101_ _3134_ _3106_ _0905_ vssd1 vssd1 vccd1 vccd1 _0906_ sky130_fd_sc_hd__a221oi_1
X_4354_ _0343_ _0369_ _0837_ vssd1 vssd1 vccd1 vccd1 _0838_ sky130_fd_sc_hd__o21ai_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ _2457_ vssd1 vssd1 vccd1 vccd1 _0245_ sky130_fd_sc_hd__clkbuf_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _0767_ _3111_ _0768_ vssd1 vssd1 vccd1 vccd1 _0769_ sky130_fd_sc_hd__o21ai_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6857_ net55 _0260_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[19\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6788_ net142 _0191_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[104\]
+ sky130_fd_sc_hd__dfxtp_1
X_5808_ _3245_ _3282_ vssd1 vssd1 vccd1 vccd1 _2280_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ _0848_ _0439_ _2211_ vssd1 vssd1 vccd1 vccd1 _2212_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4070_ _0555_ vssd1 vssd1 vccd1 vccd1 _0556_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4972_ _3010_ _3303_ _3013_ _3307_ _1450_ vssd1 vssd1 vccd1 vccd1 _1451_ sky130_fd_sc_hd__a221oi_1
X_3923_ _0406_ _0408_ vssd1 vssd1 vccd1 vccd1 _0409_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3854_ _0338_ _0339_ vssd1 vssd1 vccd1 vccd1 _0340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6573_ _2893_ _2905_ vssd1 vssd1 vccd1 vccd1 _2906_ sky130_fd_sc_hd__nand2_1
X_3785_ _3109_ _3300_ vssd1 vssd1 vccd1 vccd1 _3319_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5524_ _0494_ _0556_ vssd1 vssd1 vccd1 vccd1 _1999_ sky130_fd_sc_hd__or2_1
X_5455_ _1928_ _1929_ vssd1 vssd1 vccd1 vccd1 _1930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _0890_ sky130_fd_sc_hd__inv_2
X_5386_ _0474_ _0372_ vssd1 vssd1 vccd1 vccd1 _1862_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _3344_ _3314_ vssd1 vssd1 vccd1 vccd1 _0821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4268_ _0552_ vssd1 vssd1 vccd1 vccd1 _0753_ sky130_fd_sc_hd__inv_2
X_6007_ net8 _0521_ _2414_ vssd1 vssd1 vccd1 vccd1 _2445_ sky130_fd_sc_hd__mux2_1
X_4199_ _0329_ _0328_ _0376_ _0332_ _0683_ vssd1 vssd1 vccd1 vccd1 _0684_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6909_ net107 _0312_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[113\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3570_ _3103_ _3065_ vssd1 vssd1 vccd1 vccd1 _3104_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _1715_ _1716_ vssd1 vssd1 vccd1 vccd1 _1717_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5171_ _1618_ _1635_ _1648_ vssd1 vssd1 vccd1 vccd1 _1649_ sky130_fd_sc_hd__and3_1
X_4122_ _0606_ _0607_ vssd1 vssd1 vccd1 vccd1 _0608_ sky130_fd_sc_hd__nand2_1
X_4053_ _0485_ _0502_ _0520_ _0538_ vssd1 vssd1 vccd1 vccd1 _0539_ sky130_fd_sc_hd__and4_1
Xinput3 la_data_in_58_43[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _0807_ _3238_ _0940_ _3241_ vssd1 vssd1 vccd1 vccd1 _1434_ sky130_fd_sc_hd__o22ai_1
X_3906_ _0376_ _0379_ _0380_ _0383_ _0391_ vssd1 vssd1 vccd1 vccd1 _0392_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_46_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4886_ _0700_ _0440_ _1365_ vssd1 vssd1 vccd1 vccd1 _1366_ sky130_fd_sc_hd__o21ai_1
X_3837_ egd_top.BitStream_buffer.BS_buffer\[42\] vssd1 vssd1 vccd1 vccd1 _0323_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6556_ _2841_ _2840_ _2867_ vssd1 vssd1 vccd1 vccd1 _2890_ sky130_fd_sc_hd__nand3_1
X_3768_ _3301_ vssd1 vssd1 vccd1 vccd1 _3302_ sky130_fd_sc_hd__buf_1
X_5507_ _0478_ _0346_ _0481_ _0353_ vssd1 vssd1 vccd1 vccd1 _1982_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6487_ _2716_ _2650_ _2667_ vssd1 vssd1 vccd1 vccd1 _2825_ sky130_fd_sc_hd__or3_1
X_3699_ _3072_ _3228_ vssd1 vssd1 vccd1 vccd1 _3233_ sky130_fd_sc_hd__and2_1
X_5438_ _0742_ _3190_ _1912_ vssd1 vssd1 vccd1 vccd1 _1913_ sky130_fd_sc_hd__o21ai_1
X_5369_ _1835_ _1838_ _1841_ _1844_ vssd1 vssd1 vccd1 vccd1 _1845_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6652__140 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__inv_2
XFILLER_0_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4740_ _0695_ _0328_ _0437_ _0332_ _1220_ vssd1 vssd1 vccd1 vccd1 _1221_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4671_ _1143_ _1147_ _1149_ _1152_ vssd1 vssd1 vccd1 vccd1 _1153_ sky130_fd_sc_hd__and4_1
X_6410_ _2741_ _2752_ vssd1 vssd1 vccd1 vccd1 _2753_ sky130_fd_sc_hd__nor2_1
X_3622_ egd_top.BitStream_buffer.BS_buffer\[77\] vssd1 vssd1 vccd1 vccd1 _3156_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6341_ _2655_ _2665_ _2652_ vssd1 vssd1 vccd1 vccd1 _2684_ sky130_fd_sc_hd__a21o_1
X_3553_ _2962_ _3078_ vssd1 vssd1 vccd1 vccd1 _3087_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6272_ _2625_ vssd1 vssd1 vccd1 vccd1 _0171_ sky130_fd_sc_hd__clkbuf_1
X_3484_ _3027_ vssd1 vssd1 vccd1 vccd1 _0307_ sky130_fd_sc_hd__clkbuf_1
X_5223_ _3310_ _3321_ _3297_ _3324_ _1699_ vssd1 vssd1 vccd1 vccd1 _1700_ sky130_fd_sc_hd__a221oi_1
X_5154_ _0534_ _0691_ vssd1 vssd1 vccd1 vccd1 _1632_ sky130_fd_sc_hd__nand2_1
X_4105_ _0590_ vssd1 vssd1 vccd1 vccd1 _0591_ sky130_fd_sc_hd__dlymetal6s2s_1
X_5085_ _3258_ _3225_ vssd1 vssd1 vccd1 vccd1 _1563_ sky130_fd_sc_hd__nand2_1
X_4036_ _3145_ _0469_ vssd1 vssd1 vccd1 vccd1 _0522_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5987_ _2431_ _2423_ vssd1 vssd1 vccd1 vccd1 _2432_ sky130_fd_sc_hd__and2_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4938_ _1159_ _3124_ _1414_ _1415_ _1416_ vssd1 vssd1 vccd1 vccd1 _1417_ sky130_fd_sc_hd__o2111a_1
X_4869_ _1347_ _1348_ vssd1 vssd1 vccd1 vccd1 _1349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6539_ _2866_ _2959_ _2839_ vssd1 vssd1 vccd1 vccd1 _2873_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6703__31 clknet_1_1__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__inv_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__2914_ clknet_0__2914_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2914_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5910_ _2378_ vssd1 vssd1 vccd1 vccd1 _0280_ sky130_fd_sc_hd__clkbuf_1
X_6890_ net88 _0293_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ sky130_fd_sc_hd__dfxtp_2
X_5841_ _0351_ egd_top.BitStream_buffer.BS_buffer\[52\] _0354_ egd_top.BitStream_buffer.BS_buffer\[53\]
+ vssd1 vssd1 vccd1 vccd1 _2313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5772_ _0723_ _0594_ _0862_ _0597_ vssd1 vssd1 vccd1 vccd1 _2245_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4723_ _3326_ _3314_ vssd1 vssd1 vccd1 vccd1 _1204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4654_ _0534_ _0359_ vssd1 vssd1 vccd1 vccd1 _1136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4585_ _3271_ _3225_ _3274_ _3232_ vssd1 vssd1 vccd1 vccd1 _1067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3605_ _3138_ vssd1 vssd1 vccd1 vccd1 _3139_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6324_ _2657_ _2663_ _2666_ vssd1 vssd1 vccd1 vccd1 _2667_ sky130_fd_sc_hd__a21o_1
X_3536_ _2963_ vssd1 vssd1 vccd1 vccd1 _3070_ sky130_fd_sc_hd__inv_2
X_6255_ net7 _3255_ _2613_ vssd1 vssd1 vccd1 vccd1 _2614_ sky130_fd_sc_hd__mux2_1
X_3467_ _3014_ _2933_ vssd1 vssd1 vccd1 vccd1 _3015_ sky130_fd_sc_hd__and2_1
X_5206_ _3250_ _3286_ vssd1 vssd1 vccd1 vccd1 _1683_ sky130_fd_sc_hd__nand2_1
X_6186_ _2568_ _2554_ vssd1 vssd1 vccd1 vccd1 _2569_ sky130_fd_sc_hd__and2_1
X_3398_ _2950_ _2951_ vssd1 vssd1 vccd1 vccd1 _2952_ sky130_fd_sc_hd__and2b_1
X_5137_ _3120_ _0458_ _1614_ vssd1 vssd1 vccd1 vccd1 _1615_ sky130_fd_sc_hd__o21ai_1
X_5068_ _1534_ _1537_ _1541_ _1545_ vssd1 vssd1 vccd1 vccd1 _1546_ sky130_fd_sc_hd__and4_1
X_4019_ _3122_ _0470_ vssd1 vssd1 vccd1 vccd1 _0505_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4370_ _0442_ _0433_ vssd1 vssd1 vccd1 vccd1 _0854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ net14 _0339_ _2451_ vssd1 vssd1 vccd1 vccd1 _2468_ sky130_fd_sc_hd__mux2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6873_ net71 _0276_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_5824_ _3329_ _2998_ vssd1 vssd1 vccd1 vccd1 _2296_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5755_ _0367_ _0517_ vssd1 vssd1 vccd1 vccd1 _2228_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5686_ _3348_ _3237_ _0671_ _3240_ vssd1 vssd1 vccd1 vccd1 _2159_ sky130_fd_sc_hd__o22ai_1
X_4706_ _3282_ _3231_ _3318_ _3235_ _1186_ vssd1 vssd1 vccd1 vccd1 _1187_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4637_ _0903_ _0458_ _1118_ vssd1 vssd1 vccd1 vccd1 _1119_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4568_ _3192_ _3050_ vssd1 vssd1 vccd1 vccd1 _1050_ sky130_fd_sc_hd__nand2_1
X_4499_ _0416_ _0411_ vssd1 vssd1 vccd1 vccd1 _0982_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6307_ _2648_ _2649_ vssd1 vssd1 vccd1 vccd1 _2650_ sky130_fd_sc_hd__and2_2
X_3519_ net1 _3053_ _3006_ vssd1 vssd1 vccd1 vccd1 _3054_ sky130_fd_sc_hd__mux2_1
X_6238_ _2989_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _2605_ sky130_fd_sc_hd__nand2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _2556_ vssd1 vssd1 vccd1 vccd1 _2557_ sky130_fd_sc_hd__buf_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3870_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _0356_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5540_ _3056_ _2012_ _2014_ vssd1 vssd1 vccd1 vccd1 _0286_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5471_ _3365_ _3034_ vssd1 vssd1 vccd1 vccd1 _1946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4422_ _0903_ _3111_ _0904_ vssd1 vssd1 vccd1 vccd1 _0905_ sky130_fd_sc_hd__o21ai_1
X_4353_ _0371_ _0346_ vssd1 vssd1 vccd1 vccd1 _0837_ sky130_fd_sc_hd__nand2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _3114_ _3102_ vssd1 vssd1 vccd1 vccd1 _0768_ sky130_fd_sc_hd__nand2_1
X_6023_ _2456_ _2448_ vssd1 vssd1 vccd1 vccd1 _2457_ sky130_fd_sc_hd__and2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6856_ net54 _0259_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[20\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3999_ _0468_ _0472_ _0476_ _0484_ vssd1 vssd1 vccd1 vccd1 _0485_ sky130_fd_sc_hd__o211a_1
X_6787_ net141 _0190_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[105\]
+ sky130_fd_sc_hd__dfxtp_1
X_5807_ _3314_ _3230_ _3310_ _3234_ _2278_ vssd1 vssd1 vccd1 vccd1 _2279_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5738_ _0441_ _0461_ vssd1 vssd1 vccd1 vccd1 _2211_ sky130_fd_sc_hd__nand2_1
X_6745__70 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__inv_2
XFILLER_0_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5669_ _3262_ _3123_ _2139_ _2140_ _2141_ vssd1 vssd1 vccd1 vccd1 _2142_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6594__87 clknet_1_1__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__inv_2
XFILLER_0_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4971_ _1448_ _1449_ vssd1 vssd1 vccd1 vccd1 _1450_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3922_ _0407_ vssd1 vssd1 vccd1 vccd1 _0408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3853_ egd_top.BitStream_buffer.BS_buffer\[40\] vssd1 vssd1 vccd1 vccd1 _0339_ sky130_fd_sc_hd__clkbuf_4
X_6572_ _2902_ vssd1 vssd1 vccd1 vccd1 _2905_ sky130_fd_sc_hd__inv_2
X_3784_ egd_top.BitStream_buffer.BS_buffer\[96\] vssd1 vssd1 vccd1 vccd1 _3318_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5523_ _0551_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1998_
+ sky130_fd_sc_hd__nand2_1
X_5454_ _3271_ _3322_ _3274_ _3331_ vssd1 vssd1 vccd1 vccd1 _1929_ sky130_fd_sc_hd__a22o_1
X_5385_ _1845_ _1860_ vssd1 vssd1 vccd1 vccd1 _1861_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4405_ _0753_ _0576_ _0582_ _0580_ _0888_ vssd1 vssd1 vccd1 vccd1 _0889_ sky130_fd_sc_hd__o221a_1
X_4336_ _3340_ _3345_ vssd1 vssd1 vccd1 vccd1 _0820_ sky130_fd_sc_hd__nand2_1
X_4267_ _0593_ _0561_ _0748_ _0749_ _0751_ vssd1 vssd1 vccd1 vccd1 _0752_ sky130_fd_sc_hd__o2111a_1
X_6006_ _2444_ vssd1 vssd1 vccd1 vccd1 _0250_ sky130_fd_sc_hd__clkbuf_1
X_4198_ _0681_ _0682_ vssd1 vssd1 vccd1 vccd1 _0683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6908_ net106 _0311_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[114\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6839_ net193 _0242_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[37\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6724__51 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__inv_2
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5170_ _1639_ _1643_ _1645_ _1647_ vssd1 vssd1 vccd1 vccd1 _1648_ sky130_fd_sc_hd__and4_1
X_4121_ egd_top.BitStream_buffer.BS_buffer\[0\] vssd1 vssd1 vccd1 vccd1 _0607_ sky130_fd_sc_hd__clkbuf_4
X_4052_ _0521_ _0524_ _0525_ _0528_ _0537_ vssd1 vssd1 vccd1 vccd1 _0538_ sky130_fd_sc_hd__a221oi_1
Xinput4 la_data_in_58_43[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4954_ _1424_ _1427_ _1430_ _1432_ vssd1 vssd1 vccd1 vccd1 _1433_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3905_ _0384_ _0386_ _0390_ vssd1 vssd1 vccd1 vccd1 _0391_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4885_ _0442_ _0701_ vssd1 vssd1 vccd1 vccd1 _1365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3836_ _3165_ _3224_ _3296_ _3369_ vssd1 vssd1 vccd1 vccd1 _0322_ sky130_fd_sc_hd__and4_1
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6555_ _2888_ _2714_ vssd1 vssd1 vccd1 vccd1 _2889_ sky130_fd_sc_hd__nand2_1
X_3767_ _3061_ _3300_ vssd1 vssd1 vccd1 vccd1 _3301_ sky130_fd_sc_hd__and2_1
X_5506_ _0474_ _0691_ vssd1 vssd1 vccd1 vccd1 _1981_ sky130_fd_sc_hd__nand2_1
X_3698_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _3232_ sky130_fd_sc_hd__clkbuf_4
X_6486_ _2824_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[2\]
+ sky130_fd_sc_hd__inv_2
X_5437_ _3192_ _0540_ vssd1 vssd1 vccd1 vccd1 _1912_ sky130_fd_sc_hd__nand2_1
X_5368_ _0400_ _0379_ _0701_ _0383_ _1843_ vssd1 vssd1 vccd1 vccd1 _1844_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4319_ _0651_ _3264_ _0802_ _3268_ vssd1 vssd1 vccd1 vccd1 _0803_ sky130_fd_sc_hd__o22ai_1
X_5299_ _3056_ _1773_ _1775_ vssd1 vssd1 vccd1 vccd1 _0288_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ _0493_ _0589_ _0499_ _0592_ _1151_ vssd1 vssd1 vccd1 vccd1 _1152_ sky130_fd_sc_hd__a221oi_1
X_3621_ _3154_ vssd1 vssd1 vccd1 vccd1 _3155_ sky130_fd_sc_hd__clkbuf_4
X_6340_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] _2682_ _1652_ _1774_
+ vssd1 vssd1 vccd1 vccd1 _2683_ sky130_fd_sc_hd__o211a_1
X_3552_ _3085_ vssd1 vssd1 vccd1 vccd1 _3086_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6271_ _2624_ _2581_ vssd1 vssd1 vccd1 vccd1 _2625_ sky130_fd_sc_hd__and2_1
X_3483_ _3026_ _2933_ vssd1 vssd1 vccd1 vccd1 _3027_ sky130_fd_sc_hd__and2_1
X_5222_ _1697_ _1698_ vssd1 vssd1 vccd1 vccd1 _1699_ sky130_fd_sc_hd__nand2_1
X_5153_ _0530_ _0346_ vssd1 vssd1 vccd1 vccd1 _1631_ sky130_fd_sc_hd__nand2_1
X_4104_ _2964_ _0542_ vssd1 vssd1 vccd1 vccd1 _0590_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5084_ _3254_ _0653_ vssd1 vssd1 vccd1 vccd1 _1562_ sky130_fd_sc_hd__nand2_1
X_4035_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _0521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5986_ net15 _0503_ _2415_ vssd1 vssd1 vccd1 vccd1 _2431_ sky130_fd_sc_hd__mux2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4937_ _0900_ _3141_ vssd1 vssd1 vccd1 vccd1 _1416_ sky130_fd_sc_hd__or2_1
X_4868_ _0352_ egd_top.BitStream_buffer.BS_buffer\[44\] _0355_ _0380_ vssd1 vssd1
+ vccd1 vccd1 _1348_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3819_ egd_top.BitStream_buffer.BS_buffer\[108\] vssd1 vssd1 vccd1 vccd1 _3353_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ _0606_ _0540_ vssd1 vssd1 vccd1 vccd1 _1280_ sky130_fd_sc_hd__nand2_1
X_6538_ _2871_ _2872_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__nand2_1
XFILLER_0_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6469_ _2803_ _2809_ vssd1 vssd1 vccd1 vccd1 _2810_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__2913_ clknet_0__2913_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2913_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5840_ _0853_ _0344_ _0986_ _0348_ vssd1 vssd1 vccd1 vccd1 _2312_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6659__147 clknet_1_1__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__inv_2
XFILLER_0_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5771_ _0890_ _0575_ _0756_ _0579_ _2243_ vssd1 vssd1 vccd1 vccd1 _2244_ sky130_fd_sc_hd__o221a_1
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4722_ _0675_ _3303_ _2998_ _3307_ _1202_ vssd1 vssd1 vccd1 vccd1 _1203_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4653_ _0530_ _0363_ vssd1 vssd1 vccd1 vccd1 _1135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4584_ _3236_ _3264_ _3239_ _3268_ vssd1 vssd1 vccd1 vccd1 _1066_ sky130_fd_sc_hd__o22ai_1
X_3604_ _3088_ egd_top.BitStream_buffer.pc\[2\] _3096_ vssd1 vssd1 vccd1 vccd1 _3138_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6323_ _2664_ _2665_ vssd1 vssd1 vccd1 vccd1 _2666_ sky130_fd_sc_hd__nand2_2
X_3535_ egd_top.BitStream_buffer.BS_buffer\[75\] vssd1 vssd1 vccd1 vccd1 _3069_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6254_ _2612_ vssd1 vssd1 vccd1 vccd1 _2613_ sky130_fd_sc_hd__buf_4
X_3466_ net5 _3013_ _3007_ vssd1 vssd1 vccd1 vccd1 _3014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5205_ _3246_ _3225_ vssd1 vssd1 vccd1 vccd1 _1682_ sky130_fd_sc_hd__nand2_1
X_6185_ net2 _3347_ _2557_ vssd1 vssd1 vccd1 vccd1 _2568_ sky130_fd_sc_hd__mux2_1
X_3397_ net29 net28 net30 vssd1 vssd1 vccd1 vccd1 _2951_ sky130_fd_sc_hd__a21o_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5136_ _0460_ _3134_ vssd1 vssd1 vccd1 vccd1 _1614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5067_ _3272_ _3148_ _3275_ _3152_ _1544_ vssd1 vssd1 vccd1 vccd1 _1545_ sky130_fd_sc_hd__a221oi_1
X_4018_ _0503_ vssd1 vssd1 vccd1 vccd1 _0504_ sky130_fd_sc_hd__inv_2
XFILLER_0_39_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5969_ _2419_ vssd1 vssd1 vccd1 vccd1 _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6694__23 clknet_1_0__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__inv_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6872_ net70 _0275_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5823_ _3325_ _3010_ vssd1 vssd1 vccd1 vccd1 _2295_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5754_ _0511_ _0363_ vssd1 vssd1 vccd1 vccd1 _2227_ sky130_fd_sc_hd__nand2_1
X_4705_ _3291_ _3238_ _0656_ _3241_ vssd1 vssd1 vccd1 vccd1 _1186_ sky130_fd_sc_hd__o22ai_1
X_5685_ _2149_ _2152_ _2155_ _2157_ vssd1 vssd1 vccd1 vccd1 _2158_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4636_ _0460_ _3095_ vssd1 vssd1 vccd1 vccd1 _1118_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6306_ egd_top.exp_golomb_decoding.te_range\[2\] vssd1 vssd1 vccd1 vccd1 _2649_ sky130_fd_sc_hd__inv_2
X_4567_ _3037_ _3170_ _3040_ _3173_ _1048_ vssd1 vssd1 vccd1 vccd1 _1049_ sky130_fd_sc_hd__a221oi_1
X_4498_ _0461_ vssd1 vssd1 vccd1 vccd1 _0981_ sky130_fd_sc_hd__inv_2
X_3518_ egd_top.BitStream_buffer.BS_buffer\[127\] vssd1 vssd1 vccd1 vccd1 _3053_ sky130_fd_sc_hd__clkbuf_4
X_3449_ _2948_ _2953_ vssd1 vssd1 vccd1 vccd1 _2999_ sky130_fd_sc_hd__nand2_1
X_6237_ egd_top.BitStream_buffer.pc_previous\[4\] _2600_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[4\]
+ sky130_fd_sc_hd__xor2_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _2978_ _2971_ net196 _3002_ vssd1 vssd1 vccd1 vccd1 _2556_ sky130_fd_sc_hd__or4b_2
X_5119_ _1222_ _0369_ _1596_ vssd1 vssd1 vccd1 vccd1 _1597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6099_ _2508_ _2502_ vssd1 vssd1 vccd1 vccd1 _2509_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5470_ _0786_ _3338_ _1942_ _1943_ _1944_ vssd1 vssd1 vccd1 vccd1 _1945_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4421_ _3114_ _3129_ vssd1 vssd1 vccd1 vccd1 _0904_ sky130_fd_sc_hd__nand2_1
X_4352_ _0834_ _0835_ vssd1 vssd1 vccd1 vccd1 _0836_ sky130_fd_sc_hd__nor2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4283_ _3095_ vssd1 vssd1 vccd1 vccd1 _0767_ sky130_fd_sc_hd__inv_2
X_6022_ net5 _0689_ _2451_ vssd1 vssd1 vccd1 vccd1 _2456_ sky130_fd_sc_hd__mux2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6855_ net53 _0258_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[21\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3998_ _0483_ vssd1 vssd1 vccd1 vccd1 _0484_ sky130_fd_sc_hd__inv_2
X_6786_ net140 _0189_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[106\]
+ sky130_fd_sc_hd__dfxtp_1
X_5806_ _0671_ _3237_ _3336_ _3240_ vssd1 vssd1 vccd1 vccd1 _2278_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5737_ _3077_ _0413_ _2207_ _2208_ _2209_ vssd1 vssd1 vccd1 vccd1 _2210_ sky130_fd_sc_hd__o2111a_1
X_5668_ _1654_ _3140_ vssd1 vssd1 vccd1 vccd1 _2141_ sky130_fd_sc_hd__or2_1
X_4619_ _0691_ _0362_ _0346_ _0366_ _1100_ vssd1 vssd1 vccd1 vccd1 _1101_ sky130_fd_sc_hd__a221oi_1
X_5599_ _0400_ _0327_ _0701_ _0331_ _2072_ vssd1 vssd1 vccd1 vccd1 _2073_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4970_ _3313_ _0675_ vssd1 vssd1 vccd1 vccd1 _1449_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3921_ _3122_ _0395_ vssd1 vssd1 vccd1 vccd1 _0407_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3852_ _0337_ vssd1 vssd1 vccd1 vccd1 _0338_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6571_ _2903_ _2714_ vssd1 vssd1 vccd1 vccd1 _2904_ sky130_fd_sc_hd__nand2_1
X_3783_ _3297_ _3303_ _3304_ _3307_ _3316_ vssd1 vssd1 vccd1 vccd1 _3317_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5522_ _0547_ _0489_ vssd1 vssd1 vccd1 vccd1 _1997_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5453_ _0807_ _3264_ _0940_ _3268_ vssd1 vssd1 vccd1 vccd1 _1928_ sky130_fd_sc_hd__o22ai_1
X_5384_ _1849_ _1853_ _1856_ _1859_ vssd1 vssd1 vccd1 vccd1 _1860_ sky130_fd_sc_hd__and4_1
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4404_ _0541_ _0584_ vssd1 vssd1 vccd1 vccd1 _0888_ sky130_fd_sc_hd__or2_1
X_4335_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _0819_ sky130_fd_sc_hd__inv_2
X_4266_ _0750_ _0570_ vssd1 vssd1 vccd1 vccd1 _0751_ sky130_fd_sc_hd__or2_1
X_6005_ _2443_ _2423_ vssd1 vssd1 vccd1 vccd1 _2444_ sky130_fd_sc_hd__and2_1
X_4197_ _0338_ _0335_ vssd1 vssd1 vccd1 vccd1 _0682_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6907_ net105 _0310_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[115\]
+ sky130_fd_sc_hd__dfxtp_1
X_6838_ net192 _0241_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[38\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6769_ net123 _0172_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[84\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4120_ _0605_ vssd1 vssd1 vccd1 vccd1 _0606_ sky130_fd_sc_hd__clkbuf_4
X_4051_ _0532_ _0536_ vssd1 vssd1 vccd1 vccd1 _0537_ sky130_fd_sc_hd__nand2_1
Xinput5 la_data_in_58_43[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4953_ _0540_ _3212_ _0548_ _3215_ _1431_ vssd1 vssd1 vccd1 vccd1 _1432_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3904_ _0388_ _0389_ vssd1 vssd1 vccd1 vccd1 _0390_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4884_ _0614_ _0414_ _1361_ _1362_ _1363_ vssd1 vssd1 vccd1 vccd1 _1364_ sky130_fd_sc_hd__o2111a_1
X_6623_ clknet_1_1__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2918_ sky130_fd_sc_hd__buf_1
XFILLER_0_46_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3835_ _3317_ _3334_ _3352_ _3368_ vssd1 vssd1 vccd1 vccd1 _3369_ sky130_fd_sc_hd__and4_1
X_6554_ _2886_ _2887_ vssd1 vssd1 vccd1 vccd1 _2888_ sky130_fd_sc_hd__nand2_1
X_3766_ _3299_ vssd1 vssd1 vccd1 vccd1 _3300_ sky130_fd_sc_hd__buf_2
X_6485_ _2716_ _2650_ _2685_ vssd1 vssd1 vccd1 vccd1 _2824_ sky130_fd_sc_hd__or3_1
X_5505_ _1964_ _1979_ vssd1 vssd1 vccd1 vccd1 _1980_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3697_ _3230_ vssd1 vssd1 vccd1 vccd1 _3231_ sky130_fd_sc_hd__clkbuf_4
X_5436_ _0577_ _3170_ _0573_ _3173_ _1910_ vssd1 vssd1 vccd1 vccd1 _1911_ sky130_fd_sc_hd__a221oi_1
X_5367_ _0424_ _0386_ _1842_ vssd1 vssd1 vccd1 vccd1 _1843_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4318_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _0802_ sky130_fd_sc_hd__inv_2
X_5298_ _1774_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1775_ sky130_fd_sc_hd__a21oi_1
X_4249_ _0509_ vssd1 vssd1 vccd1 vccd1 _0734_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6613__104 clknet_1_0__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__inv_2
XFILLER_0_60_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3620_ _3153_ _3065_ vssd1 vssd1 vccd1 vccd1 _3154_ sky130_fd_sc_hd__and2_1
X_3551_ egd_top.BitStream_buffer.BS_buffer\[73\] vssd1 vssd1 vccd1 vccd1 _3085_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3482_ net16 _3025_ _3007_ vssd1 vssd1 vccd1 vccd1 _3026_ sky130_fd_sc_hd__mux2_1
X_6270_ net2 _3265_ _2613_ vssd1 vssd1 vccd1 vccd1 _2624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5221_ _3330_ _3304_ vssd1 vssd1 vccd1 vccd1 _1698_ sky130_fd_sc_hd__nand2_1
X_5152_ _1497_ _0506_ _1627_ _1628_ _1629_ vssd1 vssd1 vccd1 vccd1 _1630_ sky130_fd_sc_hd__o2111a_1
X_4103_ _0588_ vssd1 vssd1 vccd1 vccd1 _0589_ sky130_fd_sc_hd__clkbuf_4
X_5083_ _3250_ _3232_ vssd1 vssd1 vccd1 vccd1 _1561_ sky130_fd_sc_hd__nand2_1
X_4034_ _0504_ _0506_ _0510_ _0514_ _0519_ vssd1 vssd1 vccd1 vccd1 _0520_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5985_ _2430_ vssd1 vssd1 vccd1 vccd1 _0257_ sky130_fd_sc_hd__clkbuf_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4936_ _3133_ _3156_ vssd1 vssd1 vccd1 vccd1 _1415_ sky130_fd_sc_hd__nand2_1
X_4867_ _1222_ _0345_ _1346_ _0349_ vssd1 vssd1 vccd1 vccd1 _1347_ sky130_fd_sc_hd__o22ai_1
XANTENNA_10 net5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _3336_ _3338_ _3342_ _3346_ _3351_ vssd1 vssd1 vccd1 vccd1 _3352_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4798_ _1248_ _1265_ _1278_ vssd1 vssd1 vccd1 vccd1 _1279_ sky130_fd_sc_hd__and3_1
X_6537_ _2839_ _2852_ vssd1 vssd1 vccd1 vccd1 _2872_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _2964_ _3227_ vssd1 vssd1 vccd1 vccd1 _3283_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6468_ _2688_ _2807_ _2781_ _2808_ vssd1 vssd1 vccd1 vccd1 _2809_ sky130_fd_sc_hd__a22o_1
X_5419_ _1894_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1895_ sky130_fd_sc_hd__a21oi_1
X_6399_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] egd_top.BitStream_buffer.BitStream_buffer_output\[11\]
+ vssd1 vssd1 vccd1 vccd1 _2742_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5770_ _1022_ _0583_ vssd1 vssd1 vccd1 vccd1 _2243_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4721_ _1200_ _1201_ vssd1 vssd1 vccd1 vccd1 _1202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4652_ _0995_ _0506_ _1131_ _1132_ _1133_ vssd1 vssd1 vccd1 vccd1 _1134_ sky130_fd_sc_hd__o2111a_1
X_3603_ _3136_ vssd1 vssd1 vccd1 vccd1 _3137_ sky130_fd_sc_hd__inv_2
X_4583_ _1061_ _1062_ _1063_ _1064_ vssd1 vssd1 vccd1 vccd1 _1065_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3534_ _3067_ vssd1 vssd1 vccd1 vccd1 _3068_ sky130_fd_sc_hd__clkbuf_4
X_6322_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] egd_top.BitStream_buffer.BitStream_buffer_output\[12\]
+ vssd1 vssd1 vccd1 vccd1 _2665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3465_ egd_top.BitStream_buffer.BS_buffer\[114\] vssd1 vssd1 vccd1 vccd1 _3013_ sky130_fd_sc_hd__clkbuf_4
X_6253_ _2978_ net198 _2972_ _3002_ vssd1 vssd1 vccd1 vccd1 _2612_ sky130_fd_sc_hd__or4b_4
X_5204_ _3327_ _3231_ _3341_ _3235_ _1680_ vssd1 vssd1 vccd1 vccd1 _1681_ sky130_fd_sc_hd__a221oi_1
X_6184_ _2567_ vssd1 vssd1 vccd1 vccd1 _0195_ sky130_fd_sc_hd__clkbuf_1
X_3396_ _2948_ _2949_ vssd1 vssd1 vccd1 vccd1 _2950_ sky130_fd_sc_hd__nor2_1
X_5135_ _0421_ _0432_ _0411_ _0436_ _1612_ vssd1 vssd1 vccd1 vccd1 _1613_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5066_ _1542_ _1543_ vssd1 vssd1 vccd1 vccd1 _1544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4017_ egd_top.BitStream_buffer.BS_buffer\[23\] vssd1 vssd1 vccd1 vccd1 _0503_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5968_ _2418_ _2396_ vssd1 vssd1 vccd1 vccd1 _2419_ sky130_fd_sc_hd__and2_1
XFILLER_0_74_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4919_ _0745_ _0576_ _0554_ _0580_ _1398_ vssd1 vssd1 vccd1 vccd1 _1399_ sky130_fd_sc_hd__o221a_1
X_5899_ _2370_ _2996_ _2937_ vssd1 vssd1 vccd1 vccd1 _2371_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6619__110 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__inv_2
XFILLER_0_53_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6665__152 clknet_1_1__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__inv_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6871_ net69 _0274_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5822_ _3031_ _3302_ _3034_ _3306_ _2293_ vssd1 vssd1 vccd1 vccd1 _2294_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5753_ _0507_ _0372_ vssd1 vssd1 vccd1 vccd1 _2226_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4704_ _1176_ _1179_ _1182_ _1184_ vssd1 vssd1 vccd1 vccd1 _1185_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5684_ egd_top.BitStream_buffer.BS_buffer\[11\] _3211_ egd_top.BitStream_buffer.BS_buffer\[12\]
+ _3214_ _2156_ vssd1 vssd1 vccd1 vccd1 _2157_ sky130_fd_sc_hd__a221oi_1
X_4635_ _0400_ _0432_ _0701_ _0436_ _1116_ vssd1 vssd1 vccd1 vccd1 _1117_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4566_ _0916_ _3176_ _1047_ _3179_ vssd1 vssd1 vccd1 vccd1 _1048_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6305_ net21 _2647_ net20 vssd1 vssd1 vccd1 vccd1 _2648_ sky130_fd_sc_hd__and3b_1
X_3517_ _3052_ vssd1 vssd1 vccd1 vccd1 _0299_ sky130_fd_sc_hd__clkbuf_1
X_4497_ _0705_ _0397_ _0977_ _0978_ _0979_ vssd1 vssd1 vccd1 vccd1 _0980_ sky130_fd_sc_hd__o2111a_1
X_3448_ egd_top.BitStream_buffer.BS_buffer\[112\] vssd1 vssd1 vccd1 vccd1 _2998_ sky130_fd_sc_hd__clkbuf_4
X_6236_ _2604_ vssd1 vssd1 vccd1 vccd1 _0182_ sky130_fd_sc_hd__inv_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ net34 net33 vssd1 vssd1 vccd1 vccd1 _2936_ sky130_fd_sc_hd__nand2_1
X_6167_ _2555_ vssd1 vssd1 vccd1 vccd1 _0200_ sky130_fd_sc_hd__clkbuf_1
X_5118_ _0371_ _0329_ vssd1 vssd1 vccd1 vccd1 _1596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ net12 _0421_ _2486_ vssd1 vssd1 vccd1 vccd1 _2508_ sky130_fd_sc_hd__mux2_1
X_5049_ _0606_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _1528_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4420_ _3102_ vssd1 vssd1 vccd1 vccd1 _0903_ sky130_fd_sc_hd__inv_2
X_4351_ _0352_ _0339_ _0355_ _0335_ vssd1 vssd1 vccd1 vccd1 _0835_ sky130_fd_sc_hd__a22o_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4282_ _3161_ _3068_ _3156_ _3075_ _0765_ vssd1 vssd1 vccd1 vccd1 _0766_ sky130_fd_sc_hd__a221oi_1
X_6021_ _2455_ vssd1 vssd1 vccd1 vccd1 _0246_ sky130_fd_sc_hd__clkbuf_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6854_ net52 _0257_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[22\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3997_ _0478_ _0479_ _0481_ _0482_ vssd1 vssd1 vccd1 vccd1 _0483_ sky130_fd_sc_hd__a22o_1
X_6785_ net139 _0188_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_5805_ _2268_ _2271_ _2274_ _2276_ vssd1 vssd1 vccd1 vccd1 _2277_ sky130_fd_sc_hd__and4_1
X_5736_ _0620_ _0425_ vssd1 vssd1 vccd1 vccd1 _2209_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5667_ _3132_ _3251_ vssd1 vssd1 vccd1 vccd1 _2140_ sky130_fd_sc_hd__nand2_1
X_4618_ _0685_ _0369_ _1099_ vssd1 vssd1 vccd1 vccd1 _1100_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5598_ _2070_ _2071_ vssd1 vssd1 vccd1 vccd1 _2072_ sky130_fd_sc_hd__nand2_1
X_4549_ _3156_ vssd1 vssd1 vccd1 vccd1 _1031_ sky130_fd_sc_hd__inv_2
X_6219_ egd_top.BitStream_buffer.pc_previous\[1\] egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ vssd1 vssd1 vccd1 vccd1 _2591_ sky130_fd_sc_hd__or2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3920_ egd_top.BitStream_buffer.BS_buffer\[55\] vssd1 vssd1 vccd1 vccd1 _0406_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3851_ _3082_ _0325_ vssd1 vssd1 vccd1 vccd1 _0337_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3782_ _3311_ _3315_ vssd1 vssd1 vccd1 vccd1 _3316_ sky130_fd_sc_hd__nand2_1
X_6570_ _2898_ _2902_ vssd1 vssd1 vccd1 vccd1 _2903_ sky130_fd_sc_hd__nand2_1
X_6585__78 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__inv_2
X_5521_ _1984_ _1987_ _1991_ _1995_ vssd1 vssd1 vccd1 vccd1 _1996_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5452_ _1923_ _1924_ _1925_ _1926_ vssd1 vssd1 vccd1 vccd1 _1927_ sky130_fd_sc_hd__and4_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4403_ _0596_ _0561_ _0884_ _0885_ _0886_ vssd1 vssd1 vccd1 vccd1 _0887_ sky130_fd_sc_hd__o2111a_1
X_5383_ _3134_ _0450_ _3119_ _0454_ _1858_ vssd1 vssd1 vccd1 vccd1 _1859_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4334_ _3331_ _3321_ _3327_ _3324_ _0817_ vssd1 vssd1 vccd1 vccd1 _0818_ sky130_fd_sc_hd__a221oi_1
X_6004_ net9 _0531_ _2414_ vssd1 vssd1 vccd1 vccd1 _2443_ sky130_fd_sc_hd__mux2_1
X_4265_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0750_ sky130_fd_sc_hd__inv_2
X_4196_ _0334_ _0323_ vssd1 vssd1 vccd1 vccd1 _0681_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6906_ net104 _0309_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[116\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6837_ net191 _0240_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[39\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6768_ net122 _0171_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[85\]
+ sky130_fd_sc_hd__dfxtp_1
X_5719_ _0701_ _0327_ _0417_ _0331_ _2191_ vssd1 vssd1 vccd1 vccd1 _2192_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4050_ _0534_ _0535_ vssd1 vssd1 vccd1 vccd1 _0536_ sky130_fd_sc_hd__nand2_1
Xinput6 la_data_in_58_43[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _0582_ _3218_ _0753_ _3221_ vssd1 vssd1 vccd1 vccd1 _1431_ sky130_fd_sc_hd__o22ai_1
X_3903_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _0389_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4883_ _0456_ _0426_ vssd1 vssd1 vccd1 vccd1 _1363_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3834_ _3353_ _3356_ _3357_ _3360_ _3367_ vssd1 vssd1 vccd1 vccd1 _3368_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6553_ _2874_ _2875_ _2884_ vssd1 vssd1 vccd1 vccd1 _2887_ sky130_fd_sc_hd__nand3_1
X_3765_ _3298_ vssd1 vssd1 vccd1 vccd1 _3299_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6715__42 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__inv_2
X_6484_ _2823_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.exp_golomb_len\[1\]
+ sky130_fd_sc_hd__inv_2
X_3696_ _3229_ vssd1 vssd1 vccd1 vccd1 _3230_ sky130_fd_sc_hd__buf_1
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5504_ _1968_ _1972_ _1975_ _1978_ vssd1 vssd1 vccd1 vccd1 _1979_ sky130_fd_sc_hd__and4_1
X_5435_ _0790_ _3176_ _0926_ _3179_ vssd1 vssd1 vccd1 vccd1 _1910_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6730__56 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__inv_2
X_5366_ _0388_ _0417_ vssd1 vssd1 vccd1 vccd1 _1842_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4317_ _0797_ _0798_ _0799_ _0800_ vssd1 vssd1 vccd1 vccd1 _0801_ sky130_fd_sc_hd__and4_1
X_5297_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] vssd1 vssd1 vccd1 vccd1
+ _1774_ sky130_fd_sc_hd__inv_2
X_4248_ _0512_ _0515_ vssd1 vssd1 vccd1 vccd1 _0733_ sky130_fd_sc_hd__nand2_1
X_4179_ _3326_ _3341_ vssd1 vssd1 vccd1 vccd1 _0664_ sky130_fd_sc_hd__nand2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3550_ _3083_ vssd1 vssd1 vccd1 vccd1 _3084_ sky130_fd_sc_hd__clkbuf_4
X_3481_ egd_top.BitStream_buffer.BS_buffer\[118\] vssd1 vssd1 vccd1 vccd1 _3025_ sky130_fd_sc_hd__clkbuf_4
X_5220_ _3326_ _3353_ vssd1 vssd1 vccd1 vccd1 _1697_ sky130_fd_sc_hd__nand2_1
X_5151_ _1249_ _0518_ vssd1 vssd1 vccd1 vccd1 _1629_ sky130_fd_sc_hd__or2_1
X_4102_ _0587_ vssd1 vssd1 vccd1 vccd1 _0588_ sky130_fd_sc_hd__buf_1
X_5082_ _3246_ _0804_ vssd1 vssd1 vccd1 vccd1 _1560_ sky130_fd_sc_hd__nand2_1
X_4033_ _0516_ _0518_ vssd1 vssd1 vccd1 vccd1 _0519_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5984_ _2429_ _2423_ vssd1 vssd1 vccd1 vccd1 _2430_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4935_ _3128_ _3069_ vssd1 vssd1 vccd1 vccd1 _1414_ sky130_fd_sc_hd__nand2_1
X_4866_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _1346_ sky130_fd_sc_hd__inv_2
XANTENNA_11 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3817_ _3348_ _3350_ vssd1 vssd1 vccd1 vccd1 _3351_ sky130_fd_sc_hd__or2_1
X_4797_ _1269_ _1273_ _1275_ _1277_ vssd1 vssd1 vccd1 vccd1 _1278_ sky130_fd_sc_hd__and4_1
X_6536_ _2868_ _2870_ _2756_ vssd1 vssd1 vccd1 vccd1 _2871_ sky130_fd_sc_hd__nand3_1
X_3748_ egd_top.BitStream_buffer.BS_buffer\[95\] vssd1 vssd1 vccd1 vccd1 _3282_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6467_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] _2737_ _2744_ vssd1
+ vssd1 vccd1 vccd1 _2808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3679_ _2964_ _3166_ vssd1 vssd1 vccd1 vccd1 _3213_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5418_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1 vssd1 vccd1 vccd1
+ _1894_ sky130_fd_sc_hd__inv_2
X_6398_ _2738_ _2740_ vssd1 vssd1 vccd1 vccd1 _2741_ sky130_fd_sc_hd__nand2_1
X_5349_ _3361_ _3350_ vssd1 vssd1 vccd1 vccd1 _1825_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4720_ _3313_ _3357_ vssd1 vssd1 vccd1 vccd1 _1201_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4651_ _0723_ _0518_ vssd1 vssd1 vccd1 vccd1 _1133_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3602_ egd_top.BitStream_buffer.BS_buffer\[69\] vssd1 vssd1 vccd1 vccd1 _3136_ sky130_fd_sc_hd__clkbuf_4
X_4582_ _3258_ _3272_ vssd1 vssd1 vccd1 vccd1 _1064_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3533_ _3066_ vssd1 vssd1 vccd1 vccd1 _3067_ sky130_fd_sc_hd__buf_1
X_6321_ _2652_ vssd1 vssd1 vccd1 vccd1 _2664_ sky130_fd_sc_hd__inv_2
X_3464_ _3012_ vssd1 vssd1 vccd1 vccd1 _0312_ sky130_fd_sc_hd__clkbuf_1
X_6252_ _2611_ vssd1 vssd1 vccd1 vccd1 _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6183_ _2566_ _2554_ vssd1 vssd1 vccd1 vccd1 _2567_ sky130_fd_sc_hd__and2_1
X_5203_ _1069_ _3238_ _1196_ _3241_ vssd1 vssd1 vccd1 vccd1 _1680_ sky130_fd_sc_hd__o22ai_1
X_5134_ _0705_ _0440_ _1611_ vssd1 vssd1 vccd1 vccd1 _1612_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3395_ net29 net28 vssd1 vssd1 vccd1 vccd1 _2949_ sky130_fd_sc_hd__nor2_1
X_5065_ _3160_ _0646_ vssd1 vssd1 vccd1 vccd1 _1543_ sky130_fd_sc_hd__nand2_1
X_4016_ egd_top.BitStream_buffer.BS_buffer\[16\] _0488_ _0489_ _0492_ _0501_ vssd1
+ vssd1 vccd1 vccd1 _0502_ sky130_fd_sc_hd__a221oi_1
X_6642__131 clknet_1_0__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__inv_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5967_ net6 _0489_ _2415_ vssd1 vssd1 vccd1 vccd1 _2418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _0568_ _0584_ vssd1 vssd1 vccd1 vccd1 _1398_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1 vccd1
+ _2370_ sky130_fd_sc_hd__inv_2
XFILLER_0_35_527 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4849_ _3330_ _3314_ vssd1 vssd1 vccd1 vccd1 _1329_ sky130_fd_sc_hd__nand2_1
X_6519_ _2844_ _2713_ vssd1 vssd1 vccd1 vccd1 _2854_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6754__2 clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__inv_2
X_6870_ net68 _0273_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5821_ _2291_ _2292_ vssd1 vssd1 vccd1 vccd1 _2293_ sky130_fd_sc_hd__nand2_1
X_5752_ _0531_ _0487_ _0521_ _0491_ _2224_ vssd1 vssd1 vccd1 vccd1 _2225_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4703_ _0581_ _3212_ _0552_ _3215_ _1183_ vssd1 vssd1 vccd1 vccd1 _1184_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5683_ _0568_ _3217_ _0750_ _3220_ vssd1 vssd1 vccd1 vccd1 _2156_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4634_ _1114_ _0440_ _1115_ vssd1 vssd1 vccd1 vccd1 _1116_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_508 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4565_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _1047_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6304_ _2646_ vssd1 vssd1 vccd1 vccd1 _2647_ sky130_fd_sc_hd__inv_2
X_3516_ _3051_ _3042_ vssd1 vssd1 vccd1 vccd1 _3052_ sky130_fd_sc_hd__and2_1
X_4496_ _0711_ _0408_ vssd1 vssd1 vccd1 vccd1 _0979_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6235_ _2989_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _2604_ sky130_fd_sc_hd__nand2_1
X_3447_ _2997_ _2987_ _2989_ vssd1 vssd1 vccd1 vccd1 _0314_ sky130_fd_sc_hd__o21ai_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _2928_ _2929_ _2931_ vssd1 vssd1 vccd1 vccd1 _2935_ sky130_fd_sc_hd__a21o_1
X_6166_ _2553_ _2554_ vssd1 vssd1 vccd1 vccd1 _2555_ sky130_fd_sc_hd__and2_1
X_5117_ _1593_ _1594_ vssd1 vssd1 vccd1 vccd1 _1595_ sky130_fd_sc_hd__nor2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _2507_ vssd1 vssd1 vccd1 vccd1 _0222_ sky130_fd_sc_hd__clkbuf_1
X_5048_ _1496_ _1513_ _1526_ vssd1 vssd1 vccd1 vccd1 _1527_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4350_ _0685_ _0345_ _0833_ _0349_ vssd1 vssd1 vccd1 vccd1 _0834_ sky130_fd_sc_hd__o22ai_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ _0611_ _3084_ _0764_ _3092_ vssd1 vssd1 vccd1 vccd1 _0765_ sky130_fd_sc_hd__o22ai_1
X_6020_ _2454_ _2448_ vssd1 vssd1 vccd1 vccd1 _2455_ sky130_fd_sc_hd__and2_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6853_ net51 _0256_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[23\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5804_ egd_top.BitStream_buffer.BS_buffer\[12\] _3211_ egd_top.BitStream_buffer.BS_buffer\[13\]
+ _3214_ _2275_ vssd1 vssd1 vccd1 vccd1 _2276_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_91_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3996_ egd_top.BitStream_buffer.BS_buffer\[27\] vssd1 vssd1 vccd1 vccd1 _0482_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6784_ net138 _0187_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[108\]
+ sky130_fd_sc_hd__dfxtp_1
X_5735_ _0419_ _3119_ vssd1 vssd1 vccd1 vccd1 _2208_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5666_ _3127_ _3247_ vssd1 vssd1 vccd1 vccd1 _2139_ sky130_fd_sc_hd__nand2_1
X_4617_ _0371_ _0356_ vssd1 vssd1 vccd1 vccd1 _1099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5597_ _0337_ _0404_ vssd1 vssd1 vccd1 vccd1 _2071_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4548_ _3056_ _1028_ _1030_ vssd1 vssd1 vccd1 vccd1 _0294_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4479_ _0334_ _0376_ vssd1 vssd1 vccd1 vccd1 _0962_ sky130_fd_sc_hd__nand2_1
X_6218_ _2590_ vssd1 vssd1 vccd1 vccd1 _0184_ sky130_fd_sc_hd__clkbuf_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6149_ net12 _3057_ _2521_ vssd1 vssd1 vccd1 vccd1 _2543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6736__62 clknet_1_0__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__inv_2
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6751__76 clknet_1_1__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__inv_2
XFILLER_0_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3850_ _0334_ _0335_ vssd1 vssd1 vccd1 vccd1 _0336_ sky130_fd_sc_hd__nand2_1
X_3781_ _3313_ _3314_ vssd1 vssd1 vccd1 vccd1 _3315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5520_ _0335_ _0524_ _0323_ _0528_ _1994_ vssd1 vssd1 vccd1 vccd1 _1995_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5451_ _3258_ _3290_ vssd1 vssd1 vccd1 vccd1 _1926_ sky130_fd_sc_hd__nand2_1
X_4402_ _0559_ _0570_ vssd1 vssd1 vccd1 vccd1 _0886_ sky130_fd_sc_hd__or2_1
X_5382_ _3086_ _0458_ _1857_ vssd1 vssd1 vccd1 vccd1 _1858_ sky130_fd_sc_hd__o21ai_1
X_4333_ _0815_ _0816_ vssd1 vssd1 vccd1 vccd1 _0817_ sky130_fd_sc_hd__nand2_1
X_4264_ _0566_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0749_
+ sky130_fd_sc_hd__nand2_1
X_6003_ _2442_ vssd1 vssd1 vccd1 vccd1 _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4195_ _0627_ _0641_ _0659_ _0679_ vssd1 vssd1 vccd1 vccd1 _0680_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6905_ net103 _0308_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[117\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6836_ net190 _0239_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[40\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6767_ net121 _0170_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[86\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5718_ _2189_ _2190_ vssd1 vssd1 vccd1 vccd1 _2191_ sky130_fd_sc_hd__nand2_1
X_3979_ _0410_ _0428_ _0446_ _0464_ vssd1 vssd1 vccd1 vccd1 _0465_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5649_ _0504_ _0560_ _2120_ _2121_ _2122_ vssd1 vssd1 vccd1 vccd1 _2123_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput7 la_data_in_58_43[15] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4951_ _3034_ _3198_ _3037_ _3201_ _1429_ vssd1 vssd1 vccd1 vccd1 _1430_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3902_ _0387_ vssd1 vssd1 vccd1 vccd1 _0388_ sky130_fd_sc_hd__clkbuf_4
X_4882_ _0420_ _3107_ vssd1 vssd1 vccd1 vccd1 _1362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3833_ _3361_ _3363_ _3366_ vssd1 vssd1 vccd1 vccd1 _3367_ sky130_fd_sc_hd__o21ai_1
X_6552_ _2876_ _2885_ vssd1 vssd1 vccd1 vccd1 _2886_ sky130_fd_sc_hd__nand2_1
X_3764_ egd_top.BitStream_buffer.pc\[4\] _2965_ _3063_ vssd1 vssd1 vccd1 vccd1 _3298_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6483_ _2716_ _2650_ _2693_ vssd1 vssd1 vccd1 vccd1 _2823_ sky130_fd_sc_hd__or3_1
X_3695_ _3061_ _3228_ vssd1 vssd1 vccd1 vccd1 _3229_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5503_ _3119_ _0450_ _3076_ _0454_ _1977_ vssd1 vssd1 vccd1 vccd1 _1978_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5434_ _1897_ _1900_ _1904_ _1908_ vssd1 vssd1 vccd1 vccd1 _1909_ sky130_fd_sc_hd__and4_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5365_ _0323_ _0362_ _0329_ _0366_ _1840_ vssd1 vssd1 vccd1 vccd1 _1841_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4316_ _3258_ _0646_ vssd1 vssd1 vccd1 vccd1 _0800_ sky130_fd_sc_hd__nand2_1
X_5296_ _1709_ _1771_ _1772_ vssd1 vssd1 vccd1 vccd1 _1773_ sky130_fd_sc_hd__nand3_1
X_4247_ _0508_ _0503_ vssd1 vssd1 vccd1 vccd1 _0732_ sky130_fd_sc_hd__nand2_1
X_4178_ _3304_ _3303_ _3353_ _3307_ _0662_ vssd1 vssd1 vccd1 vccd1 _0663_ sky130_fd_sc_hd__a221oi_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6819_ net173 _0222_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[57\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3480_ _3024_ vssd1 vssd1 vccd1 vccd1 _0308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5150_ _0512_ _0535_ vssd1 vssd1 vccd1 vccd1 _1628_ sky130_fd_sc_hd__nand2_1
X_4101_ _3145_ _0542_ vssd1 vssd1 vccd1 vccd1 _0587_ sky130_fd_sc_hd__and2_1
X_5081_ _3331_ _3231_ _3327_ _3235_ _1558_ vssd1 vssd1 vccd1 vccd1 _1559_ sky130_fd_sc_hd__a221oi_1
X_4032_ _0517_ vssd1 vssd1 vccd1 vccd1 _0518_ sky130_fd_sc_hd__buf_2
X_5983_ net16 _0509_ _2415_ vssd1 vssd1 vccd1 vccd1 _2429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4934_ _3085_ _3101_ _3057_ _3106_ _1412_ vssd1 vssd1 vccd1 vccd1 _1413_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4865_ _0437_ _0328_ _0443_ _0332_ _1344_ vssd1 vssd1 vccd1 vccd1 _1345_ sky130_fd_sc_hd__a221oi_1
XANTENNA_12 net6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4796_ _0499_ _0589_ _0513_ _0592_ _1276_ vssd1 vssd1 vccd1 vccd1 _1277_ sky130_fd_sc_hd__a221oi_1
X_3816_ _3349_ vssd1 vssd1 vccd1 vccd1 _3350_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6535_ _2854_ _2855_ _2869_ vssd1 vssd1 vccd1 vccd1 _2870_ sky130_fd_sc_hd__nand3_1
X_3747_ _3280_ vssd1 vssd1 vccd1 vccd1 _3281_ sky130_fd_sc_hd__clkbuf_4
X_6466_ _2804_ _2806_ vssd1 vssd1 vccd1 vccd1 _2807_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3678_ _3211_ vssd1 vssd1 vccd1 vccd1 _3212_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6397_ _2703_ _2666_ _2739_ vssd1 vssd1 vccd1 vccd1 _2740_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5417_ _1831_ _1891_ _1892_ vssd1 vssd1 vccd1 vccd1 _1893_ sky130_fd_sc_hd__nand3_1
X_5348_ _3344_ _2998_ vssd1 vssd1 vccd1 vccd1 _1824_ sky130_fd_sc_hd__nand2_1
X_5279_ _0356_ _0524_ _0339_ _0528_ _1755_ vssd1 vssd1 vccd1 vccd1 _1756_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _0512_ _0467_ vssd1 vssd1 vccd1 vccd1 _1132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 la_data_in_58_43[3] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3601_ _3133_ _3134_ vssd1 vssd1 vccd1 vccd1 _3135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4581_ _3254_ _0646_ vssd1 vssd1 vccd1 vccd1 _1063_ sky130_fd_sc_hd__nand2_1
X_6320_ _2662_ _2013_ vssd1 vssd1 vccd1 vccd1 _2663_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3532_ _3061_ _3065_ vssd1 vssd1 vccd1 vccd1 _3066_ sky130_fd_sc_hd__and2_1
X_3463_ _3011_ _2933_ vssd1 vssd1 vccd1 vccd1 _3012_ sky130_fd_sc_hd__and2_1
X_6251_ _2962_ _2989_ vssd1 vssd1 vccd1 vccd1 _2611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6182_ net3 _3341_ _2557_ vssd1 vssd1 vccd1 vccd1 _2566_ sky130_fd_sc_hd__mux2_1
X_5202_ _1670_ _1673_ _1676_ _1678_ vssd1 vssd1 vccd1 vccd1 _1679_ sky130_fd_sc_hd__and4_1
X_5133_ _0442_ _0423_ vssd1 vssd1 vccd1 vccd1 _1611_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3394_ net30 vssd1 vssd1 vccd1 vccd1 _2948_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5064_ _3155_ _3265_ vssd1 vssd1 vccd1 vccd1 _1542_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4015_ _0494_ _0496_ _0500_ vssd1 vssd1 vccd1 vccd1 _0501_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5966_ _2417_ vssd1 vssd1 vccd1 vccd1 _0263_ sky130_fd_sc_hd__clkbuf_1
X_5897_ _2307_ _2367_ _2368_ vssd1 vssd1 vccd1 vccd1 _2369_ sky130_fd_sc_hd__nand3_2
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4917_ _1150_ _0561_ _1394_ _1395_ _1396_ vssd1 vssd1 vccd1 vccd1 _1397_ sky130_fd_sc_hd__o2111a_1
X_4848_ _3326_ _3310_ vssd1 vssd1 vccd1 vccd1 _1328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _1123_ _0506_ _1257_ _1258_ _1259_ vssd1 vssd1 vccd1 vccd1 _1260_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_62_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6518_ _2845_ _2851_ _2853_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__o21ai_2
X_6449_ _2758_ _2786_ _2714_ vssd1 vssd1 vccd1 vccd1 _2790_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6626__116 clknet_1_0__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__inv_2
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5820_ _3312_ _3025_ vssd1 vssd1 vccd1 vccd1 _2292_ sky130_fd_sc_hd__nand2_1
X_5751_ _1497_ _0495_ _2223_ vssd1 vssd1 vccd1 vccd1 _2224_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4702_ _0578_ _3218_ _0574_ _3221_ vssd1 vssd1 vccd1 vccd1 _1183_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5682_ _3053_ _3197_ _0607_ _3200_ _2154_ vssd1 vssd1 vccd1 vccd1 _2155_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _0442_ _0703_ vssd1 vssd1 vccd1 vccd1 _1115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4564_ _1033_ _1037_ _1041_ _1045_ vssd1 vssd1 vccd1 vccd1 _1046_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6303_ net18 net17 vssd1 vssd1 vccd1 vccd1 _2646_ sky130_fd_sc_hd__nand2_1
X_3515_ net8 _3050_ _3006_ vssd1 vssd1 vccd1 vccd1 _3051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4495_ _0403_ _0701_ vssd1 vssd1 vccd1 vccd1 _0978_ sky130_fd_sc_hd__nand2_1
X_6685__15 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__inv_2
X_6234_ _2603_ _2601_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[5\] sky130_fd_sc_hd__nor2_2
XFILLER_0_12_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3446_ _2996_ vssd1 vssd1 vccd1 vccd1 _2997_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _2932_ vssd1 vssd1 vccd1 vccd1 _2554_ sky130_fd_sc_hd__clkbuf_4
X_3377_ _2934_ vssd1 vssd1 vccd1 vccd1 _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5116_ _0352_ egd_top.BitStream_buffer.BS_buffer\[46\] _0355_ _0695_ vssd1 vssd1
+ vccd1 vccd1 _1594_ sky130_fd_sc_hd__a22o_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _2506_ _2502_ vssd1 vssd1 vccd1 vccd1 _2507_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5047_ _1517_ _1521_ _1523_ _1525_ vssd1 vssd1 vccd1 vccd1 _1526_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5949_ _2405_ vssd1 vssd1 vccd1 vccd1 _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ _3069_ vssd1 vssd1 vccd1 vccd1 _0764_ sky130_fd_sc_hd__inv_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6852_ net50 _0255_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_5803_ _0750_ _3217_ _0559_ _3220_ vssd1 vssd1 vccd1 vccd1 _2275_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3995_ _0480_ vssd1 vssd1 vccd1 vccd1 _0481_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6783_ net137 _0186_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[109\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5734_ _0415_ _3136_ vssd1 vssd1 vccd1 vccd1 _2207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5665_ _3149_ _3100_ _3255_ _3105_ _2137_ vssd1 vssd1 vccd1 vccd1 _2138_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4616_ _1096_ _1097_ vssd1 vssd1 vccd1 vccd1 _1098_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5596_ _0333_ _0703_ vssd1 vssd1 vccd1 vccd1 _2070_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4547_ _1029_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1030_ sky130_fd_sc_hd__a21oi_1
X_4478_ _0915_ _0929_ _0943_ _0960_ vssd1 vssd1 vccd1 vccd1 _0961_ sky130_fd_sc_hd__and4_1
X_6217_ _2589_ _2581_ vssd1 vssd1 vccd1 vccd1 _2590_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3429_ egd_top.BitStream_buffer.pc_previous\[6\] _2965_ vssd1 vssd1 vccd1 vccd1 _2983_
+ sky130_fd_sc_hd__or2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _2542_ vssd1 vssd1 vccd1 vccd1 _0206_ sky130_fd_sc_hd__clkbuf_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ net3 _0404_ _2486_ vssd1 vssd1 vccd1 vccd1 _2495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3780_ egd_top.BitStream_buffer.BS_buffer\[104\] vssd1 vssd1 vccd1 vccd1 _3314_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5450_ _3254_ _3232_ vssd1 vssd1 vccd1 vccd1 _1925_ sky130_fd_sc_hd__nand2_1
X_4401_ _0566_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _0885_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5381_ _0460_ _3076_ vssd1 vssd1 vccd1 vccd1 _1857_ sky130_fd_sc_hd__nand2_1
X_4332_ _3330_ _3341_ vssd1 vssd1 vccd1 vccd1 _0816_ sky130_fd_sc_hd__nand2_1
X_4263_ _0563_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _0748_
+ sky130_fd_sc_hd__nand2_1
X_6002_ _2441_ _2423_ vssd1 vssd1 vccd1 vccd1 _2442_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4194_ _0663_ _0667_ _0673_ _0678_ vssd1 vssd1 vccd1 vccd1 _0679_ sky130_fd_sc_hd__and4_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6904_ net102 _0307_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[118\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6835_ net189 _0238_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[41\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3978_ _0447_ _0450_ _0451_ _0454_ _0463_ vssd1 vssd1 vccd1 vccd1 _0464_ sky130_fd_sc_hd__a221oi_1
X_6766_ net120 _0169_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[87\]
+ sky130_fd_sc_hd__dfxtp_1
X_5717_ _0337_ _0703_ vssd1 vssd1 vccd1 vccd1 _2190_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5648_ _0516_ _0569_ vssd1 vssd1 vccd1 vccd1 _2122_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5579_ _3308_ _3022_ vssd1 vssd1 vccd1 vccd1 _2053_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6590__83 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__2927_ clknet_0__2927_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2927_
+ sky130_fd_sc_hd__clkbuf_16
Xinput8 la_data_in_58_43[1] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4950_ _0780_ _3204_ _1428_ vssd1 vssd1 vccd1 vccd1 _1429_ sky130_fd_sc_hd__o21ai_1
X_3901_ _3145_ _0325_ vssd1 vssd1 vccd1 vccd1 _0387_ sky130_fd_sc_hd__and2_1
X_4881_ _0416_ _0461_ vssd1 vssd1 vccd1 vccd1 _1361_ sky130_fd_sc_hd__nand2_1
X_3832_ _3365_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _3366_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6551_ _2884_ vssd1 vssd1 vccd1 vccd1 _2885_ sky130_fd_sc_hd__inv_2
X_3763_ egd_top.BitStream_buffer.BS_buffer\[106\] vssd1 vssd1 vccd1 vccd1 _3297_ sky130_fd_sc_hd__clkbuf_4
X_5502_ _0611_ _0458_ _1976_ vssd1 vssd1 vccd1 vccd1 _1977_ sky130_fd_sc_hd__o21ai_1
X_6482_ _2820_ _2822_ vssd1 vssd1 vccd1 vccd1 egd_top.exp_golomb_decoding.te_range\[2\]
+ sky130_fd_sc_hd__nor2_1
X_3694_ _3227_ vssd1 vssd1 vccd1 vccd1 _3228_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5433_ _0804_ _3148_ _3225_ _3152_ _1907_ vssd1 vssd1 vccd1 vccd1 _1908_ sky130_fd_sc_hd__a221oi_1
X_5364_ _1470_ _0369_ _1839_ vssd1 vssd1 vccd1 vccd1 _1840_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4315_ _3254_ _3259_ vssd1 vssd1 vccd1 vccd1 _0799_ sky130_fd_sc_hd__nand2_1
X_5295_ _0606_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _1772_
+ sky130_fd_sc_hd__nand2_1
X_4246_ _0489_ _0488_ _0493_ _0492_ _0730_ vssd1 vssd1 vccd1 vccd1 _0731_ sky130_fd_sc_hd__a221oi_1
X_4177_ _0660_ _0661_ vssd1 vssd1 vccd1 vccd1 _0662_ sky130_fd_sc_hd__nand2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6818_ net172 _0221_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[58\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _0940_ _3238_ _1069_ _3241_ vssd1 vssd1 vccd1 vccd1 _1558_ sky130_fd_sc_hd__o22ai_1
X_4100_ _0574_ _0576_ _0578_ _0580_ _0585_ vssd1 vssd1 vccd1 vccd1 _0586_ sky130_fd_sc_hd__o221a_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4031_ _3139_ _0470_ vssd1 vssd1 vccd1 vccd1 _0517_ sky130_fd_sc_hd__nand2_1
X_5982_ _2428_ vssd1 vssd1 vccd1 vccd1 _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4933_ _3120_ _3111_ _1411_ vssd1 vssd1 vccd1 vccd1 _1412_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4864_ _1342_ _1343_ vssd1 vssd1 vccd1 vccd1 _1344_ sky130_fd_sc_hd__nand2_1
XANTENNA_13 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4795_ _1150_ _0595_ _0494_ _0598_ vssd1 vssd1 vccd1 vccd1 _1276_ sky130_fd_sc_hd__o22ai_1
X_3815_ _3139_ _3299_ vssd1 vssd1 vccd1 vccd1 _3349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6534_ _2867_ vssd1 vssd1 vccd1 vccd1 _2869_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3746_ _3279_ vssd1 vssd1 vccd1 vccd1 _3280_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6465_ _2805_ vssd1 vssd1 vccd1 vccd1 _2806_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5416_ _0606_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _1892_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3677_ _3210_ vssd1 vssd1 vccd1 vccd1 _3211_ sky130_fd_sc_hd__buf_1
X_6396_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2739_ sky130_fd_sc_hd__xnor2_1
X_5347_ _3340_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _1823_
+ sky130_fd_sc_hd__nand2_1
X_5278_ _1753_ _1754_ vssd1 vssd1 vccd1 vccd1 _1755_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4229_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _0714_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 la_data_in_58_43[4] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_8
X_4580_ _3250_ _3275_ vssd1 vssd1 vccd1 vccd1 _1062_ sky130_fd_sc_hd__nand2_1
X_3600_ egd_top.BitStream_buffer.BS_buffer\[70\] vssd1 vssd1 vccd1 vccd1 _3134_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3531_ _3064_ vssd1 vssd1 vccd1 vccd1 _3065_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6250_ _2610_ vssd1 vssd1 vccd1 vccd1 _0178_ sky130_fd_sc_hd__inv_2
X_3462_ net6 _3010_ _3007_ vssd1 vssd1 vccd1 vccd1 _3011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6181_ _2565_ vssd1 vssd1 vccd1 vccd1 _0196_ sky130_fd_sc_hd__clkbuf_1
X_3393_ _2947_ vssd1 vssd1 vccd1 vccd1 _0318_ sky130_fd_sc_hd__inv_2
X_5201_ egd_top.BitStream_buffer.BS_buffer\[7\] _3212_ egd_top.BitStream_buffer.BS_buffer\[8\]
+ _3215_ _1677_ vssd1 vssd1 vccd1 vccd1 _1678_ sky130_fd_sc_hd__a221oi_1
X_5132_ _0903_ _0414_ _1607_ _1608_ _1609_ vssd1 vssd1 vccd1 vccd1 _1610_ sky130_fd_sc_hd__o2111a_1
X_5063_ _1284_ _3124_ _1538_ _1539_ _1540_ vssd1 vssd1 vccd1 vccd1 _1541_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4014_ _0498_ _0499_ vssd1 vssd1 vccd1 vccd1 _0500_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6606__98 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__inv_2
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5965_ _2416_ _2396_ vssd1 vssd1 vccd1 vccd1 _2417_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5896_ _0605_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _2368_
+ sky130_fd_sc_hd__nand2_1
X_4916_ _0890_ _0570_ vssd1 vssd1 vccd1 vccd1 _1396_ sky130_fd_sc_hd__or2_1
X_4847_ _2998_ _3303_ _3010_ _3307_ _1326_ vssd1 vssd1 vccd1 vccd1 _1327_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _0862_ _0518_ vssd1 vssd1 vccd1 vccd1 _1259_ sky130_fd_sc_hd__or2_1
X_6517_ _2813_ _2852_ vssd1 vssd1 vccd1 vccd1 _2853_ sky130_fd_sc_hd__nand2_1
X_3729_ _3126_ _3228_ vssd1 vssd1 vccd1 vccd1 _3263_ sky130_fd_sc_hd__nand2_2
X_6448_ _2758_ _2760_ _2789_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__o21ai_2
X_6379_ _2707_ egd_top.BitStream_buffer.BitStream_buffer_output\[1\] vssd1 vssd1 vccd1
+ vccd1 _2722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5750_ _0497_ _0359_ vssd1 vssd1 vccd1 vccd1 _2223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4701_ _3028_ _3198_ _3031_ _3201_ _1181_ vssd1 vssd1 vccd1 vccd1 _1182_ sky130_fd_sc_hd__a221oi_2
X_5681_ _3219_ _3203_ _2153_ vssd1 vssd1 vccd1 vccd1 _2154_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4632_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _1114_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6672__159 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__inv_2
X_4563_ _3259_ _3148_ _3251_ _3152_ _1044_ vssd1 vssd1 vccd1 vccd1 _1045_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4494_ _0399_ _0423_ vssd1 vssd1 vccd1 vccd1 _0977_ sky130_fd_sc_hd__nand2_1
X_6302_ _2645_ vssd1 vssd1 vccd1 vccd1 _0161_ sky130_fd_sc_hd__clkbuf_1
X_3514_ egd_top.BitStream_buffer.BS_buffer\[126\] vssd1 vssd1 vccd1 vccd1 _3050_ sky130_fd_sc_hd__clkbuf_4
X_6233_ _2600_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2603_ sky130_fd_sc_hd__a21oi_1
X_3445_ egd_top.BitStream_buffer.BitStream_buffer_valid_n vssd1 vssd1 vccd1 vccd1
+ _2996_ sky130_fd_sc_hd__buf_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _2931_ _2933_ vssd1 vssd1 vccd1 vccd1 _2934_ sky130_fd_sc_hd__and2_1
X_6164_ net1 _3149_ _2520_ vssd1 vssd1 vccd1 vccd1 _2553_ sky130_fd_sc_hd__mux2_1
X_5115_ _1470_ _0345_ _1592_ _0349_ vssd1 vssd1 vccd1 vccd1 _1593_ sky130_fd_sc_hd__o22ai_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ net13 _0423_ _2486_ vssd1 vssd1 vccd1 vccd1 _2506_ sky130_fd_sc_hd__mux2_1
X_5046_ _0515_ _0589_ _0509_ _0592_ _1524_ vssd1 vssd1 vccd1 vccd1 _1525_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5948_ _2404_ _2396_ vssd1 vssd1 vccd1 vccd1 _2405_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5879_ _2349_ _2350_ vssd1 vssd1 vccd1 vccd1 _2351_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6851_ net49 _0254_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[25\]
+ sky130_fd_sc_hd__dfxtp_1
X_5802_ _0607_ _3197_ _0577_ _3200_ _2273_ vssd1 vssd1 vccd1 vccd1 _2274_ sky130_fd_sc_hd__a221oi_1
X_3994_ _3072_ _0469_ vssd1 vssd1 vccd1 vccd1 _0480_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6782_ net136 _0185_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[110\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5733_ _0767_ _0396_ _2203_ _2204_ _2205_ vssd1 vssd1 vccd1 vccd1 _2206_ sky130_fd_sc_hd__o2111a_1
X_5664_ _1031_ _3110_ _2136_ vssd1 vssd1 vccd1 vccd1 _2137_ sky130_fd_sc_hd__o21ai_1
X_4615_ _0352_ egd_top.BitStream_buffer.BS_buffer\[42\] _0355_ _0329_ vssd1 vssd1
+ vccd1 vccd1 _1097_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5595_ _2028_ _2039_ _2052_ _2068_ vssd1 vssd1 vccd1 vccd1 _2069_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4546_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1 vccd1 vccd1
+ _1029_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4477_ _0947_ _0951_ _0956_ _0959_ vssd1 vssd1 vccd1 vccd1 _0960_ sky130_fd_sc_hd__and4_1
X_6216_ net1 _0675_ net197 vssd1 vssd1 vccd1 vccd1 _2589_ sky130_fd_sc_hd__mux2_1
X_3428_ _2968_ _2981_ vssd1 vssd1 vccd1 vccd1 _2982_ sky130_fd_sc_hd__nand2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6609__101 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__inv_2
X_6147_ _2541_ _2529_ vssd1 vssd1 vccd1 vccd1 _2542_ sky130_fd_sc_hd__and2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ _2494_ vssd1 vssd1 vccd1 vccd1 _0228_ sky130_fd_sc_hd__clkbuf_1
X_5029_ _1373_ _0506_ _1505_ _1506_ _1507_ vssd1 vssd1 vccd1 vccd1 _1508_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6655__143 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__inv_2
XFILLER_0_35_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6742__67 clknet_1_1__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__inv_2
X_4400_ _0563_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _0884_
+ sky130_fd_sc_hd__nand2_1
X_5380_ _0447_ _0432_ _0451_ _0436_ _1855_ vssd1 vssd1 vccd1 vccd1 _1856_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4331_ _3326_ _3347_ vssd1 vssd1 vccd1 vccd1 _0815_ sky130_fd_sc_hd__nand2_1
X_4262_ _0742_ _0545_ _0743_ _0744_ _0746_ vssd1 vssd1 vccd1 vccd1 _0747_ sky130_fd_sc_hd__o2111a_1
X_6001_ net10 _0535_ _2414_ vssd1 vssd1 vccd1 vccd1 _2441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4193_ _3357_ _3356_ _0674_ _3360_ _0677_ vssd1 vssd1 vccd1 vccd1 _0678_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6903_ net101 _0306_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[119\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6834_ net188 _0237_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[42\]
+ sky130_fd_sc_hd__dfxtp_1
X_3977_ _0456_ _0458_ _0462_ vssd1 vssd1 vccd1 vccd1 _0463_ sky130_fd_sc_hd__o21ai_1
X_6765_ net119 _0168_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[88\]
+ sky130_fd_sc_hd__dfxtp_1
X_5716_ _0333_ _0400_ vssd1 vssd1 vccd1 vccd1 _2189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5647_ _0565_ _0513_ vssd1 vssd1 vccd1 vccd1 _2121_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5578_ _2041_ _2046_ _2049_ _2051_ vssd1 vssd1 vccd1 vccd1 _2052_ sky130_fd_sc_hd__and4_1
X_4529_ _0547_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _1012_
+ sky130_fd_sc_hd__nand2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__2926_ clknet_0__2926_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2926_
+ sky130_fd_sc_hd__clkbuf_16
Xinput9 la_data_in_58_43[2] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3900_ _0385_ vssd1 vssd1 vccd1 vccd1 _0386_ sky130_fd_sc_hd__clkbuf_4
X_4880_ _0412_ _0397_ _1357_ _1358_ _1359_ vssd1 vssd1 vccd1 vccd1 _1360_ sky130_fd_sc_hd__o2111a_1
X_3831_ _3364_ vssd1 vssd1 vccd1 vccd1 _3365_ sky130_fd_sc_hd__clkbuf_4
X_6550_ _2716_ _2883_ vssd1 vssd1 vccd1 vccd1 _2884_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3762_ _3243_ _3261_ _3277_ _3295_ vssd1 vssd1 vccd1 vccd1 _3296_ sky130_fd_sc_hd__and4_1
X_5501_ _0460_ _3085_ vssd1 vssd1 vccd1 vccd1 _1976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6481_ _2821_ _2647_ vssd1 vssd1 vccd1 vccd1 _2822_ sky130_fd_sc_hd__nand2_1
X_3693_ _3226_ vssd1 vssd1 vccd1 vccd1 _3227_ sky130_fd_sc_hd__inv_2
X_5432_ _1905_ _1906_ vssd1 vssd1 vccd1 vccd1 _1907_ sky130_fd_sc_hd__nand2_1
X_5363_ _0371_ _0380_ vssd1 vssd1 vccd1 vccd1 _1839_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _3250_ _3265_ vssd1 vssd1 vccd1 vccd1 _0798_ sky130_fd_sc_hd__nand2_1
X_5294_ _1740_ _1757_ _1770_ vssd1 vssd1 vccd1 vccd1 _1771_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4245_ _0728_ _0496_ _0729_ vssd1 vssd1 vccd1 vccd1 _0730_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4176_ _3313_ _3310_ vssd1 vssd1 vccd1 vccd1 _0661_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6817_ net171 _0220_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[59\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6706__34 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__inv_2
X_6721__48 clknet_1_0__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__inv_2
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4030_ _0515_ vssd1 vssd1 vccd1 vccd1 _0516_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5981_ _2427_ _2423_ vssd1 vssd1 vccd1 vccd1 _2428_ sky130_fd_sc_hd__and2_1
X_4932_ _3114_ _3076_ vssd1 vssd1 vccd1 vccd1 _1411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _0338_ _0389_ vssd1 vssd1 vccd1 vccd1 _1343_ sky130_fd_sc_hd__nand2_1
XANTENNA_14 net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _3347_ vssd1 vssd1 vccd1 vccd1 _3348_ sky130_fd_sc_hd__inv_2
X_4794_ _0554_ _0576_ _0742_ _0580_ _1274_ vssd1 vssd1 vccd1 vccd1 _1275_ sky130_fd_sc_hd__o221a_1
X_6533_ _2856_ _2867_ vssd1 vssd1 vccd1 vccd1 _2868_ sky130_fd_sc_hd__nand2_1
X_3745_ _3145_ _3227_ vssd1 vssd1 vccd1 vccd1 _3279_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6464_ _2661_ _2745_ vssd1 vssd1 vccd1 vccd1 _2805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5415_ _1861_ _1877_ _1890_ vssd1 vssd1 vccd1 vccd1 _1891_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3676_ _3145_ _3166_ vssd1 vssd1 vccd1 vccd1 _3210_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6395_ _2733_ _2737_ vssd1 vssd1 vccd1 vccd1 _2738_ sky130_fd_sc_hd__nand2_1
X_5346_ _3297_ _3321_ _3304_ _3324_ _1821_ vssd1 vssd1 vccd1 vccd1 _1822_ sky130_fd_sc_hd__a221oi_1
X_5277_ _0534_ _0346_ vssd1 vssd1 vccd1 vccd1 _1754_ sky130_fd_sc_hd__nand2_1
X_4228_ _0708_ _0414_ _0709_ _0710_ _0712_ vssd1 vssd1 vccd1 vccd1 _0713_ sky130_fd_sc_hd__o2111a_1
X_4159_ _3232_ _3231_ _3286_ _3235_ _0643_ vssd1 vssd1 vccd1 vccd1 _0644_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_65_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 la_data_in_58_43[5] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3530_ _3062_ _3063_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _3064_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3461_ egd_top.BitStream_buffer.BS_buffer\[113\] vssd1 vssd1 vccd1 vccd1 _3010_ sky130_fd_sc_hd__clkbuf_4
X_3392_ _2937_ _2942_ _2946_ vssd1 vssd1 vccd1 vccd1 _2947_ sky130_fd_sc_hd__or3_1
X_6180_ _2564_ _2554_ vssd1 vssd1 vccd1 vccd1 _2565_ sky130_fd_sc_hd__and2_1
X_5200_ _0541_ _3218_ _0742_ _3221_ vssd1 vssd1 vccd1 vccd1 _1677_ sky130_fd_sc_hd__o22ai_1
X_6700__29 clknet_1_0__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__inv_2
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5131_ _0614_ _0426_ vssd1 vssd1 vccd1 vccd1 _1609_ sky130_fd_sc_hd__or2_1
X_5062_ _1031_ _3141_ vssd1 vssd1 vccd1 vccd1 _1540_ sky130_fd_sc_hd__or2_1
X_4013_ egd_top.BitStream_buffer.BS_buffer\[19\] vssd1 vssd1 vccd1 vccd1 _0499_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5964_ net7 egd_top.BitStream_buffer.BS_buffer\[16\] _2415_ vssd1 vssd1 vccd1 vccd1
+ _2416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5895_ _2337_ _2353_ _2366_ vssd1 vssd1 vccd1 vccd1 _2367_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4915_ _0566_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1395_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4846_ _1324_ _1325_ vssd1 vssd1 vccd1 vccd1 _1326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4777_ _0512_ _0475_ vssd1 vssd1 vccd1 vccd1 _1258_ sky130_fd_sc_hd__nand2_1
X_6516_ _2760_ vssd1 vssd1 vccd1 vccd1 _2852_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3728_ egd_top.BitStream_buffer.BS_buffer\[84\] vssd1 vssd1 vccd1 vccd1 _3262_ sky130_fd_sc_hd__inv_2
X_6447_ _2787_ _2788_ _2756_ vssd1 vssd1 vccd1 vccd1 _2789_ sky130_fd_sc_hd__nand3_1
X_3659_ _3192_ _3037_ vssd1 vssd1 vccd1 vccd1 _3193_ sky130_fd_sc_hd__nand2_1
X_6378_ _2720_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2721_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5329_ _3250_ _3290_ vssd1 vssd1 vccd1 vccd1 _1805_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4700_ _3177_ _3204_ _1180_ vssd1 vssd1 vccd1 vccd1 _1181_ sky130_fd_sc_hd__o21ai_1
X_5680_ _3205_ _3050_ vssd1 vssd1 vccd1 vccd1 _2153_ sky130_fd_sc_hd__nand2_1
X_4631_ _0456_ _0414_ _1110_ _1111_ _1112_ vssd1 vssd1 vccd1 vccd1 _1113_ sky130_fd_sc_hd__o2111a_1
X_4562_ _1042_ _1043_ vssd1 vssd1 vccd1 vccd1 _1044_ sky130_fd_sc_hd__nand2_1
X_4493_ _0965_ _0969_ _0972_ _0975_ vssd1 vssd1 vccd1 vccd1 _0976_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6301_ _2644_ _2372_ vssd1 vssd1 vccd1 vccd1 _2645_ sky130_fd_sc_hd__and2_1
X_3513_ _3049_ vssd1 vssd1 vccd1 vccd1 _0300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3444_ _2994_ _2995_ _2938_ vssd1 vssd1 vccd1 vccd1 _0315_ sky130_fd_sc_hd__a21oi_1
X_6232_ _2602_ vssd1 vssd1 vccd1 vccd1 _0183_ sky130_fd_sc_hd__inv_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _2932_ vssd1 vssd1 vccd1 vccd1 _2933_ sky130_fd_sc_hd__buf_2
X_6163_ _2552_ vssd1 vssd1 vccd1 vccd1 _0201_ sky130_fd_sc_hd__clkbuf_1
X_5114_ egd_top.BitStream_buffer.BS_buffer\[45\] vssd1 vssd1 vccd1 vccd1 _1592_ sky130_fd_sc_hd__inv_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _2505_ vssd1 vssd1 vccd1 vccd1 _0223_ sky130_fd_sc_hd__clkbuf_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _0728_ _0595_ _0867_ _0598_ vssd1 vssd1 vccd1 vccd1 _1524_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5947_ net11 egd_top.BitStream_buffer.BS_buffer\[11\] _2380_ vssd1 vssd1 vccd1 vccd1
+ _2404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6748__73 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__inv_2
XFILLER_0_90_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5878_ _0533_ _0323_ vssd1 vssd1 vccd1 vccd1 _2350_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4829_ _1300_ _1303_ _1306_ _1308_ vssd1 vssd1 vccd1 vccd1 _1309_ sky130_fd_sc_hd__and4_1
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6632__122 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__inv_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net202 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_1
X_6850_ net48 _0253_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6781_ net135 _0184_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[111\]
+ sky130_fd_sc_hd__dfxtp_1
X_5801_ _0638_ _3203_ _2272_ vssd1 vssd1 vccd1 vccd1 _2273_ sky130_fd_sc_hd__o21ai_1
X_3993_ egd_top.BitStream_buffer.BS_buffer\[26\] vssd1 vssd1 vccd1 vccd1 _0479_ sky130_fd_sc_hd__clkbuf_4
X_5732_ _1034_ _0407_ vssd1 vssd1 vccd1 vccd1 _2205_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5663_ _3113_ _3144_ vssd1 vssd1 vccd1 vccd1 _2136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4614_ _0966_ _0345_ _1095_ _0349_ vssd1 vssd1 vccd1 vccd1 _1096_ sky130_fd_sc_hd__o22ai_1
X_5594_ _2056_ _2060_ _2064_ _2067_ vssd1 vssd1 vccd1 vccd1 _2068_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4545_ _0961_ _1026_ _1027_ vssd1 vssd1 vccd1 vccd1 _1028_ sky130_fd_sc_hd__nand3_1
X_4476_ _0675_ _3356_ _2998_ _3360_ _0958_ vssd1 vssd1 vccd1 vccd1 _0959_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_0_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6215_ _2588_ vssd1 vssd1 vccd1 vccd1 _0185_ sky130_fd_sc_hd__clkbuf_1
X_3427_ _2980_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ egd_top.BitStream_buffer.pc_previous\[6\] vssd1 vssd1 vccd1 vccd1 _2981_ sky130_fd_sc_hd__a31o_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ net13 _3085_ _2521_ vssd1 vssd1 vccd1 vccd1 _2541_ sky130_fd_sc_hd__mux2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ _2493_ _2475_ vssd1 vssd1 vccd1 vccd1 _2494_ sky130_fd_sc_hd__and2_1
X_5028_ _1123_ _0518_ vssd1 vssd1 vccd1 vccd1 _1507_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4330_ _3353_ _3303_ _3357_ _3307_ _0813_ vssd1 vssd1 vccd1 vccd1 _0814_ sky130_fd_sc_hd__a221oi_1
X_4261_ _0745_ _0556_ vssd1 vssd1 vccd1 vccd1 _0746_ sky130_fd_sc_hd__or2_1
X_6000_ _2440_ vssd1 vssd1 vccd1 vccd1 _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4192_ _3202_ _3363_ _0676_ vssd1 vssd1 vccd1 vccd1 _0677_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6902_ net100 _0305_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[120\]
+ sky130_fd_sc_hd__dfxtp_1
X_6833_ net187 _0236_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[43\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3976_ _0460_ _0461_ vssd1 vssd1 vccd1 vccd1 _0462_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6764_ net118 _0167_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[89\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6639__128 clknet_1_0__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__inv_2
X_5715_ _2147_ _2158_ _2171_ _2187_ vssd1 vssd1 vccd1 vccd1 _2188_ sky130_fd_sc_hd__and4_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5646_ _0562_ _0509_ vssd1 vssd1 vccd1 vccd1 _2120_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5577_ _3297_ _3280_ _3304_ _3284_ _2050_ vssd1 vssd1 vccd1 vccd1 _2051_ sky130_fd_sc_hd__a221oi_1
X_4528_ _0999_ _1002_ _1006_ _1010_ vssd1 vssd1 vccd1 vccd1 _1011_ sky130_fd_sc_hd__and4_1
X_4459_ _3322_ _3281_ _3331_ _3285_ _0941_ vssd1 vssd1 vccd1 vccd1 _0942_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ _2528_ _2529_ vssd1 vssd1 vccd1 vccd1 _2530_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2925_ clknet_0__2925_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2925_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ _3145_ _3300_ vssd1 vssd1 vccd1 vccd1 _3364_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3761_ _3278_ _3281_ _3282_ _3285_ _3294_ vssd1 vssd1 vccd1 vccd1 _3295_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5500_ _0451_ _0432_ _0461_ _0436_ _1974_ vssd1 vssd1 vccd1 vccd1 _1975_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_6_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6480_ _2817_ _2819_ _2818_ vssd1 vssd1 vccd1 vccd1 _2821_ sky130_fd_sc_hd__nand3_1
X_3692_ egd_top.BitStream_buffer.pc\[5\] _2965_ _3062_ vssd1 vssd1 vccd1 vccd1 _3226_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5431_ _3160_ _3275_ vssd1 vssd1 vccd1 vccd1 _1906_ sky130_fd_sc_hd__nand2_1
X_5362_ _1836_ _1837_ vssd1 vssd1 vccd1 vccd1 _1838_ sky130_fd_sc_hd__nor2_1
X_4313_ _3246_ _3251_ vssd1 vssd1 vccd1 vccd1 _0797_ sky130_fd_sc_hd__nand2_1
X_5293_ _1761_ _1765_ _1767_ _1769_ vssd1 vssd1 vccd1 vccd1 _1770_ sky130_fd_sc_hd__and4_1
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4244_ _0498_ _0513_ vssd1 vssd1 vccd1 vccd1 _0729_ sky130_fd_sc_hd__nand2_1
X_4175_ _3309_ _3297_ vssd1 vssd1 vccd1 vccd1 _0660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6816_ net170 _0219_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[60\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3959_ _0438_ _0440_ _0444_ vssd1 vssd1 vccd1 vccd1 _0445_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5629_ _0343_ _0471_ _2100_ _2102_ vssd1 vssd1 vccd1 vccd1 _2103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6757__5 clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__inv_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ net2 _0515_ _2415_ vssd1 vssd1 vccd1 vccd1 _2427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4931_ _3247_ _3068_ _3259_ _3075_ _1409_ vssd1 vssd1 vccd1 vccd1 _1410_ sky130_fd_sc_hd__a221oi_1
X_4862_ _0334_ _0695_ vssd1 vssd1 vccd1 vccd1 _1342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3813_ egd_top.BitStream_buffer.BS_buffer\[101\] vssd1 vssd1 vccd1 vccd1 _3347_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 _1447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _0745_ _0584_ vssd1 vssd1 vccd1 vccd1 _1274_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6532_ _2866_ _2959_ vssd1 vssd1 vccd1 vccd1 _2867_ sky130_fd_sc_hd__nand2_1
X_3744_ egd_top.BitStream_buffer.BS_buffer\[94\] vssd1 vssd1 vccd1 vccd1 _3278_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3675_ _3013_ _3198_ _3016_ _3201_ _3208_ vssd1 vssd1 vccd1 vccd1 _3209_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6463_ _1530_ _2662_ vssd1 vssd1 vccd1 vccd1 _2804_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5414_ _1881_ _1885_ _1887_ _1889_ vssd1 vssd1 vccd1 vccd1 _1890_ sky130_fd_sc_hd__and4_1
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6394_ _2735_ _2736_ vssd1 vssd1 vccd1 vccd1 _2737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5345_ _1819_ _1820_ vssd1 vssd1 vccd1 vccd1 _1821_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5276_ _0530_ _0353_ vssd1 vssd1 vccd1 vccd1 _1753_ sky130_fd_sc_hd__nand2_1
X_4227_ _0711_ _0426_ vssd1 vssd1 vccd1 vccd1 _0712_ sky130_fd_sc_hd__or2_1
X_4158_ _3239_ _3238_ _0642_ _3241_ vssd1 vssd1 vccd1 vccd1 _0643_ sky130_fd_sc_hd__o22ai_1
X_4089_ _3098_ _0543_ vssd1 vssd1 vccd1 vccd1 _0575_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__2927_ _2927_ vssd1 vssd1 vccd1 vccd1 clknet_0__2927_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_439 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput13 la_data_in_58_43[6] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6697__26 clknet_1_0__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__inv_2
X_3460_ _3009_ vssd1 vssd1 vccd1 vccd1 _0313_ sky130_fd_sc_hd__clkbuf_1
X_3391_ net31 _2945_ vssd1 vssd1 vccd1 vccd1 _2946_ sky130_fd_sc_hd__nor2_1
X_5130_ _0420_ _3095_ vssd1 vssd1 vccd1 vccd1 _1608_ sky130_fd_sc_hd__nand2_1
X_5061_ _3133_ _3144_ vssd1 vssd1 vccd1 vccd1 _1539_ sky130_fd_sc_hd__nand2_1
X_4012_ _0497_ vssd1 vssd1 vccd1 vccd1 _0498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5963_ _2414_ vssd1 vssd1 vccd1 vccd1 _2415_ sky130_fd_sc_hd__buf_4
XFILLER_0_59_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4914_ _0563_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1394_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5894_ _2357_ _2361_ _2363_ _2365_ vssd1 vssd1 vccd1 vccd1 _2366_ sky130_fd_sc_hd__and4_1
X_4845_ _3313_ _0674_ vssd1 vssd1 vccd1 vccd1 _1325_ sky130_fd_sc_hd__nand2_1
X_4776_ _0508_ _0482_ vssd1 vssd1 vccd1 vccd1 _1257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6515_ _2850_ _2756_ vssd1 vssd1 vccd1 vccd1 _2851_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3727_ _3248_ _3252_ _3256_ _3260_ vssd1 vssd1 vccd1 vccd1 _3261_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6446_ _2786_ _2758_ vssd1 vssd1 vccd1 vccd1 _2788_ sky130_fd_sc_hd__nand2_2
X_3658_ _3191_ vssd1 vssd1 vccd1 vccd1 _3192_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6377_ _2701_ _2668_ vssd1 vssd1 vccd1 vccd1 _2720_ sky130_fd_sc_hd__nand2_1
X_3589_ _3122_ _3065_ vssd1 vssd1 vccd1 vccd1 _3123_ sky130_fd_sc_hd__nand2_1
X_5328_ _3246_ _3232_ vssd1 vssd1 vccd1 vccd1 _1804_ sky130_fd_sc_hd__nand2_1
X_5259_ _0460_ _3119_ vssd1 vssd1 vccd1 vccd1 _1736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4630_ _0848_ _0426_ vssd1 vssd1 vccd1 vccd1 _1112_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6300_ net1 _3282_ net199 vssd1 vssd1 vccd1 vccd1 _2644_ sky130_fd_sc_hd__mux2_1
X_4561_ _3160_ _3255_ vssd1 vssd1 vccd1 vccd1 _1043_ sky130_fd_sc_hd__nand2_1
X_4492_ _0695_ _0379_ _0437_ _0383_ _0974_ vssd1 vssd1 vccd1 vccd1 _0975_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3512_ _3048_ _3042_ vssd1 vssd1 vccd1 vccd1 _3049_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3443_ _2988_ net28 vssd1 vssd1 vccd1 vccd1 _2995_ sky130_fd_sc_hd__nand2_1
X_6231_ _2989_ egd_top.BitStream_buffer.pc\[6\] vssd1 vssd1 vccd1 vccd1 _2602_ sky130_fd_sc_hd__nand2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _2551_ _2529_ vssd1 vssd1 vccd1 vccd1 _2552_ sky130_fd_sc_hd__and2_1
X_5113_ _0429_ _0328_ _0433_ _0332_ _1590_ vssd1 vssd1 vccd1 vccd1 _1591_ sky130_fd_sc_hd__a221oi_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ net19 vssd1 vssd1 vccd1 vccd1 _2932_ sky130_fd_sc_hd__buf_6
XFILLER_0_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ _2504_ _2502_ vssd1 vssd1 vccd1 vccd1 _2505_ sky130_fd_sc_hd__and2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _0568_ _0576_ _0745_ _0580_ _1522_ vssd1 vssd1 vccd1 vccd1 _1523_ sky130_fd_sc_hd__o221a_1
XFILLER_0_18_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5946_ _2403_ vssd1 vssd1 vccd1 vccd1 _0269_ sky130_fd_sc_hd__clkbuf_1
X_5877_ _0529_ _0329_ vssd1 vssd1 vccd1 vccd1 _2349_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4828_ _0552_ _3212_ _0540_ _3215_ _1307_ vssd1 vssd1 vccd1 vccd1 _1308_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4759_ _3108_ _0414_ _1237_ _1238_ _1239_ vssd1 vssd1 vccd1 vccd1 _1240_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6429_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] _2735_ vssd1 vssd1
+ vccd1 vccd1 _2771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold2 _2556_ vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3992_ _0477_ vssd1 vssd1 vccd1 vccd1 _0478_ sky130_fd_sc_hd__clkbuf_4
X_6780_ net134 _0183_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[6\]
+ sky130_fd_sc_hd__dfxtp_2
X_5800_ _3205_ _3053_ vssd1 vssd1 vccd1 vccd1 _2272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5731_ _0402_ _3115_ vssd1 vssd1 vccd1 vccd1 _2204_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5662_ _3275_ _3067_ _0653_ _3074_ _2134_ vssd1 vssd1 vccd1 vccd1 _2135_ sky130_fd_sc_hd__a221oi_1
X_4613_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _1095_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5593_ _3031_ _3355_ _3034_ _3359_ _2066_ vssd1 vssd1 vccd1 vccd1 _2067_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4544_ _0606_ _0581_ vssd1 vssd1 vccd1 vccd1 _1027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4475_ _0786_ _3363_ _0957_ vssd1 vssd1 vccd1 vccd1 _0958_ sky130_fd_sc_hd__o21ai_1
X_6214_ _2587_ _2581_ vssd1 vssd1 vccd1 vccd1 _2588_ sky130_fd_sc_hd__and2_1
X_3426_ egd_top.BitStream_buffer.pc_previous\[0\] egd_top.BitStream_buffer.pc_previous\[1\]
+ egd_top.BitStream_buffer.pc_previous\[2\] egd_top.BitStream_buffer.pc_previous\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2980_ sky130_fd_sc_hd__and4_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ _2540_ vssd1 vssd1 vccd1 vccd1 _0207_ sky130_fd_sc_hd__clkbuf_1
X_6076_ net4 _0433_ _2486_ vssd1 vssd1 vccd1 vccd1 _2493_ sky130_fd_sc_hd__mux2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _0512_ _0482_ vssd1 vssd1 vccd1 vccd1 _1506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6587__80 clknet_1_0__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__inv_2
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5929_ _2391_ _3042_ vssd1 vssd1 vccd1 vccd1 _2392_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6616__107 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__inv_2
XFILLER_0_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4260_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0745_ sky130_fd_sc_hd__inv_2
X_4191_ _3365_ _0675_ vssd1 vssd1 vccd1 vccd1 _0676_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6901_ net99 _0304_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[121\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6832_ net186 _0235_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[44\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3975_ egd_top.BitStream_buffer.BS_buffer\[62\] vssd1 vssd1 vccd1 vccd1 _0461_ sky130_fd_sc_hd__clkbuf_4
X_6763_ net117 _0166_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[90\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5714_ _2175_ _2179_ _2183_ _2186_ vssd1 vssd1 vccd1 vccd1 _2187_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5645_ _1150_ _0544_ _2116_ _2117_ _2118_ vssd1 vssd1 vccd1 vccd1 _2119_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5576_ _0668_ _3288_ _0819_ _3292_ vssd1 vssd1 vccd1 vccd1 _2050_ sky130_fd_sc_hd__o22ai_1
X_4527_ _0363_ _0524_ _0689_ _0528_ _1009_ vssd1 vssd1 vccd1 vccd1 _1010_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4458_ _0807_ _3289_ _0940_ _3293_ vssd1 vssd1 vccd1 vccd1 _0941_ sky130_fd_sc_hd__o22ai_1
X_3409_ _2962_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2963_ sky130_fd_sc_hd__nand2_2
X_4389_ _0504_ _0518_ vssd1 vssd1 vccd1 vccd1 _0873_ sky130_fd_sc_hd__or2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6128_ _2932_ vssd1 vssd1 vccd1 vccd1 _2529_ sky130_fd_sc_hd__buf_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ net8 _0389_ net203 vssd1 vssd1 vccd1 vccd1 _2481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__2924_ clknet_0__2924_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2924_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _3287_ _3289_ _3291_ _3293_ vssd1 vssd1 vccd1 vccd1 _3294_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3691_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _3225_ sky130_fd_sc_hd__buf_4
X_5430_ _3155_ _0653_ vssd1 vssd1 vccd1 vccd1 _1905_ sky130_fd_sc_hd__nand2_1
X_5361_ _0352_ _0437_ _0355_ _0443_ vssd1 vssd1 vccd1 vccd1 _1837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _0503_ _0589_ _0467_ _0592_ _1768_ vssd1 vssd1 vccd1 vccd1 _1769_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_10_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4312_ _3286_ _3231_ _3290_ _3235_ _0795_ vssd1 vssd1 vccd1 vccd1 _0796_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4243_ _0499_ vssd1 vssd1 vccd1 vccd1 _0728_ sky130_fd_sc_hd__inv_2
X_4174_ _0644_ _0650_ _0655_ _0658_ vssd1 vssd1 vccd1 vccd1 _0659_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6815_ net169 _0218_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[61\]
+ sky130_fd_sc_hd__dfxtp_1
X_3958_ _0442_ _0443_ vssd1 vssd1 vccd1 vccd1 _0444_ sky130_fd_sc_hd__nand2_1
X_3889_ _0359_ _0362_ _0363_ _0366_ _0374_ vssd1 vssd1 vccd1 vccd1 _0375_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5628_ _2101_ vssd1 vssd1 vccd1 vccd1 _2102_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5559_ _0552_ _3183_ _0540_ _3186_ _2032_ vssd1 vssd1 vccd1 vccd1 _2033_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6668__155 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__inv_2
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4930_ _1284_ _3084_ _1408_ _3092_ vssd1 vssd1 vccd1 vccd1 _1409_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_86_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ _1298_ _1309_ _1323_ _1340_ vssd1 vssd1 vccd1 vccd1 _1341_ sky130_fd_sc_hd__and4_1
XFILLER_0_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3812_ _3344_ _3345_ vssd1 vssd1 vccd1 vccd1 _3346_ sky130_fd_sc_hd__nand2_1
X_4792_ _1022_ _0561_ _1270_ _1271_ _1272_ vssd1 vssd1 vccd1 vccd1 _1273_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6531_ _2863_ _2865_ vssd1 vssd1 vccd1 vccd1 _2866_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3743_ _3269_ _3276_ vssd1 vssd1 vccd1 vccd1 _3277_ sky130_fd_sc_hd__nor2_1
X_3674_ _3202_ _3204_ _3207_ vssd1 vssd1 vccd1 vccd1 _3208_ sky130_fd_sc_hd__o21ai_1
X_6462_ _2733_ _2801_ _2802_ vssd1 vssd1 vccd1 vccd1 _2803_ sky130_fd_sc_hd__and3_1
X_5413_ _0467_ _0589_ _0475_ _0592_ _1888_ vssd1 vssd1 vccd1 vccd1 _1889_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_2_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6393_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2736_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5344_ _3330_ _3353_ vssd1 vssd1 vccd1 vccd1 _1820_ sky130_fd_sc_hd__nand2_1
X_5275_ _1619_ _0506_ _1749_ _1750_ _1751_ vssd1 vssd1 vccd1 vccd1 _1752_ sky130_fd_sc_hd__o2111a_1
X_4226_ _0421_ vssd1 vssd1 vccd1 vccd1 _0711_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ egd_top.BitStream_buffer.BS_buffer\[90\] vssd1 vssd1 vccd1 vccd1 _0642_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4088_ _0573_ vssd1 vssd1 vccd1 vccd1 _0574_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0__2926_ _2926_ vssd1 vssd1 vccd1 vccd1 clknet_0__2926_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 la_data_in_58_43[7] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_8
X_3390_ _2941_ vssd1 vssd1 vccd1 vccd1 _2945_ sky130_fd_sc_hd__inv_2
X_5060_ _3128_ _3161_ vssd1 vssd1 vccd1 vccd1 _1538_ sky130_fd_sc_hd__nand2_1
X_4011_ _3103_ _0470_ vssd1 vssd1 vccd1 vccd1 _0497_ sky130_fd_sc_hd__and2_1
X_5962_ egd_top.BitStream_buffer.buffer_index\[6\] egd_top.BitStream_buffer.buffer_index\[5\]
+ _2972_ _3002_ vssd1 vssd1 vccd1 vccd1 _2414_ sky130_fd_sc_hd__or4b_4
XFILLER_0_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4913_ _0559_ _0545_ _1390_ _1391_ _1392_ vssd1 vssd1 vccd1 vccd1 _1393_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5893_ _0535_ _0588_ _0531_ _0591_ _2364_ vssd1 vssd1 vccd1 vccd1 _2365_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4844_ _3309_ _0675_ vssd1 vssd1 vccd1 vccd1 _1324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4775_ _0515_ _0488_ _0509_ _0492_ _1255_ vssd1 vssd1 vccd1 vccd1 _1256_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6514_ _2848_ _2849_ _2714_ vssd1 vssd1 vccd1 vccd1 _2850_ sky130_fd_sc_hd__o21ai_1
X_3726_ _3258_ _3259_ vssd1 vssd1 vccd1 vccd1 _3260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6445_ _2758_ _2786_ vssd1 vssd1 vccd1 vccd1 _2787_ sky130_fd_sc_hd__or2_1
X_3657_ _3061_ _3167_ vssd1 vssd1 vccd1 vccd1 _3191_ sky130_fd_sc_hd__and2_1
X_6376_ net18 _2956_ vssd1 vssd1 vccd1 vccd1 _2719_ sky130_fd_sc_hd__nor2_1
X_3588_ _3121_ vssd1 vssd1 vccd1 vccd1 _3122_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5327_ _3341_ _3231_ _3347_ _3235_ _1802_ vssd1 vssd1 vccd1 vccd1 _1803_ sky130_fd_sc_hd__a221oi_1
X_5258_ _0411_ _0432_ _0447_ _0436_ _1734_ vssd1 vssd1 vccd1 vccd1 _1735_ sky130_fd_sc_hd__a221oi_1
X_4209_ _0363_ _0362_ _0689_ _0366_ _0693_ vssd1 vssd1 vccd1 vccd1 _0694_ sky130_fd_sc_hd__a221oi_1
X_5189_ _1664_ _1665_ vssd1 vssd1 vccd1 vccd1 _1666_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ _3155_ _3247_ vssd1 vssd1 vccd1 vccd1 _1042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4491_ _0853_ _0386_ _0973_ vssd1 vssd1 vccd1 vccd1 _0974_ sky130_fd_sc_hd__o21ai_1
X_3511_ net9 _3047_ _3006_ vssd1 vssd1 vccd1 vccd1 _3048_ sky130_fd_sc_hd__mux2_1
X_3442_ _2985_ _2993_ _2988_ vssd1 vssd1 vccd1 vccd1 _2994_ sky130_fd_sc_hd__o21bai_1
X_6230_ egd_top.BitStream_buffer.pc_previous\[6\] _2601_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[6\]
+ sky130_fd_sc_hd__xor2_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _2928_ _2929_ _2930_ vssd1 vssd1 vccd1 vccd1 _2931_ sky130_fd_sc_hd__o21ai_1
X_6161_ net8 _3144_ _2520_ vssd1 vssd1 vccd1 vccd1 _2551_ sky130_fd_sc_hd__mux2_1
X_5112_ _1588_ _1589_ vssd1 vssd1 vccd1 vccd1 _1590_ sky130_fd_sc_hd__nand2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ net14 _0417_ _2486_ vssd1 vssd1 vccd1 vccd1 _2504_ sky130_fd_sc_hd__mux2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _0750_ _0584_ vssd1 vssd1 vccd1 vccd1 _1522_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5945_ _2402_ _2396_ vssd1 vssd1 vccd1 vccd1 _2403_ sky130_fd_sc_hd__and2_1
X_5876_ _0347_ _0505_ _2345_ _2346_ _2347_ vssd1 vssd1 vccd1 vccd1 _2348_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _0574_ _3218_ _0582_ _3221_ vssd1 vssd1 vccd1 vccd1 _1307_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ _0981_ _0426_ vssd1 vssd1 vccd1 vccd1 _1239_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3709_ _3225_ _3231_ _3232_ _3235_ _3242_ vssd1 vssd1 vccd1 vccd1 _3243_ sky130_fd_sc_hd__a221oi_1
X_4689_ _3160_ _3247_ vssd1 vssd1 vccd1 vccd1 _1170_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6428_ _2765_ _2769_ _2710_ vssd1 vssd1 vccd1 vccd1 _2770_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6359_ _2701_ _1406_ _2666_ vssd1 vssd1 vccd1 vccd1 _2702_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 egd_top.BitStream_buffer.buffer_index\[5\] vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3991_ _3061_ _0469_ vssd1 vssd1 vccd1 vccd1 _0477_ sky130_fd_sc_hd__and2_2
XFILLER_0_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5730_ _0398_ _3102_ vssd1 vssd1 vccd1 vccd1 _2203_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5661_ _3266_ _3083_ _0651_ _3091_ vssd1 vssd1 vccd1 vccd1 _2134_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4612_ _0389_ _0328_ _0695_ _0332_ _1093_ vssd1 vssd1 vccd1 vccd1 _1094_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5592_ _3188_ _3362_ _2065_ vssd1 vssd1 vccd1 vccd1 _2066_ sky130_fd_sc_hd__o21ai_1
X_4543_ _0994_ _1011_ _1025_ vssd1 vssd1 vccd1 vccd1 _1026_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4474_ _3365_ _3010_ vssd1 vssd1 vccd1 vccd1 _0957_ sky130_fd_sc_hd__nand2_1
X_6213_ net8 _0674_ net197 vssd1 vssd1 vccd1 vccd1 _2587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3425_ _2978_ _2971_ _2972_ vssd1 vssd1 vccd1 vccd1 _2979_ sky130_fd_sc_hd__and3_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _2539_ _2529_ vssd1 vssd1 vccd1 vccd1 _2540_ sky130_fd_sc_hd__and2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _2492_ vssd1 vssd1 vccd1 vccd1 _0229_ sky130_fd_sc_hd__clkbuf_1
X_6681__11 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__inv_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _0508_ _0531_ vssd1 vssd1 vccd1 vccd1 _1505_ sky130_fd_sc_hd__nand2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5928_ net2 _0540_ _2380_ vssd1 vssd1 vccd1 vccd1 _2391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5859_ _0981_ _0439_ _2330_ vssd1 vssd1 vccd1 vccd1 _2331_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _0675_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6900_ net98 _0303_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[122\]
+ sky130_fd_sc_hd__dfxtp_1
X_6831_ net185 _0234_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[45\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6762_ net116 _0165_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[91\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _0459_ vssd1 vssd1 vccd1 vccd1 _0460_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6718__45 clknet_1_0__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__inv_2
X_5713_ _3034_ _3355_ _3037_ _3359_ _2185_ vssd1 vssd1 vccd1 vccd1 _2186_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5644_ _0728_ _0555_ vssd1 vssd1 vccd1 vccd1 _2118_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6733__59 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__inv_2
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5575_ _2047_ _2048_ vssd1 vssd1 vccd1 vccd1 _2049_ sky130_fd_sc_hd__nor2_1
X_4526_ _1007_ _1008_ vssd1 vssd1 vccd1 vccd1 _1009_ sky130_fd_sc_hd__nand2_1
X_4457_ _3318_ vssd1 vssd1 vccd1 vccd1 _0940_ sky130_fd_sc_hd__inv_2
X_3408_ _2961_ vssd1 vssd1 vccd1 vccd1 _2962_ sky130_fd_sc_hd__inv_2
X_4388_ _0512_ _0509_ vssd1 vssd1 vccd1 vccd1 _0872_ sky130_fd_sc_hd__nand2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ net4 _3102_ _2521_ vssd1 vssd1 vccd1 vccd1 _2528_ sky130_fd_sc_hd__mux2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _2480_ vssd1 vssd1 vccd1 vccd1 _0234_ sky130_fd_sc_hd__clkbuf_1
X_5009_ _0767_ _0414_ _1485_ _1486_ _1487_ vssd1 vssd1 vccd1 vccd1 _1488_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2923_ clknet_0__2923_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2923_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3690_ _3181_ _3195_ _3209_ _3223_ vssd1 vssd1 vccd1 vccd1 _3224_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5360_ _1714_ _0345_ _0384_ _0349_ vssd1 vssd1 vccd1 vccd1 _1836_ sky130_fd_sc_hd__o22ai_1
X_5291_ _0516_ _0595_ _0734_ _0598_ vssd1 vssd1 vccd1 vccd1 _1768_ sky130_fd_sc_hd__o22ai_1
X_4311_ _0642_ _3238_ _0794_ _3241_ vssd1 vssd1 vccd1 vccd1 _0795_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4242_ _0723_ _0472_ _0724_ _0726_ vssd1 vssd1 vccd1 vccd1 _0727_ sky130_fd_sc_hd__o211a_1
X_4173_ _3282_ _3281_ _3318_ _3285_ _0657_ vssd1 vssd1 vccd1 vccd1 _0658_ sky130_fd_sc_hd__a221oi_1
X_6645__134 clknet_1_1__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__inv_2
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6814_ net168 _0217_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[62\]
+ sky130_fd_sc_hd__dfxtp_1
X_3957_ egd_top.BitStream_buffer.BS_buffer\[49\] vssd1 vssd1 vccd1 vccd1 _0443_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3888_ _0367_ _0369_ _0373_ vssd1 vssd1 vccd1 vccd1 _0374_ sky130_fd_sc_hd__o21ai_1
X_5627_ _0477_ _0353_ _0480_ _0356_ vssd1 vssd1 vccd1 vccd1 _2101_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5558_ _0554_ _3189_ _2031_ vssd1 vssd1 vccd1 vccd1 _2032_ sky130_fd_sc_hd__o21ai_1
X_4509_ _0455_ _0450_ _3107_ _0454_ _0991_ vssd1 vssd1 vccd1 vccd1 _0992_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5489_ _1954_ _1957_ _1960_ _1963_ vssd1 vssd1 vccd1 vccd1 _1964_ sky130_fd_sc_hd__and4_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _1327_ _1331_ _1336_ _1339_ vssd1 vssd1 vccd1 vccd1 _1340_ sky130_fd_sc_hd__and4_1
X_3811_ egd_top.BitStream_buffer.BS_buffer\[102\] vssd1 vssd1 vccd1 vccd1 _3345_ sky130_fd_sc_hd__clkbuf_4
X_6530_ _1282_ _2806_ _2864_ _2689_ vssd1 vssd1 vccd1 vccd1 _2865_ sky130_fd_sc_hd__a211o_1
X_4791_ _0756_ _0570_ vssd1 vssd1 vccd1 vccd1 _1272_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3742_ _3271_ _3272_ _3274_ _3275_ vssd1 vssd1 vccd1 vccd1 _3276_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3673_ _3206_ _3010_ vssd1 vssd1 vccd1 vccd1 _3207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6461_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] _2771_ vssd1 vssd1
+ vccd1 vccd1 _2802_ sky130_fd_sc_hd__or2_1
X_5412_ _0734_ _0595_ _0504_ _0598_ vssd1 vssd1 vccd1 vccd1 _1888_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6392_ _2734_ vssd1 vssd1 vccd1 vccd1 _2735_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5343_ _3326_ _3357_ vssd1 vssd1 vccd1 vccd1 _1819_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5274_ _1373_ _0518_ vssd1 vssd1 vccd1 vccd1 _1751_ sky130_fd_sc_hd__or2_1
X_4225_ _0420_ _0411_ vssd1 vssd1 vccd1 vccd1 _0710_ sky130_fd_sc_hd__nand2_1
X_4156_ _0630_ _0633_ _0637_ _0640_ vssd1 vssd1 vccd1 vccd1 _0641_ sky130_fd_sc_hd__and4_1
X_4087_ egd_top.BitStream_buffer.BS_buffer\[2\] vssd1 vssd1 vccd1 vccd1 _0573_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_0__2925_ _2925_ vssd1 vssd1 vccd1 vccd1 clknet_0__2925_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4989_ _1466_ _1467_ vssd1 vssd1 vccd1 vccd1 _1468_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 la_data_in_58_43[8] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4010_ _0495_ vssd1 vssd1 vccd1 vccd1 _0496_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5961_ _2413_ vssd1 vssd1 vccd1 vccd1 _0264_ sky130_fd_sc_hd__clkbuf_1
X_4912_ _0596_ _0556_ vssd1 vssd1 vccd1 vccd1 _1392_ sky130_fd_sc_hd__or2_1
X_5892_ _0862_ _0594_ _0995_ _0597_ vssd1 vssd1 vccd1 vccd1 _2364_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4843_ _1311_ _1316_ _1319_ _1322_ vssd1 vssd1 vccd1 vccd1 _1323_ sky130_fd_sc_hd__and4_1
XFILLER_0_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4774_ _0504_ _0496_ _1254_ vssd1 vssd1 vccd1 vccd1 _1255_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6513_ _2847_ _2840_ vssd1 vssd1 vccd1 vccd1 _2849_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3725_ egd_top.BitStream_buffer.BS_buffer\[82\] vssd1 vssd1 vccd1 vccd1 _3259_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6444_ _2785_ _2959_ vssd1 vssd1 vccd1 vccd1 _2786_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3656_ _3189_ vssd1 vssd1 vccd1 vccd1 _3190_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6375_ _2717_ _2650_ vssd1 vssd1 vccd1 vccd1 _2718_ sky130_fd_sc_hd__nand2_1
X_3587_ _3070_ egd_top.BitStream_buffer.pc\[2\] _3096_ vssd1 vssd1 vccd1 vccd1 _3121_
+ sky130_fd_sc_hd__and3_1
X_5326_ _1196_ _3238_ _1320_ _3241_ vssd1 vssd1 vccd1 vccd1 _1802_ sky130_fd_sc_hd__o22ai_1
X_5257_ _0424_ _0440_ _1733_ vssd1 vssd1 vccd1 vccd1 _1734_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4208_ _0690_ _0369_ _0692_ vssd1 vssd1 vccd1 vccd1 _0693_ sky130_fd_sc_hd__o21ai_1
X_5188_ _3160_ _3265_ vssd1 vssd1 vccd1 vccd1 _1665_ sky130_fd_sc_hd__nand2_1
X_4139_ _3160_ _3156_ vssd1 vssd1 vccd1 vccd1 _0624_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ egd_top.BitStream_buffer.BS_buffer\[125\] vssd1 vssd1 vccd1 vccd1 _3047_ sky130_fd_sc_hd__clkbuf_4
X_4490_ _0388_ _0443_ vssd1 vssd1 vccd1 vccd1 _0973_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3441_ net28 _2976_ _2974_ vssd1 vssd1 vccd1 vccd1 _2993_ sky130_fd_sc_hd__o21ai_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ net34 vssd1 vssd1 vccd1 vccd1 _2930_ sky130_fd_sc_hd__inv_2
X_6160_ _2550_ vssd1 vssd1 vccd1 vccd1 _0202_ sky130_fd_sc_hd__clkbuf_1
X_5111_ _0338_ _0437_ vssd1 vssd1 vccd1 vccd1 _1589_ sky130_fd_sc_hd__nand2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _2503_ vssd1 vssd1 vccd1 vccd1 _0224_ sky130_fd_sc_hd__clkbuf_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _0494_ _0561_ _1518_ _1519_ _1520_ vssd1 vssd1 vccd1 vccd1 _1521_ sky130_fd_sc_hd__o2111a_1
X_5944_ net12 egd_top.BitStream_buffer.BS_buffer\[10\] _2380_ vssd1 vssd1 vccd1 vccd1
+ _2402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5875_ _0690_ _0517_ vssd1 vssd1 vccd1 vccd1 _2347_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _3031_ _3198_ _3034_ _3201_ _1305_ vssd1 vssd1 vccd1 vccd1 _1306_ sky130_fd_sc_hd__a221oi_1
X_6602__94 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__inv_2
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4757_ _0420_ _0455_ vssd1 vssd1 vccd1 vccd1 _1238_ sky130_fd_sc_hd__nand2_1
X_3708_ _3236_ _3238_ _3239_ _3241_ vssd1 vssd1 vccd1 vccd1 _3242_ sky130_fd_sc_hd__o22ai_1
X_4688_ _3155_ _3259_ vssd1 vssd1 vccd1 vccd1 _1169_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6427_ _2709_ _2768_ _2726_ vssd1 vssd1 vccd1 vccd1 _2769_ sky130_fd_sc_hd__nand3_1
X_3639_ _3172_ vssd1 vssd1 vccd1 vccd1 _3173_ sky130_fd_sc_hd__buf_6
X_6358_ _2700_ vssd1 vssd1 vccd1 vccd1 _2701_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5309_ _1532_ _3124_ _1782_ _1783_ _1784_ vssd1 vssd1 vccd1 vccd1 _1785_ sky130_fd_sc_hd__o2111a_1
X_6289_ _2636_ _2372_ vssd1 vssd1 vccd1 vccd1 _2637_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6739__65 clknet_1_0__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__inv_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 _2612_ vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3990_ _0474_ _0475_ vssd1 vssd1 vccd1 vccd1 _0476_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5660_ _0898_ _2131_ _2133_ vssd1 vssd1 vccd1 vccd1 _0285_ sky130_fd_sc_hd__o21a_1
X_4611_ _1091_ _1092_ vssd1 vssd1 vccd1 vccd1 _1093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5591_ _3364_ _3037_ vssd1 vssd1 vccd1 vccd1 _2065_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4542_ _1015_ _1019_ _1021_ _1024_ vssd1 vssd1 vccd1 vccd1 _1025_ sky130_fd_sc_hd__and4_1
X_4473_ _0952_ _3338_ _0953_ _0954_ _0955_ vssd1 vssd1 vccd1 vccd1 _0956_ sky130_fd_sc_hd__o2111a_1
X_6212_ _2586_ vssd1 vssd1 vccd1 vccd1 _0186_ sky130_fd_sc_hd__clkbuf_1
X_3424_ net200 vssd1 vssd1 vccd1 vccd1 _2978_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ net14 _3076_ _2521_ vssd1 vssd1 vccd1 vccd1 _2539_ sky130_fd_sc_hd__mux2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _2491_ _2475_ vssd1 vssd1 vccd1 vccd1 _2492_ sky130_fd_sc_hd__and2_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _0503_ _0488_ _0467_ _0492_ _1503_ vssd1 vssd1 vccd1 vccd1 _1504_ sky130_fd_sc_hd__a221oi_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5927_ _2390_ vssd1 vssd1 vccd1 vccd1 _0275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5858_ _0441_ _0455_ vssd1 vssd1 vccd1 vccd1 _2330_ sky130_fd_sc_hd__nand2_1
X_5789_ _3266_ _3123_ _2258_ _2259_ _2260_ vssd1 vssd1 vccd1 vccd1 _2261_ sky130_fd_sc_hd__o2111a_1
X_4809_ _3076_ _3101_ _3085_ _3106_ _1288_ vssd1 vssd1 vccd1 vccd1 _1289_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6830_ net184 _0233_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[46\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6761_ net115 _0164_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[92\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5712_ _3216_ _3362_ _2184_ vssd1 vssd1 vccd1 vccd1 _2185_ sky130_fd_sc_hd__o21ai_1
X_3973_ _3145_ _0395_ vssd1 vssd1 vccd1 vccd1 _0459_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5643_ _0550_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _2117_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5574_ _3270_ _3331_ _3273_ _3327_ vssd1 vssd1 vccd1 vccd1 _2048_ sky130_fd_sc_hd__a22o_1
X_4525_ _0534_ _0525_ vssd1 vssd1 vccd1 vccd1 _1008_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4456_ _0937_ _0938_ vssd1 vssd1 vccd1 vccd1 _0939_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4387_ _0508_ _0467_ vssd1 vssd1 vccd1 vccd1 _0871_ sky130_fd_sc_hd__nand2_1
X_3407_ _2958_ _2960_ vssd1 vssd1 vccd1 vccd1 _2961_ sky130_fd_sc_hd__nand2_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6126_ _2527_ vssd1 vssd1 vccd1 vccd1 _0213_ sky130_fd_sc_hd__clkbuf_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _2479_ _2475_ vssd1 vssd1 vccd1 vccd1 _2480_ sky130_fd_sc_hd__and2_1
X_6622__113 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__inv_2
X_5008_ _3108_ _0426_ vssd1 vssd1 vccd1 vccd1 _1487_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__2922_ clknet_0__2922_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2922_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4310_ egd_top.BitStream_buffer.BS_buffer\[91\] vssd1 vssd1 vccd1 vccd1 _0794_ sky130_fd_sc_hd__inv_2
X_5290_ _0559_ _0576_ _0750_ _0580_ _1766_ vssd1 vssd1 vccd1 vccd1 _1767_ sky130_fd_sc_hd__o221a_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4241_ _0725_ vssd1 vssd1 vccd1 vccd1 _0726_ sky130_fd_sc_hd__inv_2
X_4172_ _3291_ _3289_ _0656_ _3293_ vssd1 vssd1 vccd1 vccd1 _0657_ sky130_fd_sc_hd__o22ai_1
X_6813_ net167 _0216_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[63\]
+ sky130_fd_sc_hd__dfxtp_1
X_3956_ _0441_ vssd1 vssd1 vccd1 vccd1 _0442_ sky130_fd_sc_hd__clkbuf_4
X_6675_ clknet_1_1__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2922_ sky130_fd_sc_hd__buf_1
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5626_ _0473_ _0346_ vssd1 vssd1 vccd1 vccd1 _2100_ sky130_fd_sc_hd__nand2_1
X_3887_ _0371_ _0372_ vssd1 vssd1 vccd1 vccd1 _0373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5557_ _3191_ _0548_ vssd1 vssd1 vccd1 vccd1 _2031_ sky130_fd_sc_hd__nand2_1
X_5488_ _0701_ _0379_ _0417_ _0383_ _1962_ vssd1 vssd1 vccd1 vccd1 _1963_ sky130_fd_sc_hd__a221oi_1
X_4508_ _0767_ _0458_ _0990_ vssd1 vssd1 vccd1 vccd1 _0991_ sky130_fd_sc_hd__o21ai_1
X_4439_ egd_top.BitStream_buffer.BS_buffer\[115\] vssd1 vssd1 vccd1 vccd1 _0922_ sky130_fd_sc_hd__inv_2
X_6109_ _2515_ vssd1 vssd1 vccd1 vccd1 _0218_ sky130_fd_sc_hd__clkbuf_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6629__119 clknet_1_0__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__inv_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3810_ _3343_ vssd1 vssd1 vccd1 vccd1 _3344_ sky130_fd_sc_hd__clkbuf_4
X_4790_ _0566_ egd_top.BitStream_buffer.BS_buffer\[13\] vssd1 vssd1 vccd1 vccd1 _1271_
+ sky130_fd_sc_hd__nand2_1
X_3741_ egd_top.BitStream_buffer.BS_buffer\[87\] vssd1 vssd1 vccd1 vccd1 _3275_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3672_ _3205_ vssd1 vssd1 vccd1 vccd1 _3206_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6460_ _2771_ egd_top.BitStream_buffer.BitStream_buffer_output\[12\] vssd1 vssd1
+ vccd1 vccd1 _2801_ sky130_fd_sc_hd__nand2_1
X_6391_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ vssd1 vssd1 vccd1 vccd1 _2734_ sky130_fd_sc_hd__nor2_1
X_5411_ _0593_ _0576_ _0559_ _0580_ _1886_ vssd1 vssd1 vccd1 vccd1 _1887_ sky130_fd_sc_hd__o221a_1
X_5342_ _3019_ _3303_ _3022_ _3307_ _1817_ vssd1 vssd1 vccd1 vccd1 _1818_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5273_ _0512_ _0531_ vssd1 vssd1 vccd1 vccd1 _1750_ sky130_fd_sc_hd__nand2_1
X_4224_ _0416_ _0423_ vssd1 vssd1 vccd1 vccd1 _0709_ sky130_fd_sc_hd__nand2_1
X_4155_ _3053_ _3212_ _0607_ _3215_ _0639_ vssd1 vssd1 vccd1 vccd1 _0640_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_37_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4086_ _0559_ _0561_ _0564_ _0567_ _0571_ vssd1 vssd1 vccd1 vccd1 _0572_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2924_ _2924_ vssd1 vssd1 vccd1 vccd1 clknet_0__2924_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4988_ _0338_ _0695_ vssd1 vssd1 vccd1 vccd1 _1467_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6727_ clknet_1_0__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2926_ sky130_fd_sc_hd__buf_1
X_3939_ _3090_ _0395_ vssd1 vssd1 vccd1 vccd1 _0425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5609_ _2073_ _2076_ _2079_ _2082_ vssd1 vssd1 vccd1 vccd1 _2083_ sky130_fd_sc_hd__and4_1
X_6702__30 clknet_1_1__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__inv_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6674__161 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__inv_2
XFILLER_0_64_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 la_data_in_58_43[9] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5960_ _2412_ _2396_ vssd1 vssd1 vccd1 vccd1 _2413_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _0551_ egd_top.BitStream_buffer.BS_buffer\[10\] vssd1 vssd1 vccd1 vccd1 _1391_
+ sky130_fd_sc_hd__nand2_1
X_5891_ _1022_ _0575_ _0890_ _0579_ _2362_ vssd1 vssd1 vccd1 vccd1 _2363_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4842_ _3341_ _3281_ _3347_ _3285_ _1321_ vssd1 vssd1 vccd1 vccd1 _1322_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4773_ _0498_ _0467_ vssd1 vssd1 vccd1 vccd1 _1254_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6512_ _2840_ _2847_ vssd1 vssd1 vccd1 vccd1 _2848_ sky130_fd_sc_hd__nor2_1
X_3724_ _3257_ vssd1 vssd1 vccd1 vccd1 _3258_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6443_ _2770_ _2784_ vssd1 vssd1 vccd1 vccd1 _2785_ sky130_fd_sc_hd__nand2_1
X_3655_ _3072_ _3167_ vssd1 vssd1 vccd1 vccd1 _3189_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6374_ _2693_ _2667_ _2685_ _2716_ _2659_ vssd1 vssd1 vccd1 vccd1 _2717_ sky130_fd_sc_hd__a311o_1
X_3586_ _3119_ vssd1 vssd1 vccd1 vccd1 _3120_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5325_ _1792_ _1795_ _1798_ _1800_ vssd1 vssd1 vccd1 vccd1 _1801_ sky130_fd_sc_hd__and4_1
X_5256_ _0442_ _0421_ vssd1 vssd1 vccd1 vccd1 _1733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4207_ _0371_ _0691_ vssd1 vssd1 vccd1 vccd1 _0692_ sky130_fd_sc_hd__nand2_1
X_5187_ _3155_ _3272_ vssd1 vssd1 vccd1 vccd1 _1664_ sky130_fd_sc_hd__nand2_1
X_4138_ _3155_ _3144_ vssd1 vssd1 vccd1 vccd1 _0623_ sky130_fd_sc_hd__nand2_1
X_4069_ _3122_ _0543_ vssd1 vssd1 vccd1 vccd1 _0555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3440_ _2991_ _2988_ _2989_ _2992_ vssd1 vssd1 vccd1 vccd1 _0316_ sky130_fd_sc_hd__o211a_1
X_3371_ net32 net31 vssd1 vssd1 vccd1 vccd1 _2929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5110_ _0334_ _0443_ vssd1 vssd1 vccd1 vccd1 _1588_ sky130_fd_sc_hd__nand2_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ _2501_ _2502_ vssd1 vssd1 vccd1 vccd1 _2503_ sky130_fd_sc_hd__and2_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _1022_ _0570_ vssd1 vssd1 vccd1 vccd1 _1520_ sky130_fd_sc_hd__or2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6599__91 clknet_1_1__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__inv_2
X_5943_ _2401_ vssd1 vssd1 vccd1 vccd1 _0270_ sky130_fd_sc_hd__clkbuf_1
X_5874_ _0511_ _0689_ vssd1 vssd1 vccd1 vccd1 _2346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4825_ _0628_ _3204_ _1304_ vssd1 vssd1 vccd1 vccd1 _1305_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4756_ _0416_ _0451_ vssd1 vssd1 vccd1 vccd1 _1237_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3707_ _3240_ vssd1 vssd1 vccd1 vccd1 _3241_ sky130_fd_sc_hd__clkbuf_4
X_4687_ _0900_ _3124_ _1165_ _1166_ _1167_ vssd1 vssd1 vccd1 vccd1 _1168_ sky130_fd_sc_hd__o2111a_1
X_6426_ _2766_ _2767_ vssd1 vssd1 vccd1 vccd1 _2768_ sky130_fd_sc_hd__nand2_1
X_3638_ _3171_ vssd1 vssd1 vccd1 vccd1 _3172_ sky130_fd_sc_hd__clkbuf_2
X_6357_ _2681_ _2691_ _2686_ vssd1 vssd1 vccd1 vccd1 _2700_ sky130_fd_sc_hd__nand3_4
X_3569_ _3097_ _2963_ vssd1 vssd1 vccd1 vccd1 _3103_ sky130_fd_sc_hd__nor2_4
XFILLER_0_11_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5308_ _1284_ _3141_ vssd1 vssd1 vccd1 vccd1 _1784_ sky130_fd_sc_hd__or2_1
X_6288_ net11 _3232_ _2613_ vssd1 vssd1 vccd1 vccd1 _2636_ sky130_fd_sc_hd__mux2_1
X_5239_ _0352_ _0695_ _0355_ _0437_ vssd1 vssd1 vccd1 vccd1 _1716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 egd_top.BitStream_buffer.buffer_index\[6\] vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4610_ _0338_ _0376_ vssd1 vssd1 vccd1 vccd1 _1092_ sky130_fd_sc_hd__nand2_1
X_5590_ _0922_ _3337_ _2061_ _2062_ _2063_ vssd1 vssd1 vccd1 vccd1 _2064_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4541_ _0489_ _0589_ _0493_ _0592_ _1023_ vssd1 vssd1 vccd1 vccd1 _1024_ sky130_fd_sc_hd__a221oi_1
X_4472_ _0668_ _3350_ vssd1 vssd1 vccd1 vccd1 _0955_ sky130_fd_sc_hd__or2_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3423_ _2974_ _2976_ vssd1 vssd1 vccd1 vccd1 _2977_ sky130_fd_sc_hd__nand2_1
X_6211_ _2585_ _2581_ vssd1 vssd1 vccd1 vccd1 _2586_ sky130_fd_sc_hd__and2_1
X_6142_ _2538_ vssd1 vssd1 vccd1 vccd1 _0208_ sky130_fd_sc_hd__clkbuf_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ net5 _0429_ _2486_ vssd1 vssd1 vccd1 vccd1 _2491_ sky130_fd_sc_hd__mux2_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _0723_ _0496_ _1502_ vssd1 vssd1 vccd1 vccd1 _1503_ sky130_fd_sc_hd__o21ai_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5926_ _2389_ _3042_ vssd1 vssd1 vccd1 vccd1 _2390_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5857_ _3086_ _0413_ _2326_ _2327_ _2328_ vssd1 vssd1 vccd1 vccd1 _2329_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5788_ _1776_ _3140_ vssd1 vssd1 vccd1 vccd1 _2260_ sky130_fd_sc_hd__or2_1
X_4808_ _0620_ _3111_ _1287_ vssd1 vssd1 vccd1 vccd1 _1288_ sky130_fd_sc_hd__o21ai_1
X_4739_ _1218_ _1219_ vssd1 vssd1 vccd1 vccd1 _1220_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6409_ _2742_ _2743_ _2748_ _2751_ vssd1 vssd1 vccd1 vccd1 _2752_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6593__86 clknet_1_1__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__inv_2
XFILLER_0_34_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6760_ net114 _0163_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[93\]
+ sky130_fd_sc_hd__dfxtp_1
X_5711_ _3364_ _3040_ vssd1 vssd1 vccd1 vccd1 _2184_ sky130_fd_sc_hd__nand2_1
X_3972_ _0457_ vssd1 vssd1 vccd1 vccd1 _0458_ sky130_fd_sc_hd__clkbuf_4
X_5642_ _0546_ _0493_ vssd1 vssd1 vccd1 vccd1 _2116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5573_ _0940_ _3263_ _1069_ _3267_ vssd1 vssd1 vccd1 vccd1 _2047_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_53_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4524_ _0530_ _0359_ vssd1 vssd1 vccd1 vccd1 _1007_ sky130_fd_sc_hd__nand2_1
X_4455_ _3271_ _0804_ _3274_ _3225_ vssd1 vssd1 vccd1 vccd1 _0938_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4386_ _0493_ _0488_ _0499_ _0492_ _0869_ vssd1 vssd1 vccd1 vccd1 _0870_ sky130_fd_sc_hd__a221oi_1
X_3406_ _2959_ egd_top.BitStream_buffer.pc_previous\[0\] vssd1 vssd1 vccd1 vccd1 _2960_
+ sky130_fd_sc_hd__nand2_4
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _2526_ _2502_ vssd1 vssd1 vccd1 vccd1 _2527_ sky130_fd_sc_hd__and2_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ net9 _0380_ _2450_ vssd1 vssd1 vccd1 vccd1 _2479_ sky130_fd_sc_hd__mux2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _0420_ _3115_ vssd1 vssd1 vccd1 vccd1 _1486_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6889_ net87 _0292_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_5909_ _2377_ _2372_ _3003_ vssd1 vssd1 vccd1 vccd1 _2378_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_1__f__2921_ clknet_0__2921_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2921_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6723__50 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__inv_2
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4240_ _0478_ _0482_ _0481_ _0535_ vssd1 vssd1 vccd1 vccd1 _0725_ sky130_fd_sc_hd__a22o_1
X_4171_ _3278_ vssd1 vssd1 vccd1 vccd1 _0656_ sky130_fd_sc_hd__inv_2
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6812_ net166 _0215_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[64\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3955_ _3112_ _0395_ vssd1 vssd1 vccd1 vccd1 _0441_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3886_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _0372_ sky130_fd_sc_hd__clkbuf_4
X_5625_ _2083_ _2098_ vssd1 vssd1 vccd1 vccd1 _2099_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5556_ _0573_ _3169_ _0581_ _3172_ _2029_ vssd1 vssd1 vccd1 vccd1 _2030_ sky130_fd_sc_hd__a221oi_1
X_5487_ _0711_ _0386_ _1961_ vssd1 vssd1 vccd1 vccd1 _1962_ sky130_fd_sc_hd__o21ai_1
X_4507_ _0460_ _3115_ vssd1 vssd1 vccd1 vccd1 _0990_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4438_ _3040_ _3184_ _3044_ _3187_ _0920_ vssd1 vssd1 vccd1 vccd1 _0921_ sky130_fd_sc_hd__a221oi_1
X_4369_ egd_top.BitStream_buffer.BS_buffer\[50\] vssd1 vssd1 vccd1 vccd1 _0853_ sky130_fd_sc_hd__inv_2
X_6108_ _2514_ _2502_ vssd1 vssd1 vccd1 vccd1 _2515_ sky130_fd_sc_hd__and2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _2467_ vssd1 vssd1 vccd1 vccd1 _0240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _3273_ vssd1 vssd1 vccd1 vccd1 _3274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3671_ _3112_ _3167_ vssd1 vssd1 vccd1 vccd1 _3205_ sky130_fd_sc_hd__and2_1
X_6390_ _2701_ _2666_ vssd1 vssd1 vccd1 vccd1 _2733_ sky130_fd_sc_hd__and2_1
X_5410_ _0596_ _0584_ vssd1 vssd1 vccd1 vccd1 _1886_ sky130_fd_sc_hd__or2_1
X_5341_ _1815_ _1816_ vssd1 vssd1 vccd1 vccd1 _1817_ sky130_fd_sc_hd__nand2_1
X_5272_ _0508_ _0525_ vssd1 vssd1 vccd1 vccd1 _1749_ sky130_fd_sc_hd__nand2_1
X_4223_ _0447_ vssd1 vssd1 vccd1 vccd1 _0708_ sky130_fd_sc_hd__inv_2
X_4154_ _3219_ _3218_ _0638_ _3221_ vssd1 vssd1 vccd1 vccd1 _0639_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4085_ _0568_ _0570_ vssd1 vssd1 vccd1 vccd1 _0571_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__2923_ _2923_ vssd1 vssd1 vccd1 vccd1 clknet_0__2923_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4987_ _0334_ _0437_ vssd1 vssd1 vccd1 vccd1 _1466_ sky130_fd_sc_hd__nand2_1
X_3938_ _0423_ vssd1 vssd1 vccd1 vccd1 _0424_ sky130_fd_sc_hd__inv_2
X_3869_ _0354_ vssd1 vssd1 vccd1 vccd1 _0355_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5608_ _0417_ _0378_ _0423_ _0382_ _2081_ vssd1 vssd1 vccd1 vccd1 _2082_ sky130_fd_sc_hd__a221oi_1
X_5539_ _2013_ _2996_ _2938_ vssd1 vssd1 vccd1 vccd1 _2014_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput17 la_data_in_60_59[0] vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__buf_2
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4910_ _0547_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1390_
+ sky130_fd_sc_hd__nand2_1
X_5890_ _1150_ _0583_ vssd1 vssd1 vccd1 vccd1 _2362_ sky130_fd_sc_hd__or2_1
X_4841_ _1196_ _3289_ _1320_ _3293_ vssd1 vssd1 vccd1 vccd1 _1321_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4772_ _1249_ _0472_ _1250_ _1252_ vssd1 vssd1 vccd1 vccd1 _1253_ sky130_fd_sc_hd__o211a_1
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6511_ _2811_ _2846_ vssd1 vssd1 vccd1 vccd1 _2847_ sky130_fd_sc_hd__nand2_1
X_3723_ _3098_ _3227_ vssd1 vssd1 vccd1 vccd1 _3257_ sky130_fd_sc_hd__and2_1
X_3654_ _3040_ vssd1 vssd1 vccd1 vccd1 _3188_ sky130_fd_sc_hd__inv_2
X_6442_ _2776_ _2783_ vssd1 vssd1 vccd1 vccd1 _2784_ sky130_fd_sc_hd__nor2_1
X_6678__8 clknet_1_1__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__inv_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6373_ _2959_ vssd1 vssd1 vccd1 vccd1 _2716_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3585_ egd_top.BitStream_buffer.BS_buffer\[71\] vssd1 vssd1 vccd1 vccd1 _3119_ sky130_fd_sc_hd__clkbuf_4
X_5324_ egd_top.BitStream_buffer.BS_buffer\[8\] _3212_ egd_top.BitStream_buffer.BS_buffer\[9\]
+ _3215_ _1799_ vssd1 vssd1 vccd1 vccd1 _1800_ sky130_fd_sc_hd__a221oi_1
X_5255_ _1034_ _0414_ _1729_ _1730_ _1731_ vssd1 vssd1 vccd1 vccd1 _1732_ sky130_fd_sc_hd__o2111a_1
X_4206_ egd_top.BitStream_buffer.BS_buffer\[36\] vssd1 vssd1 vccd1 vccd1 _0691_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5186_ _1408_ _3124_ _1660_ _1661_ _1662_ vssd1 vssd1 vccd1 vccd1 _1663_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _3077_ _3124_ _0618_ _0619_ _0621_ vssd1 vssd1 vccd1 vccd1 _0622_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4068_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _0554_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6658__146 clknet_1_1__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__inv_2
XFILLER_0_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3370_ net33 vssd1 vssd1 vccd1 vccd1 _2928_ sky130_fd_sc_hd__inv_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6693__22 clknet_1_1__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__inv_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _0566_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1519_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5942_ _2400_ _2396_ vssd1 vssd1 vccd1 vccd1 _2401_ sky130_fd_sc_hd__and2_1
XFILLER_0_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5873_ _0507_ _0691_ vssd1 vssd1 vccd1 vccd1 _2345_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4824_ _3206_ _3028_ vssd1 vssd1 vccd1 vccd1 _1304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4755_ _0711_ _0397_ _1233_ _1234_ _1235_ vssd1 vssd1 vccd1 vccd1 _1236_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3706_ _3090_ _3228_ vssd1 vssd1 vccd1 vccd1 _3240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4686_ _0611_ _3141_ vssd1 vssd1 vccd1 vccd1 _1167_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6425_ _2707_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] vssd1 vssd1 vccd1
+ vccd1 _2767_ sky130_fd_sc_hd__nand2_1
X_3637_ _3122_ _3167_ vssd1 vssd1 vccd1 vccd1 _3171_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6356_ _2690_ _2698_ vssd1 vssd1 vccd1 vccd1 _2699_ sky130_fd_sc_hd__nor2_1
X_3568_ egd_top.BitStream_buffer.BS_buffer\[67\] vssd1 vssd1 vccd1 vccd1 _3102_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5307_ _3133_ _3255_ vssd1 vssd1 vccd1 vccd1 _1783_ sky130_fd_sc_hd__nand2_1
X_6287_ _2635_ vssd1 vssd1 vccd1 vccd1 _0166_ sky130_fd_sc_hd__clkbuf_1
X_3499_ _3038_ _2933_ vssd1 vssd1 vccd1 vccd1 _3039_ sky130_fd_sc_hd__and2_1
X_5238_ _1592_ _0345_ _1714_ _0349_ vssd1 vssd1 vccd1 vccd1 _1715_ sky130_fd_sc_hd__o22ai_1
X_5169_ _0509_ _0589_ _0503_ _0592_ _1646_ vssd1 vssd1 vccd1 vccd1 _1647_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold6 egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _0890_ _0595_ _1022_ _0598_ vssd1 vssd1 vccd1 vccd1 _1023_ sky130_fd_sc_hd__o22ai_1
X_4471_ _3344_ _3310_ vssd1 vssd1 vccd1 vccd1 _0954_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3422_ _2975_ vssd1 vssd1 vccd1 vccd1 _2976_ sky130_fd_sc_hd__inv_2
X_6210_ net9 _3357_ net197 vssd1 vssd1 vccd1 vccd1 _2585_ sky130_fd_sc_hd__mux2_1
X_6141_ _2537_ _2529_ vssd1 vssd1 vccd1 vccd1 _2538_ sky130_fd_sc_hd__and2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _2490_ vssd1 vssd1 vccd1 vccd1 _0230_ sky130_fd_sc_hd__clkbuf_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5023_ _0498_ _0479_ vssd1 vssd1 vccd1 vccd1 _1502_ sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5925_ net3 _0552_ _2380_ vssd1 vssd1 vccd1 vccd1 _2389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5856_ _3120_ _0425_ vssd1 vssd1 vccd1 vccd1 _2328_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4807_ _3114_ _3119_ vssd1 vssd1 vccd1 vccd1 _1287_ sky130_fd_sc_hd__nand2_1
X_5787_ _3132_ _0646_ vssd1 vssd1 vccd1 vccd1 _2259_ sky130_fd_sc_hd__nand2_1
X_4738_ _0338_ _0380_ vssd1 vssd1 vccd1 vccd1 _1219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4669_ _1022_ _0595_ _1150_ _0598_ vssd1 vssd1 vccd1 vccd1 _1151_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6408_ _2688_ _2750_ vssd1 vssd1 vccd1 vccd1 _2751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6339_ egd_top.BitStream_buffer.BitStream_buffer_output\[3\] egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ _2013_ vssd1 vssd1 vccd1 vccd1 _2682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3971_ _2967_ vssd1 vssd1 vccd1 vccd1 _0457_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5710_ _3174_ _3337_ _2180_ _2181_ _2182_ vssd1 vssd1 vccd1 vccd1 _2183_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5641_ _2103_ _2106_ _2110_ _2114_ vssd1 vssd1 vccd1 vccd1 _2115_ sky130_fd_sc_hd__and4_1
XFILLER_0_38_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5572_ _2042_ _2043_ _2044_ _2045_ vssd1 vssd1 vccd1 vccd1 _2046_ sky130_fd_sc_hd__and4_1
X_4523_ _0862_ _0506_ _1003_ _1004_ _1005_ vssd1 vssd1 vccd1 vccd1 _1006_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_31_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4454_ _0802_ _3264_ _3236_ _3268_ vssd1 vssd1 vccd1 vccd1 _0937_ sky130_fd_sc_hd__o22ai_1
X_4385_ _0867_ _0496_ _0868_ vssd1 vssd1 vccd1 vccd1 _0869_ sky130_fd_sc_hd__o21ai_1
X_3405_ _2957_ vssd1 vssd1 vccd1 vccd1 _2959_ sky130_fd_sc_hd__buf_6
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ net5 _3095_ _2521_ vssd1 vssd1 vccd1 vccd1 _2526_ sky130_fd_sc_hd__mux2_1
X_6055_ _2478_ vssd1 vssd1 vccd1 vccd1 _0235_ sky130_fd_sc_hd__clkbuf_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _0416_ _0455_ vssd1 vssd1 vccd1 vccd1 _1485_ sky130_fd_sc_hd__nand2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6709__37 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__inv_2
X_6888_ net86 _0291_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_5908_ egd_top.BitStream_buffer.buffer_index\[4\] _3002_ vssd1 vssd1 vccd1 vccd1
+ _2377_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5839_ _0417_ _0327_ _0423_ _0331_ _2310_ vssd1 vssd1 vccd1 vccd1 _2311_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_63_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__2920_ clknet_0__2920_ vssd1 vssd1 vccd1 vccd1 clknet_1_1__leaf__2920_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4170_ _0652_ _0654_ vssd1 vssd1 vccd1 vccd1 _0655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6811_ net165 _0214_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[65\]
+ sky130_fd_sc_hd__dfxtp_1
X_3954_ _0439_ vssd1 vssd1 vccd1 vccd1 _0440_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3885_ _0370_ vssd1 vssd1 vccd1 vccd1 _0371_ sky130_fd_sc_hd__clkbuf_4
X_5624_ _2087_ _2091_ _2094_ _2097_ vssd1 vssd1 vccd1 vccd1 _2098_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5555_ _0926_ _3175_ _0578_ _3178_ vssd1 vssd1 vccd1 vccd1 _2029_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ _0388_ _0423_ vssd1 vssd1 vccd1 vccd1 _1961_ sky130_fd_sc_hd__nand2_1
X_4506_ _0703_ _0432_ _0400_ _0436_ _0988_ vssd1 vssd1 vccd1 vccd1 _0989_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4437_ _0638_ _3190_ _0919_ vssd1 vssd1 vccd1 vccd1 _0920_ sky130_fd_sc_hd__o21ai_1
X_4368_ _0848_ _0414_ _0849_ _0850_ _0851_ vssd1 vssd1 vccd1 vccd1 _0852_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_67_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6107_ net9 _0451_ _2485_ vssd1 vssd1 vccd1 vccd1 _2514_ sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _3192_ _3044_ vssd1 vssd1 vccd1 vccd1 _0783_ sky130_fd_sc_hd__nand2_1
X_6038_ _2466_ _2448_ vssd1 vssd1 vccd1 vccd1 _2467_ sky130_fd_sc_hd__and2_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3670_ _3203_ vssd1 vssd1 vccd1 vccd1 _3204_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5340_ _3313_ _3013_ vssd1 vssd1 vccd1 vccd1 _1816_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6612__103 clknet_1_0__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__inv_2
XFILLER_0_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5271_ _0475_ _0488_ _0479_ _0492_ _1747_ vssd1 vssd1 vccd1 vccd1 _1748_ sky130_fd_sc_hd__a221oi_1
X_4222_ _0700_ _0397_ _0702_ _0704_ _0706_ vssd1 vssd1 vccd1 vccd1 _0707_ sky130_fd_sc_hd__o2111a_1
X_4153_ _3050_ vssd1 vssd1 vccd1 vccd1 _0638_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _0569_ vssd1 vssd1 vccd1 vccd1 _0570_ sky130_fd_sc_hd__buf_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0__2922_ _2922_ vssd1 vssd1 vccd1 vccd1 clknet_0__2922_ sky130_fd_sc_hd__clkbuf_16
X_4986_ _1422_ _1433_ _1447_ _1464_ vssd1 vssd1 vccd1 vccd1 _1465_ sky130_fd_sc_hd__and4_1
X_3937_ egd_top.BitStream_buffer.BS_buffer\[57\] vssd1 vssd1 vccd1 vccd1 _0423_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ _3122_ _0325_ vssd1 vssd1 vccd1 vccd1 _0354_ sky130_fd_sc_hd__and2_1
X_5607_ _0412_ _0385_ _2080_ vssd1 vssd1 vccd1 vccd1 _2081_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3799_ _3328_ _3332_ vssd1 vssd1 vccd1 vccd1 _3333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5538_ egd_top.BitStream_buffer.BitStream_buffer_output\[4\] vssd1 vssd1 vccd1 vccd1
+ _2013_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5469_ _3202_ _3350_ vssd1 vssd1 vccd1 vccd1 _1944_ sky130_fd_sc_hd__or2_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 la_data_in_60_59[1] vssd1 vssd1 vccd1 vccd1 net18 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6635__125 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__inv_2
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4840_ _3327_ vssd1 vssd1 vccd1 vccd1 _1320_ sky130_fd_sc_hd__inv_2
X_4771_ _1251_ vssd1 vssd1 vccd1 vccd1 _1252_ sky130_fd_sc_hd__inv_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6510_ _2755_ _2786_ vssd1 vssd1 vccd1 vccd1 _2846_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3722_ _3254_ _3255_ vssd1 vssd1 vccd1 vccd1 _3256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6441_ _2743_ _2778_ _2782_ vssd1 vssd1 vccd1 vccd1 _2783_ sky130_fd_sc_hd__o21ai_1
X_3653_ _3186_ vssd1 vssd1 vccd1 vccd1 _3187_ sky130_fd_sc_hd__buf_6
X_6372_ _2650_ _2714_ vssd1 vssd1 vccd1 vccd1 _2715_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5323_ _0742_ _3218_ _0554_ _3221_ vssd1 vssd1 vccd1 vccd1 _1799_ sky130_fd_sc_hd__o22ai_1
X_3584_ _3095_ _3101_ _3102_ _3106_ _3117_ vssd1 vssd1 vccd1 vccd1 _3118_ sky130_fd_sc_hd__a221oi_1
X_5254_ _0767_ _0426_ vssd1 vssd1 vccd1 vccd1 _1731_ sky130_fd_sc_hd__or2_1
X_4205_ egd_top.BitStream_buffer.BS_buffer\[35\] vssd1 vssd1 vccd1 vccd1 _0690_ sky130_fd_sc_hd__inv_2
X_5185_ _1159_ _3141_ vssd1 vssd1 vccd1 vccd1 _1662_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4136_ _0620_ _3141_ vssd1 vssd1 vccd1 vccd1 _0621_ sky130_fd_sc_hd__or2_1
X_4067_ _0551_ _0552_ vssd1 vssd1 vccd1 vccd1 _0553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4969_ _3309_ _2998_ vssd1 vssd1 vccd1 vccd1 _1448_ sky130_fd_sc_hd__nand2_1
XFILLER_0_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_282 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5941_ net13 egd_top.BitStream_buffer.BS_buffer\[9\] _2380_ vssd1 vssd1 vccd1 vccd1
+ _2400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5872_ _0521_ _0487_ _0525_ _0491_ _2343_ vssd1 vssd1 vccd1 vccd1 _2344_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4823_ _3050_ _3184_ _3053_ _3187_ _1302_ vssd1 vssd1 vccd1 vccd1 _1303_ sky130_fd_sc_hd__a221oi_1
X_4754_ _0708_ _0408_ vssd1 vssd1 vccd1 vccd1 _1235_ sky130_fd_sc_hd__or2_1
XFILLER_0_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3705_ egd_top.BitStream_buffer.BS_buffer\[89\] vssd1 vssd1 vccd1 vccd1 _3239_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4685_ _3133_ _3069_ vssd1 vssd1 vccd1 vccd1 _1166_ sky130_fd_sc_hd__nand2_1
X_6424_ _2669_ _2700_ egd_top.BitStream_buffer.BitStream_buffer_output\[5\] vssd1
+ vssd1 vccd1 vccd1 _2766_ sky130_fd_sc_hd__o21ai_1
X_3636_ _3169_ vssd1 vssd1 vccd1 vccd1 _3170_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6355_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _2694_ _2697_ vssd1
+ vssd1 vccd1 vccd1 _2698_ sky130_fd_sc_hd__o21ai_1
X_3567_ _3100_ vssd1 vssd1 vccd1 vccd1 _3101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6286_ _2634_ _2372_ vssd1 vssd1 vccd1 vccd1 _2635_ sky130_fd_sc_hd__and2_1
X_5306_ _3128_ _3144_ vssd1 vssd1 vccd1 vccd1 _1782_ sky130_fd_sc_hd__nand2_1
X_5237_ egd_top.BitStream_buffer.BS_buffer\[46\] vssd1 vssd1 vccd1 vccd1 _1714_ sky130_fd_sc_hd__inv_2
X_3498_ net12 _3037_ _3007_ vssd1 vssd1 vccd1 vccd1 _3038_ sky130_fd_sc_hd__mux2_1
X_6664__151 clknet_1_1__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__inv_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5168_ _0867_ _0595_ _0516_ _0598_ vssd1 vssd1 vccd1 vccd1 _1646_ sky130_fd_sc_hd__o22ai_1
X_5099_ _1575_ _1576_ vssd1 vssd1 vccd1 vccd1 _1577_ sky130_fd_sc_hd__nand2_1
X_4119_ _0604_ vssd1 vssd1 vccd1 vccd1 _0605_ sky130_fd_sc_hd__buf_1
XFILLER_0_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold7 egd_top.BitStream_buffer.buffer_index\[4\] vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4470_ _3340_ _3335_ vssd1 vssd1 vccd1 vccd1 _0953_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3421_ _2950_ _2970_ vssd1 vssd1 vccd1 vccd1 _2975_ sky130_fd_sc_hd__nor2_1
X_6140_ net15 _3119_ _2521_ vssd1 vssd1 vccd1 vccd1 _2537_ sky130_fd_sc_hd__mux2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _2489_ _2475_ vssd1 vssd1 vccd1 vccd1 _2490_ sky130_fd_sc_hd__and2_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5022_ _1497_ _0472_ _1498_ _1500_ vssd1 vssd1 vccd1 vccd1 _1501_ sky130_fd_sc_hd__o211a_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5924_ _2388_ vssd1 vssd1 vccd1 vccd1 _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5855_ _0419_ _3076_ vssd1 vssd1 vccd1 vccd1 _2327_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _3255_ _3068_ _3247_ _3075_ _1285_ vssd1 vssd1 vccd1 vccd1 _1286_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5786_ _3127_ _3259_ vssd1 vssd1 vccd1 vccd1 _2258_ sky130_fd_sc_hd__nand2_1
X_4737_ _0334_ _0389_ vssd1 vssd1 vccd1 vccd1 _1218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4668_ _0489_ vssd1 vssd1 vccd1 vccd1 _1150_ sky130_fd_sc_hd__inv_2
X_3619_ _2954_ _3087_ vssd1 vssd1 vccd1 vccd1 _3153_ sky130_fd_sc_hd__nor2_4
X_6407_ _2661_ _2749_ vssd1 vssd1 vccd1 vccd1 _2750_ sky130_fd_sc_hd__nand2_1
X_4599_ egd_top.BitStream_buffer.BS_buffer\[107\] vssd1 vssd1 vccd1 vccd1 _1081_ sky130_fd_sc_hd__inv_2
X_6338_ _2680_ _2651_ vssd1 vssd1 vccd1 vccd1 _2681_ sky130_fd_sc_hd__nand2_2
X_6269_ _2623_ vssd1 vssd1 vccd1 vccd1 _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3970_ _0455_ vssd1 vssd1 vccd1 vccd1 _0456_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5640_ _0323_ _0523_ _0329_ _0527_ _2113_ vssd1 vssd1 vccd1 vccd1 _2114_ sky130_fd_sc_hd__a221oi_1
X_5571_ _3257_ _3278_ vssd1 vssd1 vccd1 vccd1 _2045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4522_ _0468_ _0518_ vssd1 vssd1 vccd1 vccd1 _1005_ sky130_fd_sc_hd__or2_1
X_4453_ _0932_ _0933_ _0934_ _0935_ vssd1 vssd1 vccd1 vccd1 _0936_ sky130_fd_sc_hd__and4_1
X_3404_ egd_top.BitStream_buffer.pc_previous\[0\] _2957_ vssd1 vssd1 vccd1 vccd1 _2958_
+ sky130_fd_sc_hd__or2_1
X_4384_ _0498_ _0515_ vssd1 vssd1 vccd1 vccd1 _0868_ sky130_fd_sc_hd__nand2_1
X_6123_ _2525_ vssd1 vssd1 vccd1 vccd1 _0214_ sky130_fd_sc_hd__clkbuf_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _2477_ _2475_ vssd1 vssd1 vccd1 vccd1 _2478_ sky130_fd_sc_hd__and2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _0708_ _0397_ _1481_ _1482_ _1483_ vssd1 vssd1 vccd1 vccd1 _1484_ sky130_fd_sc_hd__o2111a_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5907_ _2376_ vssd1 vssd1 vccd1 vccd1 _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6887_ net85 _0290_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _2308_ _2309_ vssd1 vssd1 vccd1 vccd1 _2310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5769_ _0468_ _0560_ _2239_ _2240_ _2241_ vssd1 vssd1 vccd1 vccd1 _2242_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6810_ net164 _0213_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[66\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3953_ _3109_ _0395_ vssd1 vssd1 vccd1 vccd1 _0439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3884_ _3103_ _0325_ vssd1 vssd1 vccd1 vccd1 _0370_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5623_ _3076_ _0449_ _3085_ _0453_ _2096_ vssd1 vssd1 vccd1 vccd1 _2097_ sky130_fd_sc_hd__a221oi_1
X_5554_ _2016_ _2019_ _2023_ _2027_ vssd1 vssd1 vccd1 vccd1 _2028_ sky130_fd_sc_hd__and4_1
X_5485_ _0329_ _0362_ _0376_ _0366_ _1959_ vssd1 vssd1 vccd1 vccd1 _1960_ sky130_fd_sc_hd__a221oi_1
X_4505_ _0986_ _0440_ _0987_ vssd1 vssd1 vccd1 vccd1 _0988_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4436_ _3192_ _3047_ vssd1 vssd1 vccd1 vccd1 _0919_ sky130_fd_sc_hd__nand2_1
X_4367_ _0412_ _0426_ vssd1 vssd1 vccd1 vccd1 _0851_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6106_ _2513_ vssd1 vssd1 vccd1 vccd1 _0219_ sky130_fd_sc_hd__clkbuf_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _3031_ _3170_ _3034_ _3173_ _0781_ vssd1 vssd1 vccd1 vccd1 _0782_ sky130_fd_sc_hd__a221oi_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ net15 _0356_ _2451_ vssd1 vssd1 vccd1 vccd1 _2466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5270_ _0995_ _0496_ _1746_ vssd1 vssd1 vccd1 vccd1 _1747_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4221_ _0705_ _0408_ vssd1 vssd1 vccd1 vccd1 _0706_ sky130_fd_sc_hd__or2_1
X_4152_ _3016_ _3198_ _3019_ _3201_ _0636_ vssd1 vssd1 vccd1 vccd1 _0637_ sky130_fd_sc_hd__a221oi_1
X_4083_ _3090_ _0542_ vssd1 vssd1 vccd1 vccd1 _0569_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__2921_ _2921_ vssd1 vssd1 vccd1 vccd1 clknet_0__2921_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4985_ _1451_ _1455_ _1460_ _1463_ vssd1 vssd1 vccd1 vccd1 _1464_ sky130_fd_sc_hd__and4_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ _0420_ _0421_ vssd1 vssd1 vccd1 vccd1 _0422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3867_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0353_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5606_ _0387_ _0421_ vssd1 vssd1 vccd1 vccd1 _2080_ sky130_fd_sc_hd__nand2_1
X_3798_ _3330_ _3331_ vssd1 vssd1 vccd1 vccd1 _3332_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5537_ _1950_ _2010_ _2011_ vssd1 vssd1 vccd1 vccd1 _2012_ sky130_fd_sc_hd__nand3_1
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5468_ _3344_ _3010_ vssd1 vssd1 vccd1 vccd1 _1943_ sky130_fd_sc_hd__nand2_1
X_5399_ _1873_ _1874_ vssd1 vssd1 vccd1 vccd1 _1875_ sky130_fd_sc_hd__nand2_1
X_4419_ _3156_ _3068_ _3144_ _3075_ _0901_ vssd1 vssd1 vccd1 vccd1 _0902_ sky130_fd_sc_hd__a221oi_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 la_data_in_65 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__buf_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4770_ _0478_ _0525_ _0481_ _0359_ vssd1 vssd1 vccd1 vccd1 _1251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3721_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _3255_ sky130_fd_sc_hd__clkbuf_4
X_6440_ _2779_ _2780_ _2781_ vssd1 vssd1 vccd1 vccd1 _2782_ sky130_fd_sc_hd__o21ai_1
X_3652_ _3185_ vssd1 vssd1 vccd1 vccd1 _3186_ sky130_fd_sc_hd__clkbuf_2
X_6371_ _2713_ vssd1 vssd1 vccd1 vccd1 _2714_ sky130_fd_sc_hd__inv_2
X_3583_ _3108_ _3111_ _3116_ vssd1 vssd1 vccd1 vccd1 _3117_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5322_ _3044_ _3198_ _3047_ _3201_ _1797_ vssd1 vssd1 vccd1 vccd1 _1798_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5253_ _0420_ _3102_ vssd1 vssd1 vccd1 vccd1 _1730_ sky130_fd_sc_hd__nand2_1
X_4204_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _0689_ sky130_fd_sc_hd__clkbuf_4
X_5184_ _3133_ _3149_ vssd1 vssd1 vccd1 vccd1 _1661_ sky130_fd_sc_hd__nand2_1
X_4135_ _3134_ vssd1 vssd1 vccd1 vccd1 _0620_ sky130_fd_sc_hd__inv_2
X_4066_ egd_top.BitStream_buffer.BS_buffer\[4\] vssd1 vssd1 vccd1 vccd1 _0552_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _1435_ _1440_ _1443_ _1446_ vssd1 vssd1 vccd1 vccd1 _1447_ sky130_fd_sc_hd__and4_1
XFILLER_0_80_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3919_ _0403_ _0404_ vssd1 vssd1 vccd1 vccd1 _0405_ sky130_fd_sc_hd__nand2_1
X_4899_ _0468_ _0496_ _1378_ vssd1 vssd1 vccd1 vccd1 _1379_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6569_ _2901_ _2959_ vssd1 vssd1 vccd1 vccd1 _2902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6641__130 clknet_1_0__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__inv_2
XFILLER_0_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5940_ _2399_ vssd1 vssd1 vccd1 vccd1 _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5871_ _1619_ _0495_ _2342_ vssd1 vssd1 vccd1 vccd1 _2343_ sky130_fd_sc_hd__o21ai_1
X_4822_ _0578_ _3190_ _1301_ vssd1 vssd1 vccd1 vccd1 _1302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4753_ _0403_ _0423_ vssd1 vssd1 vccd1 vccd1 _1234_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3704_ _3237_ vssd1 vssd1 vccd1 vccd1 _3238_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6423_ _2761_ _2764_ vssd1 vssd1 vccd1 vccd1 _2765_ sky130_fd_sc_hd__nand2_1
X_4684_ _3128_ _3085_ vssd1 vssd1 vccd1 vccd1 _1165_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3635_ _3168_ vssd1 vssd1 vccd1 vccd1 _3169_ sky130_fd_sc_hd__buf_1
XFILLER_0_11_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6354_ _2696_ _2693_ _1157_ vssd1 vssd1 vccd1 vccd1 _2697_ sky130_fd_sc_hd__nand3_1
X_3566_ _3099_ vssd1 vssd1 vccd1 vccd1 _3100_ sky130_fd_sc_hd__buf_1
X_6285_ net12 _3225_ _2613_ vssd1 vssd1 vccd1 vccd1 _2634_ sky130_fd_sc_hd__mux2_1
X_3497_ egd_top.BitStream_buffer.BS_buffer\[122\] vssd1 vssd1 vccd1 vccd1 _3037_ sky130_fd_sc_hd__clkbuf_4
X_5305_ _3161_ _3101_ _3156_ _3106_ _1780_ vssd1 vssd1 vccd1 vccd1 _1781_ sky130_fd_sc_hd__a221oi_2
X_5236_ _0433_ _0328_ _0404_ _0332_ _1712_ vssd1 vssd1 vccd1 vccd1 _1713_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5167_ _0750_ _0576_ _0568_ _0580_ _1644_ vssd1 vssd1 vccd1 vccd1 _1645_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5098_ _3330_ _3297_ vssd1 vssd1 vccd1 vccd1 _1576_ sky130_fd_sc_hd__nand2_1
X_4118_ _0603_ _2965_ _3062_ _3063_ vssd1 vssd1 vccd1 vccd1 _0604_ sky130_fd_sc_hd__and4b_1
X_4049_ egd_top.BitStream_buffer.BS_buffer\[28\] vssd1 vssd1 vccd1 vccd1 _0535_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_275 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 _2450_ vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3420_ _2968_ _2970_ _2973_ vssd1 vssd1 vccd1 vccd1 _2974_ sky130_fd_sc_hd__nand3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ net6 _0443_ _2486_ vssd1 vssd1 vccd1 vccd1 _2489_ sky130_fd_sc_hd__mux2_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _1499_ vssd1 vssd1 vccd1 vccd1 _1500_ sky130_fd_sc_hd__inv_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2927_ clknet_0__2927_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2927_
+ sky130_fd_sc_hd__clkbuf_16
X_5923_ _2387_ _3042_ vssd1 vssd1 vccd1 vccd1 _2388_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5854_ _0415_ _3134_ vssd1 vssd1 vccd1 vccd1 _2326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4805_ _1159_ _3084_ _1284_ _3092_ vssd1 vssd1 vccd1 vccd1 _1285_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5785_ _3255_ _3100_ _3247_ _3105_ _2256_ vssd1 vssd1 vccd1 vccd1 _2257_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4736_ _1173_ _1185_ _1199_ _1216_ vssd1 vssd1 vccd1 vccd1 _1217_ sky130_fd_sc_hd__and4_1
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4667_ _0742_ _0576_ _0541_ _0580_ _1148_ vssd1 vssd1 vccd1 vccd1 _1149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3618_ _3151_ vssd1 vssd1 vccd1 vccd1 _3152_ sky130_fd_sc_hd__buf_4
X_6406_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2749_ sky130_fd_sc_hd__nand2_1
X_4598_ _3341_ _3321_ _3347_ _3324_ _1079_ vssd1 vssd1 vccd1 vccd1 _1080_ sky130_fd_sc_hd__a221oi_1
X_6337_ _2678_ _2679_ vssd1 vssd1 vccd1 vccd1 _2680_ sky130_fd_sc_hd__nand2_1
X_3549_ _3082_ _3065_ vssd1 vssd1 vccd1 vccd1 _3083_ sky130_fd_sc_hd__nand2_1
X_6268_ _2622_ _2581_ vssd1 vssd1 vccd1 vccd1 _2623_ sky130_fd_sc_hd__and2_1
X_5219_ _3016_ _3303_ _3019_ _3307_ _1695_ vssd1 vssd1 vccd1 vccd1 _1696_ sky130_fd_sc_hd__a221oi_1
X_6199_ _2577_ vssd1 vssd1 vccd1 vccd1 _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6735__61 clknet_1_0__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__inv_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6750__75 clknet_1_1__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__inv_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5570_ _3253_ _3286_ vssd1 vssd1 vccd1 vccd1 _2044_ sky130_fd_sc_hd__nand2_1
X_4521_ _0512_ _0503_ vssd1 vssd1 vccd1 vccd1 _1004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4452_ _3258_ _3265_ vssd1 vssd1 vccd1 vccd1 _0935_ sky130_fd_sc_hd__nand2_1
X_3403_ _2955_ _2956_ vssd1 vssd1 vccd1 vccd1 _2957_ sky130_fd_sc_hd__nand2_1
X_4383_ _0513_ vssd1 vssd1 vccd1 vccd1 _0867_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _2524_ _2502_ vssd1 vssd1 vccd1 vccd1 _2525_ sky130_fd_sc_hd__and2_1
X_6053_ net10 _0376_ _2450_ vssd1 vssd1 vccd1 vccd1 _2477_ sky130_fd_sc_hd__mux2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _0981_ _0408_ vssd1 vssd1 vccd1 vccd1 _1483_ sky130_fd_sc_hd__or2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5906_ _3004_ _2372_ _2375_ vssd1 vssd1 vccd1 vccd1 _2376_ sky130_fd_sc_hd__and3_1
X_6886_ net84 _0289_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_5837_ _0337_ _0400_ vssd1 vssd1 vccd1 vccd1 _2309_ sky130_fd_sc_hd__nand2_1
X_5768_ _0734_ _0569_ vssd1 vssd1 vccd1 vccd1 _2241_ sky130_fd_sc_hd__or2_1
X_4719_ _3309_ _0674_ vssd1 vssd1 vccd1 vccd1 _1200_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5699_ _3308_ _3025_ vssd1 vssd1 vccd1 vccd1 _2172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6740_ clknet_1_0__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2927_ sky130_fd_sc_hd__buf_1
X_3952_ _0437_ vssd1 vssd1 vccd1 vccd1 _0438_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3883_ _0368_ vssd1 vssd1 vccd1 vccd1 _0369_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_301 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5622_ _0764_ _0457_ _2095_ vssd1 vssd1 vccd1 vccd1 _2096_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5553_ _3225_ _3147_ _3232_ _3151_ _2026_ vssd1 vssd1 vccd1 vccd1 _2027_ sky130_fd_sc_hd__a221oi_1
X_4504_ _0442_ _0404_ vssd1 vssd1 vccd1 vccd1 _0987_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5484_ _1592_ _0369_ _1958_ vssd1 vssd1 vccd1 vccd1 _1959_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4435_ _3034_ _3170_ _3037_ _3173_ _0917_ vssd1 vssd1 vccd1 vccd1 _0918_ sky130_fd_sc_hd__a221oi_1
X_4366_ _0420_ _0447_ vssd1 vssd1 vccd1 vccd1 _0850_ sky130_fd_sc_hd__nand2_1
X_6105_ _2512_ _2502_ vssd1 vssd1 vccd1 vccd1 _2513_ sky130_fd_sc_hd__and2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _0628_ _3176_ _0780_ _3179_ vssd1 vssd1 vccd1 vccd1 _0781_ sky130_fd_sc_hd__o22ai_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _2465_ vssd1 vssd1 vccd1 vccd1 _0241_ sky130_fd_sc_hd__clkbuf_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6869_ net67 _0272_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4220_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0705_ sky130_fd_sc_hd__inv_2
X_4151_ _0634_ _3204_ _0635_ vssd1 vssd1 vccd1 vccd1 _0636_ sky130_fd_sc_hd__o21ai_1
X_4082_ egd_top.BitStream_buffer.BS_buffer\[9\] vssd1 vssd1 vccd1 vccd1 _0568_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_0__2920_ _2920_ vssd1 vssd1 vccd1 vccd1 clknet_0__2920_ sky130_fd_sc_hd__clkbuf_16
X_4984_ _3016_ _3356_ _3019_ _3360_ _1462_ vssd1 vssd1 vccd1 vccd1 _1463_ sky130_fd_sc_hd__a221oi_2
X_3935_ egd_top.BitStream_buffer.BS_buffer\[58\] vssd1 vssd1 vccd1 vccd1 _0421_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3866_ _0351_ vssd1 vssd1 vccd1 vccd1 _0352_ sky130_fd_sc_hd__clkbuf_4
X_5605_ _0376_ _0361_ _0380_ _0365_ _2078_ vssd1 vssd1 vccd1 vccd1 _2079_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3797_ egd_top.BitStream_buffer.BS_buffer\[98\] vssd1 vssd1 vccd1 vccd1 _3331_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5536_ _0606_ egd_top.BitStream_buffer.BS_buffer\[11\] vssd1 vssd1 vccd1 vccd1 _2011_
+ sky130_fd_sc_hd__nand2_1
X_5467_ _3340_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _1942_
+ sky130_fd_sc_hd__nand2_1
X_4418_ _0764_ _3084_ _0900_ _3092_ vssd1 vssd1 vccd1 vccd1 _0901_ sky130_fd_sc_hd__o22ai_1
X_5398_ _0534_ _0353_ vssd1 vssd1 vccd1 vccd1 _1874_ sky130_fd_sc_hd__nand2_1
X_4349_ egd_top.BitStream_buffer.BS_buffer\[39\] vssd1 vssd1 vccd1 vccd1 _0833_ sky130_fd_sc_hd__inv_2
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6019_ net6 _0363_ _2451_ vssd1 vssd1 vccd1 vccd1 _2454_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3720_ _3253_ vssd1 vssd1 vccd1 vccd1 _3254_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3651_ _3090_ _3167_ vssd1 vssd1 vccd1 vccd1 _3185_ sky130_fd_sc_hd__and2_1
X_6370_ _2712_ _2959_ vssd1 vssd1 vccd1 vccd1 _2713_ sky130_fd_sc_hd__nand2_2
X_3582_ _3114_ _3115_ vssd1 vssd1 vccd1 vccd1 _3116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5321_ _1174_ _3204_ _1796_ vssd1 vssd1 vccd1 vccd1 _1797_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5252_ _0416_ _3115_ vssd1 vssd1 vccd1 vccd1 _1729_ sky130_fd_sc_hd__nand2_1
X_4203_ _0686_ _0687_ vssd1 vssd1 vccd1 vccd1 _0688_ sky130_fd_sc_hd__nor2_1
X_5183_ _3128_ _3156_ vssd1 vssd1 vccd1 vccd1 _1660_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4134_ _3133_ _3119_ vssd1 vssd1 vccd1 vccd1 _0619_ sky130_fd_sc_hd__nand2_1
X_4065_ _0550_ vssd1 vssd1 vccd1 vccd1 _0551_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _3347_ _3281_ _3345_ _3285_ _1445_ vssd1 vssd1 vccd1 vccd1 _1446_ sky130_fd_sc_hd__a221oi_1
X_3918_ egd_top.BitStream_buffer.BS_buffer\[52\] vssd1 vssd1 vccd1 vccd1 _0404_ sky130_fd_sc_hd__clkbuf_4
X_4898_ _0498_ _0475_ vssd1 vssd1 vccd1 vccd1 _1378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3849_ egd_top.BitStream_buffer.BS_buffer\[41\] vssd1 vssd1 vccd1 vccd1 _0335_ sky130_fd_sc_hd__buf_4
XFILLER_0_46_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6568_ _2900_ vssd1 vssd1 vccd1 vccd1 _2901_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _1992_ _1993_ vssd1 vssd1 vccd1 vccd1 _1994_ sky130_fd_sc_hd__nand2_1
X_6499_ _1406_ _2806_ vssd1 vssd1 vccd1 vccd1 _2835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5870_ _0497_ _0363_ vssd1 vssd1 vccd1 vccd1 _2342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4821_ _3192_ _0607_ vssd1 vssd1 vccd1 vccd1 _1301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4752_ _0399_ _0411_ vssd1 vssd1 vccd1 vccd1 _1233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3703_ _3082_ _3228_ vssd1 vssd1 vccd1 vccd1 _3237_ sky130_fd_sc_hd__nand2_1
X_4683_ _3119_ _3101_ _3076_ _3106_ _1163_ vssd1 vssd1 vccd1 vccd1 _1164_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_50_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6422_ _2762_ _2763_ vssd1 vssd1 vccd1 vccd1 _2764_ sky130_fd_sc_hd__nand2_1
X_3634_ _3131_ _3167_ vssd1 vssd1 vccd1 vccd1 _3168_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6353_ _2695_ vssd1 vssd1 vccd1 vccd1 _2696_ sky130_fd_sc_hd__inv_2
X_3565_ _3098_ _3064_ vssd1 vssd1 vccd1 vccd1 _3099_ sky130_fd_sc_hd__and2_1
X_6684__14 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__inv_2
X_3496_ _3036_ vssd1 vssd1 vccd1 vccd1 _0304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6284_ _2633_ vssd1 vssd1 vccd1 vccd1 _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5304_ _0611_ _3111_ _1779_ vssd1 vssd1 vccd1 vccd1 _1780_ sky130_fd_sc_hd__o21ai_1
X_5235_ _1710_ _1711_ vssd1 vssd1 vccd1 vccd1 _1712_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _0559_ _0584_ vssd1 vssd1 vccd1 vccd1 _1644_ sky130_fd_sc_hd__or2_1
X_6625__115 clknet_1_0__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__inv_2
X_5097_ _3326_ _3304_ vssd1 vssd1 vccd1 vccd1 _1575_ sky130_fd_sc_hd__nand2_1
X_4117_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] egd_top.BitStream_buffer.pc\[1\]
+ _2962_ _0543_ vssd1 vssd1 vccd1 vccd1 _0603_ sky130_fd_sc_hd__o41a_1
X_4048_ _0533_ vssd1 vssd1 vccd1 vccd1 _0534_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5999_ _2439_ _2423_ vssd1 vssd1 vccd1 vccd1 _2440_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _0478_ egd_top.BitStream_buffer.BS_buffer\[33\] _0481_ _0689_ vssd1 vssd1
+ vccd1 vccd1 _1499_ sky130_fd_sc_hd__a22o_1
X_6648__137 clknet_1_1__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__inv_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2926_ clknet_0__2926_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2926_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ net4 _0581_ _2380_ vssd1 vssd1 vccd1 vccd1 _2387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5853_ _0903_ _0396_ _2322_ _2323_ _2324_ vssd1 vssd1 vccd1 vccd1 _2325_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5784_ _1159_ _3110_ _2255_ vssd1 vssd1 vccd1 vccd1 _2256_ sky130_fd_sc_hd__o21ai_1
X_4804_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _1284_ sky130_fd_sc_hd__inv_2
X_4735_ _1203_ _1207_ _1212_ _1215_ vssd1 vssd1 vccd1 vccd1 _1216_ sky130_fd_sc_hd__and4_1
XFILLER_0_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4666_ _0554_ _0584_ vssd1 vssd1 vccd1 vccd1 _1148_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4597_ _1077_ _1078_ vssd1 vssd1 vccd1 vccd1 _1079_ sky130_fd_sc_hd__nand2_1
X_3617_ _3150_ vssd1 vssd1 vccd1 vccd1 _3151_ sky130_fd_sc_hd__clkbuf_2
X_6405_ _2692_ _2693_ _2747_ vssd1 vssd1 vccd1 vccd1 _2748_ sky130_fd_sc_hd__nand3_1
X_3548_ _3081_ vssd1 vssd1 vccd1 vccd1 _3082_ sky130_fd_sc_hd__clkbuf_4
X_6336_ _1029_ egd_top.BitStream_buffer.BitStream_buffer_output\[11\] egd_top.BitStream_buffer.BitStream_buffer_output\[13\]
+ vssd1 vssd1 vccd1 vccd1 _2679_ sky130_fd_sc_hd__a21oi_1
X_3479_ _3023_ _2933_ vssd1 vssd1 vccd1 vccd1 _3024_ sky130_fd_sc_hd__and2_1
X_6267_ net3 _0646_ _2613_ vssd1 vssd1 vccd1 vccd1 _2622_ sky130_fd_sc_hd__mux2_1
X_5218_ _1693_ _1694_ vssd1 vssd1 vccd1 vccd1 _1695_ sky130_fd_sc_hd__nand2_1
X_6198_ _2576_ _2554_ vssd1 vssd1 vccd1 vccd1 _2577_ sky130_fd_sc_hd__and2_1
X_5149_ _0508_ _0521_ vssd1 vssd1 vccd1 vccd1 _1627_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4520_ _0508_ _0475_ vssd1 vssd1 vccd1 vccd1 _1003_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4451_ _3254_ _3251_ vssd1 vssd1 vccd1 vccd1 _0934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3402_ net17 vssd1 vssd1 vccd1 vccd1 _2956_ sky130_fd_sc_hd__inv_2
X_4382_ _0862_ _0472_ _0863_ _0865_ vssd1 vssd1 vccd1 vccd1 _0866_ sky130_fd_sc_hd__o211a_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ net6 _3115_ _2521_ vssd1 vssd1 vccd1 vccd1 _2524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _2476_ vssd1 vssd1 vccd1 vccd1 _0236_ sky130_fd_sc_hd__clkbuf_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5003_ _0403_ _0411_ vssd1 vssd1 vccd1 vccd1 _1482_ sky130_fd_sc_hd__nand2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5905_ _3003_ _2971_ vssd1 vssd1 vccd1 vccd1 _2375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6885_ net83 _0288_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_5836_ _0333_ _0701_ vssd1 vssd1 vccd1 vccd1 _2308_ sky130_fd_sc_hd__nand2_1
X_5767_ _0565_ _0515_ vssd1 vssd1 vccd1 vccd1 _2240_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4718_ _1187_ _1192_ _1195_ _1198_ vssd1 vssd1 vccd1 vccd1 _1199_ sky130_fd_sc_hd__and4_1
X_5698_ _2160_ _2165_ _2168_ _2170_ vssd1 vssd1 vccd1 vccd1 _2171_ sky130_fd_sc_hd__and4_1
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4649_ _0508_ _0479_ vssd1 vssd1 vccd1 vccd1 _1131_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6319_ egd_top.BitStream_buffer.BitStream_buffer_output\[7\] _2661_ vssd1 vssd1 vccd1
+ vccd1 _2662_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3951_ egd_top.BitStream_buffer.BS_buffer\[48\] vssd1 vssd1 vccd1 vccd1 _0437_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3882_ _3098_ _0325_ vssd1 vssd1 vccd1 vccd1 _0368_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5621_ _0459_ _3057_ vssd1 vssd1 vccd1 vccd1 _2095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5552_ _2024_ _2025_ vssd1 vssd1 vccd1 vccd1 _2026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4503_ egd_top.BitStream_buffer.BS_buffer\[51\] vssd1 vssd1 vccd1 vccd1 _0986_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483_ _0371_ _0389_ vssd1 vssd1 vccd1 vccd1 _1958_ sky130_fd_sc_hd__nand2_1
X_4434_ _0780_ _3176_ _0916_ _3179_ vssd1 vssd1 vccd1 vccd1 _0917_ sky130_fd_sc_hd__o22ai_1
X_4365_ _0416_ _0421_ vssd1 vssd1 vccd1 vccd1 _0849_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6104_ net10 _0447_ _2485_ vssd1 vssd1 vccd1 vccd1 _2512_ sky130_fd_sc_hd__mux2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _2464_ _2448_ vssd1 vssd1 vccd1 vccd1 _2465_ sky130_fd_sc_hd__and2_1
X_4296_ egd_top.BitStream_buffer.BS_buffer\[119\] vssd1 vssd1 vccd1 vccd1 _0780_ sky130_fd_sc_hd__inv_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6868_ net66 _0271_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5819_ _3308_ _3028_ vssd1 vssd1 vccd1 vccd1 _2291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6799_ net153 _0202_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[77\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4150_ _3206_ _3013_ vssd1 vssd1 vccd1 vccd1 _0635_ sky130_fd_sc_hd__nand2_1
X_4081_ _0566_ egd_top.BitStream_buffer.BS_buffer\[8\] vssd1 vssd1 vccd1 vccd1 _0567_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4983_ _0628_ _3363_ _1461_ vssd1 vssd1 vccd1 vccd1 _1462_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3934_ _0419_ vssd1 vssd1 vccd1 vccd1 _0420_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3865_ _3131_ _0325_ vssd1 vssd1 vccd1 vccd1 _0351_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5604_ _1714_ _0368_ _2077_ vssd1 vssd1 vccd1 vccd1 _2078_ sky130_fd_sc_hd__o21ai_1
X_6584_ clknet_1_1__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2915_ sky130_fd_sc_hd__buf_1
X_3796_ _3329_ vssd1 vssd1 vccd1 vccd1 _3330_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5535_ _1980_ _1996_ _2009_ vssd1 vssd1 vccd1 vccd1 _2010_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ _3304_ _3321_ _3353_ _3324_ _1940_ vssd1 vssd1 vccd1 vccd1 _1941_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4417_ _3161_ vssd1 vssd1 vccd1 vccd1 _0900_ sky130_fd_sc_hd__inv_2
X_5397_ _0530_ _0356_ vssd1 vssd1 vccd1 vccd1 _1873_ sky130_fd_sc_hd__nand2_1
X_4348_ _0376_ _0328_ _0380_ _0332_ _0831_ vssd1 vssd1 vccd1 vccd1 _0832_ sky130_fd_sc_hd__a221oi_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ _3056_ _0762_ _0763_ vssd1 vssd1 vccd1 vccd1 _0296_ sky130_fd_sc_hd__o21a_1
X_6018_ _2453_ vssd1 vssd1 vccd1 vccd1 _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ _3183_ vssd1 vssd1 vccd1 vccd1 _3184_ sky130_fd_sc_hd__buf_4
X_3581_ egd_top.BitStream_buffer.BS_buffer\[65\] vssd1 vssd1 vccd1 vccd1 _3115_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _3206_ _3040_ vssd1 vssd1 vccd1 vccd1 _1796_ sky130_fd_sc_hd__nand2_1
X_5251_ _0981_ _0397_ _1725_ _1726_ _1727_ vssd1 vssd1 vccd1 vccd1 _1728_ sky130_fd_sc_hd__o2111a_1
X_4202_ _0352_ _0356_ _0355_ _0339_ vssd1 vssd1 vccd1 vccd1 _0687_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5182_ _3069_ _3101_ _3161_ _3106_ _1658_ vssd1 vssd1 vccd1 vccd1 _1659_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4133_ _3128_ _3136_ vssd1 vssd1 vccd1 vccd1 _0618_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _3126_ _0543_ vssd1 vssd1 vccd1 vccd1 _0550_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6605__97 clknet_1_0__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__inv_2
XFILLER_0_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4966_ _1320_ _3289_ _1444_ _3293_ vssd1 vssd1 vccd1 vccd1 _1445_ sky130_fd_sc_hd__o22ai_1
X_4897_ _1373_ _0472_ _1374_ _1376_ vssd1 vssd1 vccd1 vccd1 _1377_ sky130_fd_sc_hd__o211a_1
X_3917_ _0402_ vssd1 vssd1 vccd1 vccd1 _0403_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3848_ _0333_ vssd1 vssd1 vccd1 vccd1 _0334_ sky130_fd_sc_hd__buf_4
X_6636_ clknet_1_1__leaf__2914_ vssd1 vssd1 vccd1 vccd1 _2919_ sky130_fd_sc_hd__buf_1
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6567_ _2899_ _2707_ vssd1 vssd1 vccd1 vccd1 _2900_ sky130_fd_sc_hd__nand2_1
X_3779_ _3312_ vssd1 vssd1 vccd1 vccd1 _3313_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5518_ _0534_ _0356_ vssd1 vssd1 vccd1 vccd1 _1993_ sky130_fd_sc_hd__nand2_1
X_6498_ egd_top.BitStream_buffer.BitStream_buffer_output\[9\] _2805_ vssd1 vssd1 vccd1
+ vccd1 _2834_ sky130_fd_sc_hd__nor2_1
X_5449_ _3250_ _3278_ vssd1 vssd1 vccd1 vccd1 _1924_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ _3044_ _3170_ _3047_ _3173_ _1299_ vssd1 vssd1 vccd1 vccd1 _1300_ sky130_fd_sc_hd__a221oi_1
X_4751_ _1221_ _1225_ _1228_ _1231_ vssd1 vssd1 vccd1 vccd1 _1232_ sky130_fd_sc_hd__and4_1
XFILLER_0_83_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3702_ egd_top.BitStream_buffer.BS_buffer\[88\] vssd1 vssd1 vccd1 vccd1 _3236_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4682_ _3137_ _3111_ _1162_ vssd1 vssd1 vccd1 vccd1 _1163_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6421_ _2707_ _2132_ vssd1 vssd1 vccd1 vccd1 _2763_ sky130_fd_sc_hd__nand2_1
X_3633_ _3166_ vssd1 vssd1 vccd1 vccd1 _3167_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3564_ _3097_ _3058_ vssd1 vssd1 vccd1 vccd1 _3098_ sky130_fd_sc_hd__nor2_4
X_6352_ _2691_ _2666_ vssd1 vssd1 vccd1 vccd1 _2695_ sky130_fd_sc_hd__nand2_1
X_3495_ _3035_ _2933_ vssd1 vssd1 vccd1 vccd1 _3036_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6283_ _2632_ _2372_ vssd1 vssd1 vccd1 vccd1 _2633_ sky130_fd_sc_hd__and2_1
X_5303_ _3114_ _3069_ vssd1 vssd1 vccd1 vccd1 _1779_ sky130_fd_sc_hd__nand2_1
X_5234_ _0338_ _0443_ vssd1 vssd1 vccd1 vccd1 _1711_ sky130_fd_sc_hd__nand2_1
X_5165_ _0728_ _0561_ _1640_ _1641_ _1642_ vssd1 vssd1 vccd1 vccd1 _1643_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4116_ _0466_ _0539_ _0601_ vssd1 vssd1 vccd1 vccd1 _0602_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5096_ _3013_ _3303_ _3016_ _3307_ _1573_ vssd1 vssd1 vccd1 vccd1 _1574_ sky130_fd_sc_hd__a221oi_1
X_4047_ _3158_ _0470_ vssd1 vssd1 vccd1 vccd1 _0533_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5998_ net11 _0482_ _2415_ vssd1 vssd1 vccd1 vccd1 _2439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4949_ _3206_ _3031_ vssd1 vssd1 vccd1 vccd1 _1428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6671__158 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__inv_2
XFILLER_0_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2925_ clknet_0__2925_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2925_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5921_ _2386_ vssd1 vssd1 vccd1 vccd1 _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5852_ _3137_ _0407_ vssd1 vssd1 vccd1 vccd1 _2324_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5783_ _3113_ _3149_ vssd1 vssd1 vccd1 vccd1 _2255_ sky130_fd_sc_hd__nand2_1
X_4803_ _3056_ _1281_ _1283_ vssd1 vssd1 vccd1 vccd1 _0292_ sky130_fd_sc_hd__o21a_1
X_4734_ _3010_ _3356_ _3013_ _3360_ _1214_ vssd1 vssd1 vccd1 vccd1 _1215_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4665_ _0890_ _0561_ _1144_ _1145_ _1146_ vssd1 vssd1 vccd1 vccd1 _1147_ sky130_fd_sc_hd__o2111a_1
X_4596_ _3330_ _3345_ vssd1 vssd1 vccd1 vccd1 _1078_ sky130_fd_sc_hd__nand2_1
X_3616_ _2964_ _3064_ vssd1 vssd1 vccd1 vccd1 _3150_ sky130_fd_sc_hd__and2_1
X_6404_ _2745_ _2746_ vssd1 vssd1 vccd1 vccd1 _2747_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6335_ _2677_ _2656_ vssd1 vssd1 vccd1 vccd1 _2678_ sky130_fd_sc_hd__nand2_1
X_3547_ _3080_ _3060_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3081_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3478_ net2 _3022_ _3007_ vssd1 vssd1 vccd1 vccd1 _3023_ sky130_fd_sc_hd__mux2_1
X_6266_ _2621_ vssd1 vssd1 vccd1 vccd1 _0173_ sky130_fd_sc_hd__clkbuf_1
X_5217_ _3313_ _3010_ vssd1 vssd1 vccd1 vccd1 _1694_ sky130_fd_sc_hd__nand2_1
X_6197_ net13 _3310_ _2557_ vssd1 vssd1 vccd1 vccd1 _2576_ sky130_fd_sc_hd__mux2_1
X_5148_ _0467_ _0488_ _0475_ _0492_ _1625_ vssd1 vssd1 vccd1 vccd1 _1626_ sky130_fd_sc_hd__a221oi_1
X_5079_ _1548_ _1551_ _1554_ _1556_ vssd1 vssd1 vccd1 vccd1 _1557_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6608__100 clknet_1_1__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__inv_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6654__142 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__inv_2
XFILLER_0_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _3250_ _3272_ vssd1 vssd1 vccd1 vccd1 _0933_ sky130_fd_sc_hd__nand2_1
X_4381_ _0864_ vssd1 vssd1 vccd1 vccd1 _0865_ sky130_fd_sc_hd__inv_2
X_6741__66 clknet_1_1__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__inv_2
X_3401_ net18 vssd1 vssd1 vccd1 vccd1 _2955_ sky130_fd_sc_hd__inv_2
X_6120_ _2523_ vssd1 vssd1 vccd1 vccd1 _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _2474_ _2475_ vssd1 vssd1 vccd1 vccd1 _2476_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _0399_ _0451_ vssd1 vssd1 vccd1 vccd1 _1481_ sky130_fd_sc_hd__nand2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6884_ net82 _0287_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ sky130_fd_sc_hd__dfxtp_2
X_5904_ _2374_ vssd1 vssd1 vccd1 vccd1 _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5835_ _2266_ _2277_ _2290_ _2306_ vssd1 vssd1 vccd1 vccd1 _2307_ sky130_fd_sc_hd__and4_1
XFILLER_0_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5766_ _0562_ _0503_ vssd1 vssd1 vccd1 vccd1 _2239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4717_ _3327_ _3281_ _3341_ _3285_ _1197_ vssd1 vssd1 vccd1 vccd1 _1198_ sky130_fd_sc_hd__a221oi_1
X_5697_ _3304_ _3280_ _3353_ _3284_ _2169_ vssd1 vssd1 vccd1 vccd1 _2170_ sky130_fd_sc_hd__a221oi_1
X_4648_ _0513_ _0488_ _0515_ _0492_ _1129_ vssd1 vssd1 vccd1 vccd1 _1130_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4579_ _3246_ _3265_ vssd1 vssd1 vccd1 vccd1 _1061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6318_ _2660_ vssd1 vssd1 vccd1 vccd1 _2661_ sky130_fd_sc_hd__inv_2
X_6249_ _2989_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _2610_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3950_ _0435_ vssd1 vssd1 vccd1 vccd1 _0436_ sky130_fd_sc_hd__clkbuf_4
X_3881_ egd_top.BitStream_buffer.BS_buffer\[34\] vssd1 vssd1 vccd1 vccd1 _0367_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5620_ _0461_ _0431_ _0455_ _0435_ _2093_ vssd1 vssd1 vccd1 vccd1 _2094_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5551_ _3159_ _0653_ vssd1 vssd1 vccd1 vccd1 _2025_ sky130_fd_sc_hd__nand2_1
X_4502_ _0981_ _0414_ _0982_ _0983_ _0984_ vssd1 vssd1 vccd1 vccd1 _0985_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5482_ _1955_ _1956_ vssd1 vssd1 vccd1 vccd1 _1957_ sky130_fd_sc_hd__nor2_1
X_4433_ egd_top.BitStream_buffer.BS_buffer\[120\] vssd1 vssd1 vccd1 vccd1 _0916_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4364_ _0451_ vssd1 vssd1 vccd1 vccd1 _0848_ sky130_fd_sc_hd__inv_2
X_6103_ _2511_ vssd1 vssd1 vccd1 vccd1 _0220_ sky130_fd_sc_hd__clkbuf_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _0766_ _0770_ _0774_ _0778_ vssd1 vssd1 vccd1 vccd1 _0779_ sky130_fd_sc_hd__and4_1
X_6034_ net16 _0353_ _2451_ vssd1 vssd1 vccd1 vccd1 _2464_ sky130_fd_sc_hd__mux2_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ net65 _0270_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5818_ _2279_ _2284_ _2287_ _2289_ vssd1 vssd1 vccd1 vccd1 _2290_ sky130_fd_sc_hd__and4_1
X_6798_ net152 _0201_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[78\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5749_ _0347_ _0471_ _2219_ _2221_ vssd1 vssd1 vccd1 vccd1 _2222_ sky130_fd_sc_hd__o211a_1
X_6705__33 clknet_1_1__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__inv_2
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6720__47 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__inv_2
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4080_ _0565_ vssd1 vssd1 vccd1 vccd1 _0566_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _3365_ _3022_ vssd1 vssd1 vccd1 vccd1 _1461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3933_ _3061_ _0395_ vssd1 vssd1 vccd1 vccd1 _0419_ sky130_fd_sc_hd__and2_1
X_3864_ _0343_ _0345_ _0347_ _0349_ vssd1 vssd1 vccd1 vccd1 _0350_ sky130_fd_sc_hd__o22ai_1
X_5603_ _0370_ _0695_ vssd1 vssd1 vccd1 vccd1 _2077_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6583_ clknet_1_1__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2914_ sky130_fd_sc_hd__buf_1
X_3795_ _3098_ _3300_ vssd1 vssd1 vccd1 vccd1 _3329_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5534_ _2000_ _2004_ _2006_ _2008_ vssd1 vssd1 vccd1 vccd1 _2009_ sky130_fd_sc_hd__and4_1
X_5465_ _1938_ _1939_ vssd1 vssd1 vccd1 vccd1 _1940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4416_ _3056_ _0896_ _0899_ vssd1 vssd1 vccd1 vccd1 _0295_ sky130_fd_sc_hd__o21a_1
X_5396_ _1741_ _0506_ _1869_ _1870_ _1871_ vssd1 vssd1 vccd1 vccd1 _1872_ sky130_fd_sc_hd__o2111a_1
X_4347_ _0829_ _0830_ vssd1 vssd1 vccd1 vccd1 _0831_ sky130_fd_sc_hd__nand2_1
X_4278_ egd_top.BitStream_buffer.BitStream_buffer_output\[14\] _2997_ _2989_ vssd1
+ vssd1 vccd1 vccd1 _0763_ sky130_fd_sc_hd__o21a_1
X_6017_ _2452_ _2448_ vssd1 vssd1 vccd1 vccd1 _2453_ sky130_fd_sc_hd__and2_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3580_ _3113_ vssd1 vssd1 vccd1 vccd1 _3114_ sky130_fd_sc_hd__clkbuf_4
X_5250_ _3108_ _0408_ vssd1 vssd1 vccd1 vccd1 _1727_ sky130_fd_sc_hd__or2_1
X_4201_ _0347_ _0345_ _0685_ _0349_ vssd1 vssd1 vccd1 vccd1 _0686_ sky130_fd_sc_hd__o22ai_1
X_5181_ _3086_ _3111_ _1657_ vssd1 vssd1 vccd1 vccd1 _1658_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4132_ _3102_ _3101_ _3129_ _3106_ _0616_ vssd1 vssd1 vccd1 vccd1 _0617_ sky130_fd_sc_hd__a221oi_1
X_4063_ _0547_ _0548_ vssd1 vssd1 vccd1 vccd1 _0549_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4965_ egd_top.BitStream_buffer.BS_buffer\[100\] vssd1 vssd1 vccd1 vccd1 _1444_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3916_ _3126_ _0395_ vssd1 vssd1 vccd1 vccd1 _0402_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4896_ _1375_ vssd1 vssd1 vccd1 vccd1 _1376_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3847_ _3090_ _0325_ vssd1 vssd1 vccd1 vccd1 _0333_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6566_ _2879_ _2878_ vssd1 vssd1 vccd1 vccd1 _2899_ sky130_fd_sc_hd__or2_1
X_3778_ _3082_ _3300_ vssd1 vssd1 vccd1 vccd1 _3312_ sky130_fd_sc_hd__and2_1
X_5517_ _0530_ _0339_ vssd1 vssd1 vccd1 vccd1 _1992_ sky130_fd_sc_hd__nand2_1
X_6497_ _2830_ _2832_ _2710_ vssd1 vssd1 vccd1 vccd1 _2833_ sky130_fd_sc_hd__nand3_1
X_5448_ _3246_ _3286_ vssd1 vssd1 vccd1 vccd1 _1923_ sky130_fd_sc_hd__nand2_1
X_5379_ _0711_ _0440_ _1854_ vssd1 vssd1 vccd1 vccd1 _1855_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4750_ _0443_ _0379_ _0429_ _0383_ _1230_ vssd1 vssd1 vccd1 vccd1 _1231_ sky130_fd_sc_hd__a221oi_2
X_3701_ _3234_ vssd1 vssd1 vccd1 vccd1 _3235_ sky130_fd_sc_hd__buf_4
X_4681_ _3114_ _3134_ vssd1 vssd1 vccd1 vccd1 _1162_ sky130_fd_sc_hd__nand2_1
X_6420_ _2669_ _2700_ _1894_ vssd1 vssd1 vccd1 vccd1 _2762_ sky130_fd_sc_hd__o21ai_1
X_3632_ egd_top.BitStream_buffer.pc\[6\] egd_top.BitStream_buffer.pc\[4\] egd_top.BitStream_buffer.pc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _3166_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6351_ _2692_ _2693_ vssd1 vssd1 vccd1 vccd1 _2694_ sky130_fd_sc_hd__nand2_1
X_3563_ _3060_ _3096_ vssd1 vssd1 vccd1 vccd1 _3097_ sky130_fd_sc_hd__nand2_4
X_5302_ _0646_ _3068_ _3265_ _3075_ _1777_ vssd1 vssd1 vccd1 vccd1 _1778_ sky130_fd_sc_hd__a221oi_1
X_3494_ net13 _3034_ _3007_ vssd1 vssd1 vccd1 vccd1 _3035_ sky130_fd_sc_hd__mux2_1
X_6282_ net13 _0804_ _2613_ vssd1 vssd1 vccd1 vccd1 _2632_ sky130_fd_sc_hd__mux2_1
X_5233_ _0334_ _0429_ vssd1 vssd1 vccd1 vccd1 _1710_ sky130_fd_sc_hd__nand2_1
X_5164_ _1150_ _0570_ vssd1 vssd1 vccd1 vccd1 _1642_ sky130_fd_sc_hd__or2_1
X_4115_ _0558_ _0572_ _0586_ _0600_ vssd1 vssd1 vccd1 vccd1 _0601_ sky130_fd_sc_hd__and4_1
X_5095_ _1571_ _1572_ vssd1 vssd1 vccd1 vccd1 _1573_ sky130_fd_sc_hd__nand2_1
X_4046_ _0530_ _0531_ vssd1 vssd1 vccd1 vccd1 _0532_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5997_ _2438_ vssd1 vssd1 vccd1 vccd1 _0253_ sky130_fd_sc_hd__clkbuf_1
X_6747__72 clknet_1_0__leaf__2927_ vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__inv_2
X_4948_ _3053_ _3184_ _0607_ _3187_ _1426_ vssd1 vssd1 vccd1 vccd1 _1427_ sky130_fd_sc_hd__a221oi_1
X_4879_ _0848_ _0408_ vssd1 vssd1 vccd1 vccd1 _1359_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6549_ _2881_ _2710_ _2882_ vssd1 vssd1 vccd1 vccd1 _2883_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6690__19 clknet_1_1__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__inv_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6596__89 clknet_1_1__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__inv_2
XFILLER_0_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6755__3 clknet_1_0__leaf__2914_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__2924_ clknet_0__2924_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2924_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5920_ _2385_ _3042_ vssd1 vssd1 vccd1 vccd1 _2386_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5851_ _0402_ _3095_ vssd1 vssd1 vccd1 vccd1 _2323_ sky130_fd_sc_hd__nand2_1
X_5782_ _0653_ _3067_ _0804_ _3074_ _2253_ vssd1 vssd1 vccd1 vccd1 _2254_ sky130_fd_sc_hd__a221oi_1
X_4802_ _1282_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1283_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4733_ _3174_ _3363_ _1213_ vssd1 vssd1 vccd1 vccd1 _1214_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6403_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2746_ sky130_fd_sc_hd__nand2_1
X_4664_ _0596_ _0570_ vssd1 vssd1 vccd1 vccd1 _1146_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ _3326_ _3335_ vssd1 vssd1 vccd1 vccd1 _1077_ sky130_fd_sc_hd__nand2_1
X_3615_ egd_top.BitStream_buffer.BS_buffer\[79\] vssd1 vssd1 vccd1 vccd1 _3149_ sky130_fd_sc_hd__clkbuf_4
X_6631__121 clknet_1_1__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__inv_2
XFILLER_0_3_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6334_ _2676_ _1406_ vssd1 vssd1 vccd1 vccd1 _2677_ sky130_fd_sc_hd__nand2_1
X_3546_ _3079_ vssd1 vssd1 vccd1 vccd1 _3080_ sky130_fd_sc_hd__inv_2
X_6265_ _2620_ _2581_ vssd1 vssd1 vccd1 vccd1 _2621_ sky130_fd_sc_hd__and2_1
X_5216_ _3309_ _3013_ vssd1 vssd1 vccd1 vccd1 _1693_ sky130_fd_sc_hd__nand2_1
X_3477_ egd_top.BitStream_buffer.BS_buffer\[117\] vssd1 vssd1 vccd1 vccd1 _3022_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6196_ _2575_ vssd1 vssd1 vccd1 vccd1 _0191_ sky130_fd_sc_hd__clkbuf_1
X_5147_ _0862_ _0496_ _1624_ vssd1 vssd1 vccd1 vccd1 _1625_ sky130_fd_sc_hd__o21ai_1
X_5078_ _0548_ _3212_ egd_top.BitStream_buffer.BS_buffer\[7\] _3215_ _1555_ vssd1
+ vssd1 vccd1 vccd1 _1556_ sky130_fd_sc_hd__a221oi_1
X_4029_ egd_top.BitStream_buffer.BS_buffer\[21\] vssd1 vssd1 vccd1 vccd1 _0515_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6726__53 clknet_1_1__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__inv_2
XFILLER_0_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4380_ _0478_ _0535_ _0481_ _0531_ vssd1 vssd1 vccd1 vccd1 _0864_ sky130_fd_sc_hd__a22o_1
X_3400_ egd_top.BitStream_buffer.pc\[2\] egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1
+ vccd1 vccd1 _2954_ sky130_fd_sc_hd__nand2_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ _2932_ vssd1 vssd1 vccd1 vccd1 _2475_ sky130_fd_sc_hd__buf_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _1469_ _1473_ _1476_ _1479_ vssd1 vssd1 vccd1 vccd1 _1480_ sky130_fd_sc_hd__and4_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5903_ _3007_ _2372_ _2373_ vssd1 vssd1 vccd1 vccd1 _2374_ sky130_fd_sc_hd__and3_1
X_6883_ net81 _0286_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5834_ _2294_ _2298_ _2302_ _2305_ vssd1 vssd1 vccd1 vccd1 _2306_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5765_ _0494_ _0544_ _2235_ _2236_ _2237_ vssd1 vssd1 vccd1 vccd1 _2238_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4716_ _1069_ _3289_ _1196_ _3293_ vssd1 vssd1 vccd1 vccd1 _1197_ sky130_fd_sc_hd__o22ai_1
X_5696_ _0819_ _3288_ _0952_ _3292_ vssd1 vssd1 vccd1 vccd1 _2169_ sky130_fd_sc_hd__o22ai_1
X_4647_ _0734_ _0496_ _1128_ vssd1 vssd1 vccd1 vccd1 _1129_ sky130_fd_sc_hd__o21ai_1
X_4578_ _3278_ _3231_ _3282_ _3235_ _1059_ vssd1 vssd1 vccd1 vccd1 _1060_ sky130_fd_sc_hd__a221oi_1
X_6317_ egd_top.BitStream_buffer.BitStream_buffer_output\[6\] egd_top.BitStream_buffer.BitStream_buffer_output\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2660_ sky130_fd_sc_hd__nor2_1
X_3529_ egd_top.BitStream_buffer.pc\[5\] vssd1 vssd1 vccd1 vccd1 _3063_ sky130_fd_sc_hd__inv_2
X_6248_ _2960_ _2593_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[1\] sky130_fd_sc_hd__xor2_4
X_6179_ net4 _3327_ _2557_ vssd1 vssd1 vccd1 vccd1 _2564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6638__127 clknet_1_0__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__inv_2
XFILLER_0_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _0365_ vssd1 vssd1 vccd1 vccd1 _0366_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5550_ _3154_ _0804_ vssd1 vssd1 vccd1 vccd1 _2024_ sky130_fd_sc_hd__nand2_1
X_5481_ _0352_ _0443_ _0355_ _0429_ vssd1 vssd1 vccd1 vccd1 _1956_ sky130_fd_sc_hd__a22o_1
X_4501_ _0708_ _0426_ vssd1 vssd1 vccd1 vccd1 _0984_ sky130_fd_sc_hd__or2_1
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4432_ _0902_ _0906_ _0910_ _0914_ vssd1 vssd1 vccd1 vccd1 _0915_ sky130_fd_sc_hd__and4_1
X_4363_ _0406_ _0397_ _0844_ _0845_ _0846_ vssd1 vssd1 vccd1 vccd1 _0847_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6102_ _2510_ _2502_ vssd1 vssd1 vccd1 vccd1 _2511_ sky130_fd_sc_hd__and2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4294_ _3255_ _3148_ _3247_ _3152_ _0777_ vssd1 vssd1 vccd1 vccd1 _0778_ sky130_fd_sc_hd__a221oi_1
X_6033_ _2463_ vssd1 vssd1 vccd1 vccd1 _0242_ sky130_fd_sc_hd__clkbuf_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6866_ net64 _0269_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[10\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_91_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5817_ _3353_ _3280_ _3357_ _3284_ _2288_ vssd1 vssd1 vccd1 vccd1 _2289_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6797_ net151 _0200_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[79\]
+ sky130_fd_sc_hd__dfxtp_1
X_5748_ _2220_ vssd1 vssd1 vccd1 vccd1 _2221_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5679_ _0540_ _3183_ _0548_ _3186_ _2151_ vssd1 vssd1 vccd1 vccd1 _2152_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_40_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ _1456_ _3338_ _1457_ _1458_ _1459_ vssd1 vssd1 vccd1 vccd1 _1460_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3932_ _0416_ _0417_ vssd1 vssd1 vccd1 vccd1 _0418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3863_ _0348_ vssd1 vssd1 vccd1 vccd1 _0349_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5602_ _2074_ _2075_ vssd1 vssd1 vccd1 vccd1 _2076_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6582_ wb_clk_i vssd1 vssd1 vccd1 vccd1 _2913_ sky130_fd_sc_hd__buf_1
X_5533_ _0475_ _0589_ _0479_ _0592_ _2007_ vssd1 vssd1 vccd1 vccd1 _2008_ sky130_fd_sc_hd__a221oi_1
X_3794_ _3326_ _3327_ vssd1 vssd1 vccd1 vccd1 _3328_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5464_ _3330_ _3357_ vssd1 vssd1 vccd1 vccd1 _1939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5395_ _1497_ _0518_ vssd1 vssd1 vccd1 vccd1 _1871_ sky130_fd_sc_hd__or2_1
X_4415_ _0897_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _0899_ sky130_fd_sc_hd__a21oi_1
X_4346_ _0338_ _0323_ vssd1 vssd1 vccd1 vccd1 _0830_ sky130_fd_sc_hd__nand2_1
X_4277_ _0680_ _0760_ _0761_ vssd1 vssd1 vccd1 vccd1 _0762_ sky130_fd_sc_hd__nand3_1
X_6016_ net7 _0359_ _2451_ vssd1 vssd1 vccd1 vccd1 _2452_ sky130_fd_sc_hd__mux2_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6918_ net39 _0321_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6849_ net47 _0252_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[27\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6696__25 clknet_1_0__leaf__2923_ vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__inv_2
X_4200_ egd_top.BitStream_buffer.BS_buffer\[38\] vssd1 vssd1 vccd1 vccd1 _0685_ sky130_fd_sc_hd__inv_2
X_5180_ _3114_ _3057_ vssd1 vssd1 vccd1 vccd1 _1657_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4131_ _0614_ _3111_ _0615_ vssd1 vssd1 vccd1 vccd1 _0616_ sky130_fd_sc_hd__o21ai_1
X_4062_ egd_top.BitStream_buffer.BS_buffer\[6\] vssd1 vssd1 vccd1 vccd1 _0548_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4964_ _1441_ _1442_ vssd1 vssd1 vccd1 vccd1 _1443_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3915_ _0399_ _0400_ vssd1 vssd1 vccd1 vccd1 _0401_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4895_ _0478_ _0359_ _0481_ _0363_ vssd1 vssd1 vccd1 vccd1 _1375_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3846_ _0331_ vssd1 vssd1 vccd1 vccd1 _0332_ sky130_fd_sc_hd__buf_6
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3777_ _3309_ _3310_ vssd1 vssd1 vccd1 vccd1 _3311_ sky130_fd_sc_hd__nand2_1
X_6565_ _2848_ _2884_ _2869_ vssd1 vssd1 vccd1 vccd1 _2898_ sky130_fd_sc_hd__nand3_1
X_5516_ _0367_ _0506_ _1988_ _1989_ _1990_ vssd1 vssd1 vccd1 vccd1 _1991_ sky130_fd_sc_hd__o2111a_1
X_6496_ _2831_ _2828_ vssd1 vssd1 vccd1 vccd1 _2832_ sky130_fd_sc_hd__nand2_1
X_5447_ _3347_ _3231_ _3345_ _3235_ _1921_ vssd1 vssd1 vccd1 vccd1 _1922_ sky130_fd_sc_hd__a221oi_1
X_5378_ _0442_ _0411_ vssd1 vssd1 vccd1 vccd1 _1854_ sky130_fd_sc_hd__nand2_1
X_4329_ _0811_ _0812_ vssd1 vssd1 vccd1 vccd1 _0813_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3700_ _3233_ vssd1 vssd1 vccd1 vccd1 _3234_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4680_ _3149_ _3068_ _3255_ _3075_ _1160_ vssd1 vssd1 vccd1 vccd1 _1161_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3631_ _3094_ _3118_ _3143_ _3164_ vssd1 vssd1 vccd1 vccd1 _3165_ sky130_fd_sc_hd__and4_1
XFILLER_0_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6350_ _2681_ _2686_ vssd1 vssd1 vccd1 vccd1 _2693_ sky130_fd_sc_hd__nand2_2
X_3562_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3096_ sky130_fd_sc_hd__inv_2
X_5301_ _1654_ _3084_ _1776_ _3092_ vssd1 vssd1 vccd1 vccd1 _1777_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3493_ egd_top.BitStream_buffer.BS_buffer\[121\] vssd1 vssd1 vccd1 vccd1 _3034_ sky130_fd_sc_hd__clkbuf_4
X_6281_ _2631_ vssd1 vssd1 vccd1 vccd1 _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5232_ _1668_ _1679_ _1692_ _1708_ vssd1 vssd1 vccd1 vccd1 _1709_ sky130_fd_sc_hd__and4_1
X_5163_ _0566_ egd_top.BitStream_buffer.BS_buffer\[16\] vssd1 vssd1 vccd1 vccd1 _1641_
+ sky130_fd_sc_hd__nand2_1
X_4114_ egd_top.BitStream_buffer.BS_buffer\[14\] _0589_ egd_top.BitStream_buffer.BS_buffer\[15\]
+ _0592_ _0599_ vssd1 vssd1 vccd1 vccd1 _0600_ sky130_fd_sc_hd__a221oi_1
X_5094_ _3313_ _2998_ vssd1 vssd1 vccd1 vccd1 _1572_ sky130_fd_sc_hd__nand2_1
X_4045_ egd_top.BitStream_buffer.BS_buffer\[29\] vssd1 vssd1 vccd1 vccd1 _0531_ sky130_fd_sc_hd__clkbuf_4
X_5996_ _2437_ _2423_ vssd1 vssd1 vccd1 vccd1 _2438_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4947_ _0574_ _3190_ _1425_ vssd1 vssd1 vccd1 vccd1 _1426_ sky130_fd_sc_hd__o21ai_1
X_4878_ _0403_ _0421_ vssd1 vssd1 vccd1 vccd1 _1358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _3362_ vssd1 vssd1 vccd1 vccd1 _3363_ sky130_fd_sc_hd__clkbuf_4
X_6548_ _2831_ _2877_ _2879_ vssd1 vssd1 vccd1 vccd1 _2882_ sky130_fd_sc_hd__nand3_1
X_6479_ _2817_ _2818_ _2819_ vssd1 vssd1 vccd1 vccd1 _2820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2923_ clknet_0__2923_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2923_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5850_ _0398_ _3129_ vssd1 vssd1 vccd1 vccd1 _2322_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5781_ _0651_ _3083_ _0802_ _3091_ vssd1 vssd1 vccd1 vccd1 _2253_ sky130_fd_sc_hd__o22ai_1
X_4801_ egd_top.BitStream_buffer.BitStream_buffer_output\[10\] vssd1 vssd1 vccd1 vccd1
+ _1282_ sky130_fd_sc_hd__inv_2
X_4732_ _3365_ _3016_ vssd1 vssd1 vccd1 vccd1 _1213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _0566_ egd_top.BitStream_buffer.BS_buffer\[12\] vssd1 vssd1 vccd1 vccd1 _1145_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3614_ _3147_ vssd1 vssd1 vccd1 vccd1 _3148_ sky130_fd_sc_hd__buf_4
X_6402_ _2744_ vssd1 vssd1 vccd1 vccd1 _2745_ sky130_fd_sc_hd__inv_2
X_4594_ _0674_ _3303_ _0675_ _3307_ _1075_ vssd1 vssd1 vccd1 vccd1 _1076_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6333_ _2675_ _1530_ vssd1 vssd1 vccd1 vccd1 _2676_ sky130_fd_sc_hd__nand2_1
X_3545_ _2961_ _3078_ vssd1 vssd1 vccd1 vccd1 _3079_ sky130_fd_sc_hd__nand2_2
X_3476_ _3021_ vssd1 vssd1 vccd1 vccd1 _0309_ sky130_fd_sc_hd__clkbuf_1
X_6264_ net4 _3251_ _2613_ vssd1 vssd1 vccd1 vccd1 _2620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ _1681_ _1686_ _1689_ _1691_ vssd1 vssd1 vccd1 vccd1 _1692_ sky130_fd_sc_hd__and4_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6195_ _2574_ _2554_ vssd1 vssd1 vccd1 vccd1 _2575_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5146_ _0498_ _0482_ vssd1 vssd1 vccd1 vccd1 _1624_ sky130_fd_sc_hd__nand2_1
X_5077_ _0753_ _3218_ _0541_ _3221_ vssd1 vssd1 vccd1 vccd1 _1555_ sky130_fd_sc_hd__o22ai_1
X_4028_ _0512_ _0513_ vssd1 vssd1 vccd1 vccd1 _0514_ sky130_fd_sc_hd__nand2_1
X_5979_ _2426_ vssd1 vssd1 vccd1 vccd1 _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6615__106 clknet_1_0__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__inv_2
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _0433_ _0379_ _0404_ _0383_ _1478_ vssd1 vssd1 vccd1 vccd1 _1479_ sky130_fd_sc_hd__a221oi_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6882_ net80 _0285_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_5902_ _3004_ _2978_ vssd1 vssd1 vccd1 vccd1 _2373_ sky130_fd_sc_hd__nand2_1
X_5833_ _3037_ _3355_ _3040_ _3359_ _2304_ vssd1 vssd1 vccd1 vccd1 _2305_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_29_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5764_ _0867_ _0555_ vssd1 vssd1 vccd1 vccd1 _2237_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4715_ _3331_ vssd1 vssd1 vccd1 vccd1 _1196_ sky130_fd_sc_hd__inv_2
X_5695_ _2166_ _2167_ vssd1 vssd1 vccd1 vccd1 _2168_ sky130_fd_sc_hd__nor2_1
X_4646_ _0498_ _0503_ vssd1 vssd1 vccd1 vccd1 _1128_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4577_ _3287_ _3238_ _3291_ _3241_ vssd1 vssd1 vccd1 vccd1 _1059_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6316_ _2652_ _2658_ vssd1 vssd1 vccd1 vccd1 _2659_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ egd_top.BitStream_buffer.pc\[4\] vssd1 vssd1 vccd1 vccd1 _3062_ sky130_fd_sc_hd__inv_2
X_3459_ _3008_ _2933_ vssd1 vssd1 vccd1 vccd1 _3009_ sky130_fd_sc_hd__and2_1
X_6247_ _2609_ vssd1 vssd1 vccd1 vccd1 _0179_ sky130_fd_sc_hd__inv_2
X_6178_ _2563_ vssd1 vssd1 vccd1 vccd1 _0197_ sky130_fd_sc_hd__clkbuf_1
X_5129_ _0416_ _3107_ vssd1 vssd1 vccd1 vccd1 _1607_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480_ _0384_ _0345_ _0438_ _0349_ vssd1 vssd1 vccd1 vccd1 _1955_ sky130_fd_sc_hd__o22ai_1
X_4500_ _0420_ _0451_ vssd1 vssd1 vccd1 vccd1 _0983_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431_ _3247_ _3148_ _3259_ _3152_ _0913_ vssd1 vssd1 vccd1 vccd1 _0914_ sky130_fd_sc_hd__a221oi_1
XANTENNA_1 _1217_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4362_ _0424_ _0408_ vssd1 vssd1 vccd1 vccd1 _0846_ sky130_fd_sc_hd__or2_1
X_6101_ net11 _0411_ _2486_ vssd1 vssd1 vccd1 vccd1 _2510_ sky130_fd_sc_hd__mux2_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _0775_ _0776_ vssd1 vssd1 vccd1 vccd1 _0777_ sky130_fd_sc_hd__nand2_1
X_6032_ _2462_ _2448_ vssd1 vssd1 vccd1 vccd1 _2463_ sky130_fd_sc_hd__and2_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6865_ net63 _0268_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[11\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6796_ net150 _0199_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[96\]
+ sky130_fd_sc_hd__dfxtp_1
X_5816_ _0952_ _3288_ _1081_ _3292_ vssd1 vssd1 vccd1 vccd1 _2288_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5747_ _0477_ egd_top.BitStream_buffer.BS_buffer\[39\] _0480_ _0339_ vssd1 vssd1
+ vccd1 vccd1 _2220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5678_ _0745_ _3189_ _2150_ vssd1 vssd1 vccd1 vccd1 _2151_ sky130_fd_sc_hd__o21ai_1
X_4629_ _0420_ _0461_ vssd1 vssd1 vccd1 vccd1 _1111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4980_ _1208_ _3350_ vssd1 vssd1 vccd1 vccd1 _1459_ sky130_fd_sc_hd__or2_1
X_3931_ egd_top.BitStream_buffer.BS_buffer\[56\] vssd1 vssd1 vccd1 vccd1 _0417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3862_ _3139_ _0325_ vssd1 vssd1 vccd1 vccd1 _0348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5601_ _0351_ _0429_ _0354_ _0433_ vssd1 vssd1 vccd1 vccd1 _2075_ sky130_fd_sc_hd__a22o_1
X_6581_ _2756_ _2907_ _2912_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__a21bo_1
X_5532_ _0504_ _0595_ _0468_ _0598_ vssd1 vssd1 vccd1 vccd1 _2007_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_5_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3793_ egd_top.BitStream_buffer.BS_buffer\[99\] vssd1 vssd1 vccd1 vccd1 _3327_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5463_ _3326_ _0674_ vssd1 vssd1 vccd1 vccd1 _1938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5394_ _0512_ _0521_ vssd1 vssd1 vccd1 vccd1 _1870_ sky130_fd_sc_hd__nand2_1
X_4414_ _2996_ vssd1 vssd1 vccd1 vccd1 _0898_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4345_ _0334_ _0329_ vssd1 vssd1 vccd1 vccd1 _0829_ sky130_fd_sc_hd__nand2_1
X_6667__154 clknet_1_1__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__inv_2
X_4276_ _0606_ _0577_ vssd1 vssd1 vccd1 vccd1 _0761_ sky130_fd_sc_hd__nand2_1
X_6015_ _2450_ vssd1 vssd1 vccd1 vccd1 _2451_ sky130_fd_sc_hd__buf_4
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6917_ net38 _0320_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__dfxtp_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6848_ net46 _0251_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6779_ net133 _0182_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4130_ _3114_ _3095_ vssd1 vssd1 vccd1 vccd1 _0615_ sky130_fd_sc_hd__nand2_1
X_4061_ _0546_ vssd1 vssd1 vccd1 vccd1 _0547_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4963_ _3271_ _3290_ _3274_ _3278_ vssd1 vssd1 vccd1 vccd1 _1442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3914_ egd_top.BitStream_buffer.BS_buffer\[54\] vssd1 vssd1 vccd1 vccd1 _0400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4894_ _0474_ _0525_ vssd1 vssd1 vccd1 vccd1 _1374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3845_ _0330_ vssd1 vssd1 vccd1 vccd1 _0331_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3776_ egd_top.BitStream_buffer.BS_buffer\[105\] vssd1 vssd1 vccd1 vccd1 _3310_ sky130_fd_sc_hd__clkbuf_4
X_6564_ _2896_ _2897_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__nand2_1
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5515_ _1619_ _0518_ vssd1 vssd1 vccd1 vccd1 _1990_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6495_ _2761_ _2826_ vssd1 vssd1 vccd1 vccd1 _2831_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5446_ _1320_ _3238_ _1444_ _3241_ vssd1 vssd1 vccd1 vccd1 _1921_ sky130_fd_sc_hd__o22ai_1
X_5377_ _3137_ _0414_ _1850_ _1851_ _1852_ vssd1 vssd1 vccd1 vccd1 _1853_ sky130_fd_sc_hd__o2111a_1
X_4328_ _3313_ _3297_ vssd1 vssd1 vccd1 vccd1 _0812_ sky130_fd_sc_hd__nand2_1
X_4259_ _0551_ _0540_ vssd1 vssd1 vccd1 vccd1 _0744_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _3144_ _3148_ _3149_ _3152_ _3163_ vssd1 vssd1 vccd1 vccd1 _3164_ sky130_fd_sc_hd__a221oi_1
X_3561_ egd_top.BitStream_buffer.BS_buffer\[66\] vssd1 vssd1 vccd1 vccd1 _3095_ sky130_fd_sc_hd__clkbuf_4
X_5300_ egd_top.BitStream_buffer.BS_buffer\[83\] vssd1 vssd1 vccd1 vccd1 _1776_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3492_ _3033_ vssd1 vssd1 vccd1 vccd1 _0305_ sky130_fd_sc_hd__clkbuf_1
X_6280_ _2630_ _2372_ vssd1 vssd1 vccd1 vccd1 _2631_ sky130_fd_sc_hd__and2_1
X_5231_ _1696_ _1700_ _1704_ _1707_ vssd1 vssd1 vccd1 vccd1 _1708_ sky130_fd_sc_hd__and4_1
X_5162_ _0563_ _0493_ vssd1 vssd1 vccd1 vccd1 _1640_ sky130_fd_sc_hd__nand2_1
X_5093_ _3309_ _3010_ vssd1 vssd1 vccd1 vccd1 _1571_ sky130_fd_sc_hd__nand2_1
X_4113_ _0593_ _0595_ _0596_ _0598_ vssd1 vssd1 vccd1 vccd1 _0599_ sky130_fd_sc_hd__o22ai_1
X_4044_ _0529_ vssd1 vssd1 vccd1 vccd1 _0530_ sky130_fd_sc_hd__clkbuf_4
X_5995_ net12 _0479_ _2415_ vssd1 vssd1 vccd1 vccd1 _2437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4946_ _3192_ _0577_ vssd1 vssd1 vccd1 vccd1 _1425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _0399_ _0447_ vssd1 vssd1 vccd1 vccd1 _1357_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3828_ _2964_ _3300_ vssd1 vssd1 vccd1 vccd1 _3362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6547_ _2878_ _2880_ vssd1 vssd1 vccd1 vccd1 _2881_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3759_ _3292_ vssd1 vssd1 vccd1 vccd1 _3293_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6478_ net20 net21 vssd1 vssd1 vccd1 vccd1 _2819_ sky130_fd_sc_hd__nand2_1
X_5429_ _1654_ _3124_ _1901_ _1902_ _1903_ vssd1 vssd1 vccd1 vccd1 _1904_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2922_ clknet_0__2922_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2922_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4800_ _1217_ _1279_ _1280_ vssd1 vssd1 vccd1 vccd1 _1281_ sky130_fd_sc_hd__nand3_1
X_5780_ _0898_ _2250_ _2252_ vssd1 vssd1 vccd1 vccd1 _0284_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4731_ _1208_ _3338_ _1209_ _1210_ _1211_ vssd1 vssd1 vccd1 vccd1 _1212_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4662_ _0563_ egd_top.BitStream_buffer.BS_buffer\[14\] vssd1 vssd1 vccd1 vccd1 _1144_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3613_ _3146_ vssd1 vssd1 vccd1 vccd1 _3147_ sky130_fd_sc_hd__clkbuf_2
X_6401_ egd_top.BitStream_buffer.BitStream_buffer_output\[8\] egd_top.BitStream_buffer.BitStream_buffer_output\[7\]
+ vssd1 vssd1 vccd1 vccd1 _2744_ sky130_fd_sc_hd__nor2_1
X_4593_ _1073_ _1074_ vssd1 vssd1 vccd1 vccd1 _1075_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6332_ _2674_ _1652_ vssd1 vssd1 vccd1 vccd1 _2675_ sky130_fd_sc_hd__nand2_1
X_3544_ egd_top.BitStream_buffer.pc\[1\] vssd1 vssd1 vccd1 vccd1 _3078_ sky130_fd_sc_hd__inv_2
X_3475_ _3020_ _2933_ vssd1 vssd1 vccd1 vccd1 _3021_ sky130_fd_sc_hd__and2_1
X_6263_ _2619_ vssd1 vssd1 vccd1 vccd1 _0174_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5214_ _3335_ _3281_ _3314_ _3285_ _1690_ vssd1 vssd1 vccd1 vccd1 _1691_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_86_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6194_ net14 _3314_ _2557_ vssd1 vssd1 vccd1 vccd1 _2574_ sky130_fd_sc_hd__mux2_1
X_5145_ _1619_ _0472_ _1620_ _1622_ vssd1 vssd1 vccd1 vccd1 _1623_ sky130_fd_sc_hd__o211a_1
X_6680__10 clknet_1_1__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__inv_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5076_ _3037_ _3198_ _3040_ _3201_ _1553_ vssd1 vssd1 vccd1 vccd1 _1554_ sky130_fd_sc_hd__a221oi_1
X_4027_ egd_top.BitStream_buffer.BS_buffer\[20\] vssd1 vssd1 vccd1 vccd1 _0513_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5978_ _2425_ _2423_ vssd1 vssd1 vccd1 vccd1 _2426_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4929_ egd_top.BitStream_buffer.BS_buffer\[80\] vssd1 vssd1 vccd1 vccd1 _1408_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6661__149 clknet_1_1__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__inv_2
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5901_ net19 vssd1 vssd1 vccd1 vccd1 _2372_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6881_ net79 _0284_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5832_ _3219_ _3362_ _2303_ vssd1 vssd1 vccd1 vccd1 _2304_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5763_ _0550_ _0489_ vssd1 vssd1 vccd1 vccd1 _2236_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4714_ _1193_ _1194_ vssd1 vssd1 vccd1 vccd1 _1195_ sky130_fd_sc_hd__nor2_1
X_6717__44 clknet_1_0__leaf__2925_ vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__inv_2
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5694_ _3270_ _3327_ _3273_ _3341_ vssd1 vssd1 vccd1 vccd1 _2167_ sky130_fd_sc_hd__a22o_1
X_4645_ _1123_ _0472_ _1124_ _1126_ vssd1 vssd1 vccd1 vccd1 _1127_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4576_ _1049_ _1052_ _1055_ _1057_ vssd1 vssd1 vccd1 vccd1 _1058_ sky130_fd_sc_hd__and4_1
X_6732__58 clknet_1_1__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__inv_2
X_6315_ _2657_ vssd1 vssd1 vccd1 vccd1 _2658_ sky130_fd_sc_hd__inv_2
X_3527_ _3059_ _3060_ egd_top.BitStream_buffer.pc\[3\] vssd1 vssd1 vccd1 vccd1 _3061_
+ sky130_fd_sc_hd__and3_4
X_3458_ net7 _2998_ _3007_ vssd1 vssd1 vccd1 vccd1 _3008_ sky130_fd_sc_hd__mux2_1
X_6246_ _2989_ egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _2609_ sky130_fd_sc_hd__nand2_1
X_3389_ _2944_ vssd1 vssd1 vccd1 vccd1 _0319_ sky130_fd_sc_hd__clkbuf_1
X_6177_ _2562_ _2554_ vssd1 vssd1 vccd1 vccd1 _2563_ sky130_fd_sc_hd__and2_1
X_5128_ _0848_ _0397_ _1603_ _1604_ _1605_ vssd1 vssd1 vccd1 vccd1 _1606_ sky130_fd_sc_hd__o2111a_1
X_5059_ _3057_ _3101_ _3069_ _3106_ _1536_ vssd1 vssd1 vccd1 vccd1 _1537_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4430_ _0911_ _0912_ vssd1 vssd1 vccd1 vccd1 _0913_ sky130_fd_sc_hd__nand2_1
XANTENNA_2 _1635_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6100_ _2509_ vssd1 vssd1 vccd1 vccd1 _0221_ sky130_fd_sc_hd__clkbuf_1
X_4361_ _0403_ _0400_ vssd1 vssd1 vccd1 vccd1 _0845_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _3160_ _3144_ vssd1 vssd1 vccd1 vccd1 _0776_ sky130_fd_sc_hd__nand2_1
X_6031_ net2 _0346_ _2451_ vssd1 vssd1 vccd1 vccd1 _2462_ sky130_fd_sc_hd__mux2_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6864_ net62 _0267_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[12\]
+ sky130_fd_sc_hd__dfxtp_4
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5815_ _2285_ _2286_ vssd1 vssd1 vccd1 vccd1 _2287_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6795_ net149 _0198_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[97\]
+ sky130_fd_sc_hd__dfxtp_1
X_5746_ _0473_ _0353_ vssd1 vssd1 vccd1 vccd1 _2219_ sky130_fd_sc_hd__nand2_1
X_5677_ _3191_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _2150_
+ sky130_fd_sc_hd__nand2_1
X_4628_ _0416_ _0447_ vssd1 vssd1 vccd1 vccd1 _1110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4559_ _0764_ _3124_ _1038_ _1039_ _1040_ vssd1 vssd1 vccd1 vccd1 _1041_ sky130_fd_sc_hd__o2111a_1
X_6229_ _2600_ egd_top.BitStream_buffer.pc_previous\[4\] egd_top.BitStream_buffer.pc_previous\[5\]
+ vssd1 vssd1 vccd1 vccd1 _2601_ sky130_fd_sc_hd__and3_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6644__133 clknet_1_1__leaf__2919_ vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__inv_2
XFILLER_0_86_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6711__39 clknet_1_0__leaf__2924_ vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__inv_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3930_ _0415_ vssd1 vssd1 vccd1 vccd1 _0416_ sky130_fd_sc_hd__buf_4
X_3861_ _0346_ vssd1 vssd1 vccd1 vccd1 _0347_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5600_ _0438_ _0344_ _0714_ _0348_ vssd1 vssd1 vccd1 vccd1 _2074_ sky130_fd_sc_hd__o22ai_1
X_6580_ net18 _2650_ _2956_ _2900_ vssd1 vssd1 vccd1 vccd1 _2912_ sky130_fd_sc_hd__a211o_1
X_3792_ _3325_ vssd1 vssd1 vccd1 vccd1 _3326_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5531_ _0596_ _0576_ _0593_ _0580_ _2005_ vssd1 vssd1 vccd1 vccd1 _2006_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5462_ _3022_ _3303_ _3025_ _3307_ _1936_ vssd1 vssd1 vccd1 vccd1 _1937_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5393_ _0508_ _0359_ vssd1 vssd1 vccd1 vccd1 _1869_ sky130_fd_sc_hd__nand2_1
X_4413_ egd_top.BitStream_buffer.BitStream_buffer_output\[13\] vssd1 vssd1 vccd1 vccd1
+ _0897_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4344_ _0779_ _0793_ _0810_ _0827_ vssd1 vssd1 vccd1 vccd1 _0828_ sky130_fd_sc_hd__and4_1
X_4275_ _0722_ _0741_ _0759_ vssd1 vssd1 vccd1 vccd1 _0760_ sky130_fd_sc_hd__and3_1
X_6014_ net200 _2971_ net196 _3002_ vssd1 vssd1 vccd1 vccd1 _2450_ sky130_fd_sc_hd__or4b_4
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ net37 _0319_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__dfxtp_2
X_6847_ net45 _0250_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[29\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6778_ net132 _0181_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[4\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _2192_ _2195_ _2198_ _2201_ vssd1 vssd1 vccd1 vccd1 _2202_ sky130_fd_sc_hd__and4_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _3131_ _0543_ vssd1 vssd1 vccd1 vccd1 _0546_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4962_ _0794_ _3264_ _3287_ _3268_ vssd1 vssd1 vccd1 vccd1 _1441_ sky130_fd_sc_hd__o22ai_1
X_4893_ egd_top.BitStream_buffer.BS_buffer\[30\] vssd1 vssd1 vccd1 vccd1 _1373_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6701_ clknet_1_0__leaf__2913_ vssd1 vssd1 vccd1 vccd1 _2924_ sky130_fd_sc_hd__buf_1
X_3913_ _0398_ vssd1 vssd1 vccd1 vccd1 _0399_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3844_ _3072_ _0325_ vssd1 vssd1 vccd1 vccd1 _0330_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6563_ _2866_ _2852_ vssd1 vssd1 vccd1 vccd1 _2897_ sky130_fd_sc_hd__nand2_1
X_3775_ _3308_ vssd1 vssd1 vccd1 vccd1 _3309_ sky130_fd_sc_hd__buf_4
X_5514_ _0512_ _0525_ vssd1 vssd1 vccd1 vccd1 _1989_ sky130_fd_sc_hd__nand2_1
X_6494_ _2761_ _2826_ _2829_ vssd1 vssd1 vccd1 vccd1 _2830_ sky130_fd_sc_hd__o21ai_1
X_5445_ _1911_ _1914_ _1917_ _1919_ vssd1 vssd1 vccd1 vccd1 _1920_ sky130_fd_sc_hd__and4_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5376_ _0903_ _0426_ vssd1 vssd1 vccd1 vccd1 _1852_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4327_ _3309_ _3304_ vssd1 vssd1 vccd1 vccd1 _0811_ sky130_fd_sc_hd__nand2_1
X_4258_ _0547_ egd_top.BitStream_buffer.BS_buffer\[7\] vssd1 vssd1 vccd1 vccd1 _0743_
+ sky130_fd_sc_hd__nand2_1
X_4189_ egd_top.BitStream_buffer.BS_buffer\[110\] vssd1 vssd1 vccd1 vccd1 _0674_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3560_ _3057_ _3068_ _3069_ _3075_ _3093_ vssd1 vssd1 vccd1 vccd1 _3094_ sky130_fd_sc_hd__a221oi_1
X_3491_ _3032_ _2933_ vssd1 vssd1 vccd1 vccd1 _3033_ sky130_fd_sc_hd__and2_1
X_5230_ _3022_ _3356_ _3025_ _3360_ _1706_ vssd1 vssd1 vccd1 vccd1 _1707_ sky130_fd_sc_hd__a221oi_1
X_5161_ _0596_ _0545_ _1636_ _1637_ _1638_ vssd1 vssd1 vccd1 vccd1 _1639_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4112_ _0597_ vssd1 vssd1 vccd1 vccd1 _0598_ sky130_fd_sc_hd__clkbuf_4
X_5092_ _1559_ _1564_ _1567_ _1569_ vssd1 vssd1 vccd1 vccd1 _1570_ sky130_fd_sc_hd__and4_1
X_4043_ _3153_ _0470_ vssd1 vssd1 vccd1 vccd1 _0529_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5994_ _2436_ vssd1 vssd1 vccd1 vccd1 _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4945_ _3047_ _3170_ _3050_ _3173_ _1423_ vssd1 vssd1 vccd1 vccd1 _1424_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_86_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4876_ _1345_ _1349_ _1352_ _1355_ vssd1 vssd1 vccd1 vccd1 _1356_ sky130_fd_sc_hd__and4_1
X_6601__93 clknet_1_1__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__inv_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3827_ egd_top.BitStream_buffer.BS_buffer\[111\] vssd1 vssd1 vccd1 vccd1 _3361_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6546_ _2879_ vssd1 vssd1 vccd1 vccd1 _2880_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3758_ _3153_ _3228_ vssd1 vssd1 vccd1 vccd1 _3292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6477_ _2760_ _2786_ vssd1 vssd1 vccd1 vccd1 _2818_ sky130_fd_sc_hd__or2_1
X_3689_ _3050_ _3212_ _3053_ _3215_ _3222_ vssd1 vssd1 vccd1 vccd1 _3223_ sky130_fd_sc_hd__a221oi_1
X_5428_ _1408_ _3141_ vssd1 vssd1 vccd1 vccd1 _1903_ sky130_fd_sc_hd__or2_1
X_5359_ _0404_ _0328_ _0703_ _0332_ _1834_ vssd1 vssd1 vccd1 vccd1 _1835_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6738__64 clknet_1_0__leaf__2926_ vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__inv_2
XFILLER_0_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2921_ clknet_0__2921_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2921_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4730_ _0952_ _3350_ vssd1 vssd1 vccd1 vccd1 _1211_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4661_ _0568_ _0545_ _1140_ _1141_ _1142_ vssd1 vssd1 vccd1 vccd1 _1143_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ _3145_ _3064_ vssd1 vssd1 vccd1 vccd1 _3146_ sky130_fd_sc_hd__and2_1
X_6400_ _2696_ _2693_ vssd1 vssd1 vccd1 vccd1 _2743_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4592_ _3313_ _3353_ vssd1 vssd1 vccd1 vccd1 _1074_ sky130_fd_sc_hd__nand2_1
X_6331_ _2673_ _1774_ vssd1 vssd1 vccd1 vccd1 _2674_ sky130_fd_sc_hd__nand2_1
X_3543_ _3076_ vssd1 vssd1 vccd1 vccd1 _3077_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3474_ net3 _3019_ _3007_ vssd1 vssd1 vccd1 vccd1 _3020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6262_ _2618_ _2581_ vssd1 vssd1 vccd1 vccd1 _2619_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6193_ _2573_ vssd1 vssd1 vccd1 vccd1 _0192_ sky130_fd_sc_hd__clkbuf_1
X_5213_ _3348_ _3289_ _0671_ _3293_ vssd1 vssd1 vccd1 vccd1 _1690_ sky130_fd_sc_hd__o22ai_1
X_5144_ _1621_ vssd1 vssd1 vccd1 vccd1 _1622_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _0916_ _3204_ _1552_ vssd1 vssd1 vccd1 vccd1 _1553_ sky130_fd_sc_hd__o21ai_1
X_4026_ _0511_ vssd1 vssd1 vccd1 vccd1 _0512_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5977_ net3 _0513_ _2415_ vssd1 vssd1 vccd1 vccd1 _2425_ sky130_fd_sc_hd__mux2_1
X_4928_ _3056_ _1405_ _1407_ vssd1 vssd1 vccd1 vccd1 _0291_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4859_ _3013_ _3356_ _3016_ _3360_ _1338_ vssd1 vssd1 vccd1 vccd1 _1339_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6529_ _2737_ _2806_ vssd1 vssd1 vccd1 vccd1 _2864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5900_ _0898_ _2369_ _2371_ vssd1 vssd1 vccd1 vccd1 _0283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6880_ net78 _0283_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BitStream_buffer_output\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5831_ _3364_ _3044_ vssd1 vssd1 vccd1 vccd1 _2303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5762_ _0546_ _0499_ vssd1 vssd1 vccd1 vccd1 _2235_ sky130_fd_sc_hd__nand2_1
X_4713_ _3271_ _3232_ _3274_ _3286_ vssd1 vssd1 vccd1 vccd1 _1194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5693_ _1069_ _3263_ _1196_ _3267_ vssd1 vssd1 vccd1 vccd1 _2166_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_56_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4644_ _1125_ vssd1 vssd1 vccd1 vccd1 _1126_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4575_ _0573_ _3212_ _0581_ _3215_ _1056_ vssd1 vssd1 vccd1 vccd1 _1057_ sky130_fd_sc_hd__a221oi_1
X_6314_ _2656_ _1406_ _1530_ vssd1 vssd1 vccd1 vccd1 _2657_ sky130_fd_sc_hd__and3_1
X_3526_ egd_top.BitStream_buffer.pc\[2\] vssd1 vssd1 vccd1 vccd1 _3060_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6245_ _2608_ _2594_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc\[2\] sky130_fd_sc_hd__xnor2_4
X_3457_ _3006_ vssd1 vssd1 vccd1 vccd1 _3007_ sky130_fd_sc_hd__buf_4
X_6176_ net5 _3331_ _2557_ vssd1 vssd1 vccd1 vccd1 _2562_ sky130_fd_sc_hd__mux2_1
X_3388_ net32 _2942_ _2943_ vssd1 vssd1 vccd1 vccd1 _2944_ sky130_fd_sc_hd__o21ba_1
X_5127_ _0456_ _0408_ vssd1 vssd1 vccd1 vccd1 _1605_ sky130_fd_sc_hd__or2_1
X_5058_ _3077_ _3111_ _1535_ vssd1 vssd1 vccd1 vccd1 _1536_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4009_ _3098_ _0470_ vssd1 vssd1 vccd1 vccd1 _0495_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6621__112 clknet_1_1__leaf__2917_ vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__inv_2
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_3 _1692_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _0399_ _0417_ vssd1 vssd1 vccd1 vccd1 _0844_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _3155_ _3149_ vssd1 vssd1 vccd1 vccd1 _0775_ sky130_fd_sc_hd__nand2_1
X_6030_ _2461_ vssd1 vssd1 vccd1 vccd1 _0243_ sky130_fd_sc_hd__clkbuf_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6863_ net61 _0266_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_5814_ _3270_ _3341_ _3273_ _3347_ vssd1 vssd1 vccd1 vccd1 _2286_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6794_ net148 _0197_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[98\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5745_ _2202_ _2217_ vssd1 vssd1 vccd1 vccd1 _2218_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5676_ _0581_ _3169_ _0552_ _3172_ _2148_ vssd1 vssd1 vccd1 vccd1 _2149_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4627_ _0424_ _0397_ _1106_ _1107_ _1108_ vssd1 vssd1 vccd1 vccd1 _1109_ sky130_fd_sc_hd__o2111a_1
X_4558_ _3086_ _3141_ vssd1 vssd1 vccd1 vccd1 _1040_ sky130_fd_sc_hd__or2_1
X_4489_ _0372_ _0362_ _0691_ _0366_ _0971_ vssd1 vssd1 vccd1 vccd1 _0972_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ _3046_ vssd1 vssd1 vccd1 vccd1 _0301_ sky130_fd_sc_hd__clkbuf_1
X_6228_ _2597_ _2598_ _2599_ vssd1 vssd1 vccd1 vccd1 _2600_ sky130_fd_sc_hd__a21bo_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _2549_ _2529_ vssd1 vssd1 vccd1 vccd1 _2550_ sky130_fd_sc_hd__and2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3860_ egd_top.BitStream_buffer.BS_buffer\[37\] vssd1 vssd1 vccd1 vccd1 _0346_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3791_ _3103_ _3300_ vssd1 vssd1 vccd1 vccd1 _3325_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5530_ _0756_ _0584_ vssd1 vssd1 vccd1 vccd1 _2005_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5461_ _1934_ _1935_ vssd1 vssd1 vccd1 vccd1 _1936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4412_ _0828_ _0894_ _0895_ vssd1 vssd1 vccd1 vccd1 _0896_ sky130_fd_sc_hd__nand3_1
XFILLER_0_41_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5392_ _0479_ _0488_ _0482_ _0492_ _1867_ vssd1 vssd1 vccd1 vccd1 _1868_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4343_ _0814_ _0818_ _0823_ _0826_ vssd1 vssd1 vccd1 vccd1 _0827_ sky130_fd_sc_hd__and4_1
X_4274_ _0747_ _0752_ _0755_ _0758_ vssd1 vssd1 vccd1 vccd1 _0759_ sky130_fd_sc_hd__and4_1
X_6013_ _2449_ vssd1 vssd1 vccd1 vccd1 _0248_ sky130_fd_sc_hd__clkbuf_1
X_6628__118 clknet_1_0__leaf__2918_ vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__inv_2
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6915_ net36 _0318_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6846_ net44 _0249_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[30\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6777_ net131 _0180_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.pc_previous\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_5728_ _0423_ _0378_ _0421_ _0382_ _2200_ vssd1 vssd1 vccd1 vccd1 _2201_ sky130_fd_sc_hd__a221oi_1
X_3989_ egd_top.BitStream_buffer.BS_buffer\[25\] vssd1 vssd1 vccd1 vccd1 _0475_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5659_ _2132_ _2996_ _2937_ vssd1 vssd1 vccd1 vccd1 _2133_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4961_ _1436_ _1437_ _1438_ _1439_ vssd1 vssd1 vccd1 vccd1 _1440_ sky130_fd_sc_hd__and4_1
X_4892_ _1356_ _1371_ vssd1 vssd1 vccd1 vccd1 _1372_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3912_ _3131_ _0395_ vssd1 vssd1 vccd1 vccd1 _0398_ sky130_fd_sc_hd__and2_1
X_3843_ egd_top.BitStream_buffer.BS_buffer\[43\] vssd1 vssd1 vccd1 vccd1 _0329_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6673__160 clknet_1_0__leaf__2921_ vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__inv_2
X_6562_ _2889_ _2895_ _2756_ vssd1 vssd1 vccd1 vccd1 _2896_ sky130_fd_sc_hd__nand3_1
X_3774_ _3090_ _3300_ vssd1 vssd1 vccd1 vccd1 _3308_ sky130_fd_sc_hd__and2_1
X_5513_ _0508_ _0363_ vssd1 vssd1 vccd1 vccd1 _1988_ sky130_fd_sc_hd__nand2_1
X_6493_ _2828_ vssd1 vssd1 vccd1 vccd1 _2829_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6687__17 clknet_1_0__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__inv_2
X_5444_ egd_top.BitStream_buffer.BS_buffer\[9\] _3212_ egd_top.BitStream_buffer.BS_buffer\[10\]
+ _3215_ _1918_ vssd1 vssd1 vccd1 vccd1 _1919_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5375_ _0420_ _3129_ vssd1 vssd1 vccd1 vccd1 _1851_ sky130_fd_sc_hd__nand2_1
X_4326_ _0796_ _0801_ _0806_ _0809_ vssd1 vssd1 vccd1 vccd1 _0810_ sky130_fd_sc_hd__and4_1
X_4257_ _0548_ vssd1 vssd1 vccd1 vccd1 _0742_ sky130_fd_sc_hd__inv_2
X_4188_ _0668_ _3338_ _0669_ _0670_ _0672_ vssd1 vssd1 vccd1 vccd1 _0673_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6829_ net183 _0232_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[47\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3490_ net14 _3031_ _3007_ vssd1 vssd1 vccd1 vccd1 _3032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5160_ _0890_ _0556_ vssd1 vssd1 vccd1 vccd1 _1638_ sky130_fd_sc_hd__or2_1
X_4111_ _3153_ _0543_ vssd1 vssd1 vccd1 vccd1 _0597_ sky130_fd_sc_hd__nand2_1
X_5091_ _3345_ _3281_ _3335_ _3285_ _1568_ vssd1 vssd1 vccd1 vccd1 _1569_ sky130_fd_sc_hd__a221oi_1
X_4042_ _0527_ vssd1 vssd1 vccd1 vccd1 _0528_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _2435_ _2423_ vssd1 vssd1 vccd1 vccd1 _2436_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _3188_ _3176_ _3216_ _3179_ vssd1 vssd1 vccd1 vccd1 _1423_ sky130_fd_sc_hd__o22ai_1
X_6598__90 clknet_1_1__leaf__2916_ vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__inv_2
XFILLER_0_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4875_ _0429_ _0379_ _0433_ _0383_ _1354_ vssd1 vssd1 vccd1 vccd1 _1355_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3826_ _3359_ vssd1 vssd1 vccd1 vccd1 _3360_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ _3290_ vssd1 vssd1 vccd1 vccd1 _3291_ sky130_fd_sc_hd__inv_2
X_6545_ _1652_ _2720_ _1406_ vssd1 vssd1 vccd1 vccd1 _2879_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6476_ _2816_ _2756_ vssd1 vssd1 vccd1 vccd1 _2817_ sky130_fd_sc_hd__nand2_1
X_3688_ _3216_ _3218_ _3219_ _3221_ vssd1 vssd1 vccd1 vccd1 _3222_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5427_ _3133_ _3247_ vssd1 vssd1 vccd1 vccd1 _1902_ sky130_fd_sc_hd__nand2_1
X_5358_ _1832_ _1833_ vssd1 vssd1 vccd1 vccd1 _1834_ sky130_fd_sc_hd__nand2_1
X_4309_ _0782_ _0785_ _0789_ _0792_ vssd1 vssd1 vccd1 vccd1 _0793_ sky130_fd_sc_hd__and4_1
X_5289_ _0593_ _0584_ vssd1 vssd1 vccd1 vccd1 _1766_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__2920_ clknet_0__2920_ vssd1 vssd1 vccd1 vccd1 clknet_1_0__leaf__2920_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4660_ _0559_ _0556_ vssd1 vssd1 vccd1 vccd1 _1142_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3611_ _2954_ _3058_ vssd1 vssd1 vccd1 vccd1 _3145_ sky130_fd_sc_hd__nor2_2
XFILLER_0_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4591_ _3309_ _3357_ vssd1 vssd1 vccd1 vccd1 _1073_ sky130_fd_sc_hd__nand2_1
X_6330_ _2672_ _1894_ vssd1 vssd1 vccd1 vccd1 _2673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3542_ egd_top.BitStream_buffer.BS_buffer\[72\] vssd1 vssd1 vccd1 vccd1 _3076_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3473_ egd_top.BitStream_buffer.BS_buffer\[116\] vssd1 vssd1 vccd1 vccd1 _3019_ sky130_fd_sc_hd__clkbuf_4
X_6261_ net5 _3259_ _2613_ vssd1 vssd1 vccd1 vccd1 _2618_ sky130_fd_sc_hd__mux2_1
X_6192_ _2572_ _2554_ vssd1 vssd1 vccd1 vccd1 _2573_ sky130_fd_sc_hd__and2_1
X_5212_ _1687_ _1688_ vssd1 vssd1 vccd1 vccd1 _1689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5143_ _0478_ _0689_ _0481_ _0372_ vssd1 vssd1 vccd1 vccd1 _1621_ sky130_fd_sc_hd__a22o_1
X_5074_ _3206_ _3034_ vssd1 vssd1 vccd1 vccd1 _1552_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4025_ _3126_ _0470_ vssd1 vssd1 vccd1 vccd1 _0511_ sky130_fd_sc_hd__and2_1
X_5976_ _2424_ vssd1 vssd1 vccd1 vccd1 _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4927_ _1406_ _0898_ _2938_ vssd1 vssd1 vccd1 vccd1 _1407_ sky130_fd_sc_hd__a21oi_1
X_4858_ _3177_ _3363_ _1337_ vssd1 vssd1 vccd1 vccd1 _1338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3809_ _3131_ _3300_ vssd1 vssd1 vccd1 vccd1 _3343_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4789_ _0563_ egd_top.BitStream_buffer.BS_buffer\[15\] vssd1 vssd1 vccd1 vccd1 _1270_
+ sky130_fd_sc_hd__nand2_1
X_6528_ _2861_ _2862_ _2710_ vssd1 vssd1 vccd1 vccd1 _2863_ sky130_fd_sc_hd__nand3_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6459_ _2795_ _2799_ _2710_ vssd1 vssd1 vccd1 vccd1 _2800_ sky130_fd_sc_hd__nand3_1
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6592__85 clknet_1_1__leaf__2915_ vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__inv_2
XFILLER_0_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5830_ _3177_ _3337_ _2299_ _2300_ _2301_ vssd1 vssd1 vccd1 vccd1 _2302_ sky130_fd_sc_hd__o2111a_1
X_5761_ _2222_ _2225_ _2229_ _2233_ vssd1 vssd1 vccd1 vccd1 _2234_ sky130_fd_sc_hd__and4_1
XFILLER_0_71_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4712_ _3239_ _3264_ _0642_ _3268_ vssd1 vssd1 vccd1 vccd1 _1193_ sky130_fd_sc_hd__o22ai_1
X_5692_ _2161_ _2162_ _2163_ _2164_ vssd1 vssd1 vccd1 vccd1 _2165_ sky130_fd_sc_hd__and4_1
X_4643_ _0478_ _0521_ _0481_ _0525_ vssd1 vssd1 vccd1 vccd1 _1125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4574_ _0926_ _3218_ _0578_ _3221_ vssd1 vssd1 vccd1 vccd1 _1056_ sky130_fd_sc_hd__o22ai_1
X_3525_ _3058_ vssd1 vssd1 vccd1 vccd1 _3059_ sky130_fd_sc_hd__inv_2
X_6313_ _2655_ vssd1 vssd1 vccd1 vccd1 _2656_ sky130_fd_sc_hd__inv_2
X_6676__6 clknet_1_1__leaf__2922_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__inv_2
XFILLER_0_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _2595_ _2596_ vssd1 vssd1 vccd1 vccd1 _2608_ sky130_fd_sc_hd__nand2_2
X_3456_ _3005_ vssd1 vssd1 vccd1 vccd1 _3006_ sky130_fd_sc_hd__buf_2
X_6175_ _2561_ vssd1 vssd1 vccd1 vccd1 _0198_ sky130_fd_sc_hd__clkbuf_1
X_3387_ _2942_ net32 _2937_ vssd1 vssd1 vccd1 vccd1 _2943_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5126_ _0403_ _0447_ vssd1 vssd1 vccd1 vccd1 _1604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5057_ _3114_ _3085_ vssd1 vssd1 vccd1 vccd1 _1535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4008_ _0493_ vssd1 vssd1 vccd1 vccd1 _0494_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5959_ net1 egd_top.BitStream_buffer.BS_buffer\[15\] _2379_ vssd1 vssd1 vccd1 vccd1
+ _2412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _1814_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4290_ _3086_ _3124_ _0771_ _0772_ _0773_ vssd1 vssd1 vccd1 vccd1 _0774_ sky130_fd_sc_hd__o2111a_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6862_ net60 _0265_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_5813_ _1196_ _3263_ _1320_ _3267_ vssd1 vssd1 vccd1 vccd1 _2285_ sky130_fd_sc_hd__o22ai_1
X_6793_ net147 _0196_ vssd1 vssd1 vccd1 vccd1 egd_top.BitStream_buffer.BS_buffer\[99\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5744_ _2206_ _2210_ _2213_ _2216_ vssd1 vssd1 vccd1 vccd1 _2217_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5675_ _0578_ _3175_ _0574_ _3178_ vssd1 vssd1 vccd1 vccd1 _2148_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4626_ _0412_ _0408_ vssd1 vssd1 vccd1 vccd1 _1108_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4557_ _3133_ _3057_ vssd1 vssd1 vccd1 vccd1 _1039_ sky130_fd_sc_hd__nand2_1
X_4488_ _0347_ _0369_ _0970_ vssd1 vssd1 vccd1 vccd1 _0971_ sky130_fd_sc_hd__o21ai_1
X_3508_ _3045_ _3042_ vssd1 vssd1 vccd1 vccd1 _3046_ sky130_fd_sc_hd__and2_1
X_3439_ _2988_ _2953_ vssd1 vssd1 vccd1 vccd1 _2992_ sky130_fd_sc_hd__nand2_1
X_6227_ egd_top.BitStream_buffer.pc_previous\[3\] egd_top.BitStream_buffer.exp_golomb_len\[3\]
+ vssd1 vssd1 vccd1 vccd1 _2599_ sky130_fd_sc_hd__nand2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ net9 _3156_ _2520_ vssd1 vssd1 vccd1 vccd1 _2549_ sky130_fd_sc_hd__mux2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _1546_ _1557_ _1570_ _1586_ vssd1 vssd1 vccd1 vccd1 _1587_ sky130_fd_sc_hd__and4_1
X_6089_ _2932_ vssd1 vssd1 vccd1 vccd1 _2502_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6651__139 clknet_1_0__leaf__2920_ vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__inv_2
XFILLER_0_16_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 la_data_out_26_24[2] sky130_fd_sc_hd__buf_12
XFILLER_0_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3790_ _3323_ vssd1 vssd1 vccd1 vccd1 _3324_ sky130_fd_sc_hd__clkbuf_4
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5460_ _3313_ _3016_ vssd1 vssd1 vccd1 vccd1 _1935_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4411_ _0606_ _0573_ vssd1 vssd1 vccd1 vccd1 _0895_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5391_ _1123_ _0496_ _1866_ vssd1 vssd1 vccd1 vccd1 _1867_ sky130_fd_sc_hd__o21ai_1
X_4342_ _0674_ _3356_ _0675_ _3360_ _0825_ vssd1 vssd1 vccd1 vccd1 _0826_ sky130_fd_sc_hd__a221oi_1
X_4273_ egd_top.BitStream_buffer.BS_buffer\[15\] _0589_ egd_top.BitStream_buffer.BS_buffer\[16\]
+ _0592_ _0757_ vssd1 vssd1 vccd1 vccd1 _0758_ sky130_fd_sc_hd__a221oi_1
X_6012_ _2447_ _2448_ vssd1 vssd1 vccd1 vccd1 _2449_ sky130_fd_sc_hd__and2_1
.ends

