magic
tech sky130B
magscale 1 2
timestamp 1676037725
<< via4 >>
rect 1355 33227 1591 33463
rect 1675 33227 1911 33463
rect 1995 33227 2231 33463
rect 2315 33227 2551 33463
rect 2635 33227 2871 33463
rect 2955 33227 3191 33463
rect 3275 33227 3511 33463
rect 3595 33227 3831 33463
rect 3915 33227 4151 33463
rect 4235 33227 4471 33463
rect 4555 33227 4791 33463
rect 4875 33227 5111 33463
rect 5195 33227 5431 33463
rect 5515 33227 5751 33463
rect 5835 33227 6071 33463
rect 6155 33227 6391 33463
rect 6475 33227 6711 33463
rect 6795 33227 7031 33463
rect 7115 33227 7351 33463
rect 7435 33227 7671 33463
rect 7755 33227 7991 33463
rect 8075 33227 8311 33463
rect 8395 33227 8631 33463
rect 8715 33227 8951 33463
rect 9035 33227 9271 33463
rect 9355 33227 9591 33463
rect 9675 33227 9911 33463
rect 9995 33227 10231 33463
rect 10315 33227 10551 33463
rect 10635 33227 10871 33463
rect 10955 33227 11191 33463
rect 11275 33227 11511 33463
rect 11595 33227 11831 33463
rect 11915 33227 12151 33463
rect 12235 33227 12471 33463
rect 12555 33227 12791 33463
rect 12875 33227 13111 33463
rect 13195 33227 13431 33463
rect 13515 33227 13751 33463
rect 992 32958 1228 33194
rect 13838 32904 14074 33140
rect 672 32638 908 32874
rect 14158 32584 14394 32820
rect 352 32318 588 32554
rect 14478 32264 14714 32500
rect -10 31956 226 32192
rect 14786 31942 15022 32178
rect -10 31636 226 31872
rect 14786 31622 15022 31858
rect -10 31316 226 31552
rect 14786 31302 15022 31538
rect -10 30996 226 31232
rect 14786 30982 15022 31218
rect -10 30676 226 30912
rect 14786 30662 15022 30898
rect -10 30356 226 30592
rect 14786 30342 15022 30578
rect -10 30036 226 30272
rect 14786 30022 15022 30258
rect -10 29716 226 29952
rect 14786 29702 15022 29938
rect -10 29396 226 29632
rect 14786 29382 15022 29618
rect -10 29076 226 29312
rect 14786 29062 15022 29298
rect -10 28756 226 28992
rect 14786 28742 15022 28978
rect -10 28436 226 28672
rect 14786 28422 15022 28658
rect -10 28116 226 28352
rect 14786 28102 15022 28338
rect -10 27796 226 28032
rect 14786 27782 15022 28018
rect -10 27476 226 27712
rect 14786 27462 15022 27698
rect -10 27156 226 27392
rect 14786 27142 15022 27378
rect -10 26836 226 27072
rect 14786 26822 15022 27058
rect -10 26516 226 26752
rect 14786 26502 15022 26738
rect -10 26196 226 26432
rect 14786 26182 15022 26418
rect -10 25876 226 26112
rect 14786 25862 15022 26098
rect -10 25556 226 25792
rect 14786 25542 15022 25778
rect -10 25236 226 25472
rect 14786 25222 15022 25458
rect -10 24916 226 25152
rect 14786 24902 15022 25138
rect -10 24596 226 24832
rect 14786 24582 15022 24818
rect -10 24276 226 24512
rect 14786 24262 15022 24498
rect -10 23956 226 24192
rect 14786 23942 15022 24178
rect -10 23636 226 23872
rect 14786 23622 15022 23858
rect -10 23316 226 23552
rect 14786 23302 15022 23538
rect -10 22996 226 23232
rect 14786 22982 15022 23218
rect -10 22676 226 22912
rect 14786 22662 15022 22898
rect -10 22356 226 22592
rect 14786 22342 15022 22578
rect -10 22036 226 22272
rect 14786 22022 15022 22258
rect -10 21716 226 21952
rect 14786 21702 15022 21938
rect 298 21394 534 21630
rect 14424 21340 14660 21576
rect 618 21074 854 21310
rect 14104 21020 14340 21256
rect 938 20754 1174 20990
rect 13784 20700 14020 20936
rect 1261 20431 1497 20667
rect 1581 20431 1817 20667
rect 1901 20431 2137 20667
rect 2221 20431 2457 20667
rect 2541 20431 2777 20667
rect 2861 20431 3097 20667
rect 3181 20431 3417 20667
rect 3501 20431 3737 20667
rect 3821 20431 4057 20667
rect 4141 20431 4377 20667
rect 4461 20431 4697 20667
rect 4781 20431 5017 20667
rect 5101 20431 5337 20667
rect 5421 20431 5657 20667
rect 5741 20431 5977 20667
rect 6061 20431 6297 20667
rect 6381 20431 6617 20667
rect 6701 20431 6937 20667
rect 7021 20431 7257 20667
rect 7341 20431 7577 20667
rect 7661 20431 7897 20667
rect 7981 20431 8217 20667
rect 8301 20431 8537 20667
rect 8621 20431 8857 20667
rect 8941 20431 9177 20667
rect 9261 20431 9497 20667
rect 9581 20431 9817 20667
rect 9901 20431 10137 20667
rect 10221 20431 10457 20667
rect 10541 20431 10777 20667
rect 10861 20431 11097 20667
rect 11181 20431 11417 20667
rect 11501 20431 11737 20667
rect 11821 20431 12057 20667
rect 12141 20431 12377 20667
rect 12461 20431 12697 20667
rect 12781 20431 13017 20667
rect 13101 20431 13337 20667
rect 13421 20431 13657 20667
use sky130_fd_pr__padplhp__example_559591418080  sky130_fd_pr__padplhp__example_559591418080_0
timestamp 1676037725
transform 0 -1 14506 1 0 20947
box -540 -540 12540 14540
<< properties >>
string GDS_END 31364778
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31364688
<< end >>
